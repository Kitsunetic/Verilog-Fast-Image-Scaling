
module bufferram (
  input [15:0] addra,      
  output reg [15:0] douta 
);

always@(*) begin
  case(addra)
0: douta=16'h6457;
1: douta=16'h53f5;
2: douta=16'h9517;
3: douta=16'h5311;
4: douta=16'had98;
5: douta=16'h8455;
6: douta=16'h8c95;
7: douta=16'h84d7;
8: douta=16'hbdd8;
9: douta=16'ha598;
10: douta=16'hbdb6;
11: douta=16'h73f2;
12: douta=16'h73b2;
13: douta=16'h4333;
14: douta=16'hbe7a;
15: douta=16'h9d36;
16: douta=16'hd658;
17: douta=16'hd6b9;
18: douta=16'h3b11;
19: douta=16'hc5f8;
20: douta=16'hc67a;
21: douta=16'h2af0;
22: douta=16'h9d58;
23: douta=16'h8c95;
24: douta=16'h84d6;
25: douta=16'h8538;
26: douta=16'h9599;
27: douta=16'hbe39;
28: douta=16'h3b32;
29: douta=16'hce59;
30: douta=16'ha536;
31: douta=16'h21cd;
32: douta=16'had55;
33: douta=16'h2188;
34: douta=16'ha555;
35: douta=16'h5aee;
36: douta=16'h9cd3;
37: douta=16'h8c51;
38: douta=16'h634e;
39: douta=16'hbdb5;
40: douta=16'h8c71;
41: douta=16'h636f;
42: douta=16'h73d0;
43: douta=16'h6391;
44: douta=16'h2989;
45: douta=16'h9cf3;
46: douta=16'h2105;
47: douta=16'h3a4c;
48: douta=16'h52ce;
49: douta=16'h7bf1;
50: douta=16'h9d37;
51: douta=16'h2a2d;
52: douta=16'hbdb7;
53: douta=16'h4b31;
54: douta=16'h6c34;
55: douta=16'h19ee;
56: douta=16'h4b31;
57: douta=16'h8d18;
58: douta=16'h21ce;
59: douta=16'h8d18;
60: douta=16'h6435;
61: douta=16'h5c15;
62: douta=16'h53d5;
63: douta=16'h5bf7;
64: douta=16'h4bf6;
65: douta=16'h7cd8;
66: douta=16'h5351;
67: douta=16'had98;
68: douta=16'h5bd3;
69: douta=16'h6bf1;
70: douta=16'h9d78;
71: douta=16'h5372;
72: douta=16'he6da;
73: douta=16'h9495;
74: douta=16'had97;
75: douta=16'hbdd8;
76: douta=16'h7c53;
77: douta=16'ha4f5;
78: douta=16'h6415;
79: douta=16'he73a;
80: douta=16'h5c36;
81: douta=16'h9515;
82: douta=16'hce7a;
83: douta=16'h63f3;
84: douta=16'ha557;
85: douta=16'heed9;
86: douta=16'h84f7;
87: douta=16'h8d38;
88: douta=16'h7c14;
89: douta=16'h7454;
90: douta=16'h6c98;
91: douta=16'h7434;
92: douta=16'h9577;
93: douta=16'h5331;
94: douta=16'h9536;
95: douta=16'had76;
96: douta=16'h3a4c;
97: douta=16'hef3a;
98: douta=16'h0885;
99: douta=16'h738f;
100: douta=16'hce14;
101: douta=16'ha512;
102: douta=16'h31ec;
103: douta=16'had75;
104: douta=16'h8433;
105: douta=16'h0063;
106: douta=16'ha575;
107: douta=16'h21cb;
108: douta=16'h63f2;
109: douta=16'h8473;
110: douta=16'h18a3;
111: douta=16'h2189;
112: douta=16'h7c12;
113: douta=16'h52cd;
114: douta=16'hff58;
115: douta=16'h3a4c;
116: douta=16'h9d57;
117: douta=16'h9539;
118: douta=16'h3aaf;
119: douta=16'h5bf5;
120: douta=16'h3af0;
121: douta=16'hc639;
122: douta=16'h32d2;
123: douta=16'h8d19;
124: douta=16'h63f5;
125: douta=16'h7497;
126: douta=16'h5438;
127: douta=16'ha5da;
128: douta=16'h53f6;
129: douta=16'h6436;
130: douta=16'h7414;
131: douta=16'hadfb;
132: douta=16'h8452;
133: douta=16'hce59;
134: douta=16'h5352;
135: douta=16'had56;
136: douta=16'h8474;
137: douta=16'hb598;
138: douta=16'h7413;
139: douta=16'h83f2;
140: douta=16'he6ba;
141: douta=16'h4aee;
142: douta=16'hbd95;
143: douta=16'had75;
144: douta=16'h6370;
145: douta=16'hb5b7;
146: douta=16'hbe18;
147: douta=16'hbdf9;
148: douta=16'h1a0e;
149: douta=16'ha5b9;
150: douta=16'h95ba;
151: douta=16'h4b51;
152: douta=16'had97;
153: douta=16'h6c96;
154: douta=16'h9d78;
155: douta=16'hb619;
156: douta=16'h4b74;
157: douta=16'h9d36;
158: douta=16'h6bd1;
159: douta=16'h7c53;
160: douta=16'hb5b8;
161: douta=16'h530e;
162: douta=16'h424a;
163: douta=16'h18e3;
164: douta=16'h29a8;
165: douta=16'ha4f4;
166: douta=16'h320b;
167: douta=16'hbd33;
168: douta=16'h7c31;
169: douta=16'hce37;
170: douta=16'h3a2c;
171: douta=16'ha536;
172: douta=16'h5b70;
173: douta=16'hbdd7;
174: douta=16'h1083;
175: douta=16'h7413;
176: douta=16'h73f3;
177: douta=16'h5350;
178: douta=16'h94d4;
179: douta=16'h328f;
180: douta=16'h42ad;
181: douta=16'h9517;
182: douta=16'h6392;
183: douta=16'h7436;
184: douta=16'h7cda;
185: douta=16'h2a2d;
186: douta=16'h84f9;
187: douta=16'h5b93;
188: douta=16'h5b52;
189: douta=16'h118b;
190: douta=16'h5bb5;
191: douta=16'h3b33;
192: douta=16'h6498;
193: douta=16'h4352;
194: douta=16'h8518;
195: douta=16'h426e;
196: douta=16'hc5d7;
197: douta=16'h8cb4;
198: douta=16'h6bd2;
199: douta=16'hbe38;
200: douta=16'h5b30;
201: douta=16'hf75a;
202: douta=16'h9493;
203: douta=16'hdeb9;
204: douta=16'h8c11;
205: douta=16'h8c30;
206: douta=16'h83f2;
207: douta=16'h8451;
208: douta=16'hd657;
209: douta=16'h4350;
210: douta=16'h9d98;
211: douta=16'h9517;
212: douta=16'hd67a;
213: douta=16'h32f3;
214: douta=16'h84d7;
215: douta=16'hce7b;
216: douta=16'h6c77;
217: douta=16'h8495;
218: douta=16'hbe9c;
219: douta=16'hbe5b;
220: douta=16'hc639;
221: douta=16'h6bd2;
222: douta=16'h6391;
223: douta=16'hd5f8;
224: douta=16'h8473;
225: douta=16'h5b70;
226: douta=16'h1926;
227: douta=16'h2124;
228: douta=16'h5b0e;
229: douta=16'h634e;
230: douta=16'h9492;
231: douta=16'h8cb3;
232: douta=16'h6370;
233: douta=16'h1127;
234: douta=16'h0863;
235: douta=16'h08a4;
236: douta=16'h10c4;
237: douta=16'h0884;
238: douta=16'h0883;
239: douta=16'h0863;
240: douta=16'h0062;
241: douta=16'h0001;
242: douta=16'h42ad;
243: douta=16'h6436;
244: douta=16'h2a2d;
245: douta=16'hd67a;
246: douta=16'h3af2;
247: douta=16'h222e;
248: douta=16'h7476;
249: douta=16'h5351;
250: douta=16'h9517;
251: douta=16'h32f1;
252: douta=16'h6416;
253: douta=16'h3b13;
254: douta=16'h959c;
255: douta=16'h2ad2;
256: douta=16'h3af1;
257: douta=16'h84f9;
258: douta=16'h5331;
259: douta=16'h6350;
260: douta=16'ha555;
261: douta=16'h7413;
262: douta=16'ha576;
263: douta=16'h9516;
264: douta=16'h9cf3;
265: douta=16'hd699;
266: douta=16'ha514;
267: douta=16'hded9;
268: douta=16'hce16;
269: douta=16'h8411;
270: douta=16'hc5d4;
271: douta=16'h8431;
272: douta=16'h94b2;
273: douta=16'hbd75;
274: douta=16'h4b50;
275: douta=16'ha5b8;
276: douta=16'hb577;
277: douta=16'hb63b;
278: douta=16'h7497;
279: douta=16'h32b0;
280: douta=16'h9578;
281: douta=16'ha61b;
282: douta=16'h7c96;
283: douta=16'h8518;
284: douta=16'hadfa;
285: douta=16'h9cd3;
286: douta=16'h8d37;
287: douta=16'h5330;
288: douta=16'h8d77;
289: douta=16'h7cb5;
290: douta=16'h5b72;
291: douta=16'h6b4d;
292: douta=16'h5b0d;
293: douta=16'h4aac;
294: douta=16'h10e4;
295: douta=16'h10e5;
296: douta=16'h0862;
297: douta=16'h3a2b;
298: douta=16'h5b72;
299: douta=16'h63f6;
300: douta=16'h6c57;
301: douta=16'h6c98;
302: douta=16'h7cf9;
303: douta=16'h6c57;
304: douta=16'h5b93;
305: douta=16'h322d;
306: douta=16'h10e5;
307: douta=16'h0883;
308: douta=16'h08c4;
309: douta=16'h29e9;
310: douta=16'h6c54;
311: douta=16'h1128;
312: douta=16'h63f3;
313: douta=16'h5b72;
314: douta=16'h116a;
315: douta=16'h7455;
316: douta=16'h5b92;
317: douta=16'h5c58;
318: douta=16'h6cb9;
319: douta=16'h959b;
320: douta=16'h6416;
321: douta=16'h42cf;
322: douta=16'h6371;
323: douta=16'h8c74;
324: douta=16'ha536;
325: douta=16'hd658;
326: douta=16'h6c34;
327: douta=16'h7433;
328: douta=16'hef3a;
329: douta=16'hd678;
330: douta=16'hd698;
331: douta=16'hce37;
332: douta=16'hef5a;
333: douta=16'h83ae;
334: douta=16'he6b8;
335: douta=16'h4aad;
336: douta=16'hc5d4;
337: douta=16'h9450;
338: douta=16'h8431;
339: douta=16'h5b50;
340: douta=16'had96;
341: douta=16'hc658;
342: douta=16'h6bd3;
343: douta=16'h6477;
344: douta=16'h5c15;
345: douta=16'h4b73;
346: douta=16'h855a;
347: douta=16'h53d4;
348: douta=16'h3aaf;
349: douta=16'hbe59;
350: douta=16'hbe3a;
351: douta=16'h4aad;
352: douta=16'h7c96;
353: douta=16'h3a4e;
354: douta=16'h6c35;
355: douta=16'h1127;
356: douta=16'h1905;
357: douta=16'h39c8;
358: douta=16'h7c55;
359: douta=16'h855a;
360: douta=16'ha61c;
361: douta=16'h74d9;
362: douta=16'h6c98;
363: douta=16'h6478;
364: douta=16'h6458;
365: douta=16'h6c98;
366: douta=16'h74d9;
367: douta=16'h74d9;
368: douta=16'h8d9b;
369: douta=16'h751a;
370: douta=16'h6498;
371: douta=16'h7d3b;
372: douta=16'h74fa;
373: douta=16'h29eb;
374: douta=16'h10c5;
375: douta=16'h0064;
376: douta=16'h7c53;
377: douta=16'h8cb6;
378: douta=16'h6bd3;
379: douta=16'h5b72;
380: douta=16'h3ad0;
381: douta=16'h6c56;
382: douta=16'h53d5;
383: douta=16'h53d4;
384: douta=16'h6415;
385: douta=16'h6c57;
386: douta=16'h6bd4;
387: douta=16'h6bf4;
388: douta=16'h5b92;
389: douta=16'had97;
390: douta=16'hb5b7;
391: douta=16'hffdb;
392: douta=16'ha534;
393: douta=16'hff7b;
394: douta=16'h4acd;
395: douta=16'hde98;
396: douta=16'hce57;
397: douta=16'hbd74;
398: douta=16'ha4d0;
399: douta=16'h5b0c;
400: douta=16'h840f;
401: douta=16'h94b2;
402: douta=16'hde77;
403: douta=16'h5aaa;
404: douta=16'h3a2a;
405: douta=16'h324d;
406: douta=16'h5bb3;
407: douta=16'h5372;
408: douta=16'h4311;
409: douta=16'h4bd6;
410: douta=16'h5395;
411: douta=16'h53d5;
412: douta=16'h53f5;
413: douta=16'h42b0;
414: douta=16'h4b11;
415: douta=16'ha578;
416: douta=16'h324e;
417: douta=16'h5b71;
418: douta=16'h2966;
419: douta=16'h7b6e;
420: douta=16'h8519;
421: douta=16'h851a;
422: douta=16'h851a;
423: douta=16'h851a;
424: douta=16'h8d5b;
425: douta=16'h8d7b;
426: douta=16'h8d7b;
427: douta=16'h6cb9;
428: douta=16'h6c99;
429: douta=16'h7d3b;
430: douta=16'h7d3a;
431: douta=16'h7d3a;
432: douta=16'h855a;
433: douta=16'h6c99;
434: douta=16'h7d1a;
435: douta=16'h7d1a;
436: douta=16'h751a;
437: douta=16'h74d9;
438: douta=16'h751a;
439: douta=16'h29aa;
440: douta=16'h1107;
441: douta=16'h42ee;
442: douta=16'h19ab;
443: douta=16'h9d79;
444: douta=16'h5c38;
445: douta=16'h6c97;
446: douta=16'h6c57;
447: douta=16'h3b12;
448: douta=16'h7457;
449: douta=16'h5373;
450: douta=16'h7455;
451: douta=16'h73f3;
452: douta=16'h9d56;
453: douta=16'ha557;
454: douta=16'hc5f7;
455: douta=16'hb575;
456: douta=16'hbdb5;
457: douta=16'hde98;
458: douta=16'h73f0;
459: douta=16'hef19;
460: douta=16'hd655;
461: douta=16'hff38;
462: douta=16'hb510;
463: douta=16'h62cb;
464: douta=16'h18e5;
465: douta=16'h73ae;
466: douta=16'had32;
467: douta=16'h9cb0;
468: douta=16'h5b4e;
469: douta=16'h4a4b;
470: douta=16'h1082;
471: douta=16'h3aaf;
472: douta=16'h5393;
473: douta=16'h6c56;
474: douta=16'h4b53;
475: douta=16'h6bf2;
476: douta=16'h5352;
477: douta=16'h32b1;
478: douta=16'h63d3;
479: douta=16'ha599;
480: douta=16'h4aad;
481: douta=16'h41a6;
482: douta=16'h84f8;
483: douta=16'h7c97;
484: douta=16'h84f9;
485: douta=16'h84f9;
486: douta=16'h8d7b;
487: douta=16'h8d5a;
488: douta=16'h84d9;
489: douta=16'h8d5b;
490: douta=16'h74b8;
491: douta=16'h957b;
492: douta=16'h95bc;
493: douta=16'h74da;
494: douta=16'h859c;
495: douta=16'h8dbc;
496: douta=16'h855b;
497: douta=16'h859c;
498: douta=16'h7d3b;
499: douta=16'h8d9b;
500: douta=16'h7d3a;
501: douta=16'h753a;
502: douta=16'h7d7c;
503: douta=16'h74fa;
504: douta=16'h753b;
505: douta=16'h21a8;
506: douta=16'h32af;
507: douta=16'h63f5;
508: douta=16'haddb;
509: douta=16'h2a90;
510: douta=16'h8518;
511: douta=16'h8d5a;
512: douta=16'h4312;
513: douta=16'h2a70;
514: douta=16'h6bd4;
515: douta=16'h6bd2;
516: douta=16'h8c94;
517: douta=16'h8453;
518: douta=16'hd657;
519: douta=16'ha4d2;
520: douta=16'hf738;
521: douta=16'hc5b5;
522: douta=16'hde76;
523: douta=16'hce16;
524: douta=16'hb551;
525: douta=16'hde96;
526: douta=16'h62ca;
527: douta=16'h2167;
528: douta=16'h2988;
529: douta=16'h0084;
530: douta=16'h530c;
531: douta=16'h7bce;
532: douta=16'h4b31;
533: douta=16'h9472;
534: douta=16'h4b0f;
535: douta=16'h1061;
536: douta=16'h1061;
537: douta=16'h00e7;
538: douta=16'h3b31;
539: douta=16'h29ec;
540: douta=16'h4b31;
541: douta=16'h74b8;
542: douta=16'h6bd2;
543: douta=16'h52f0;
544: douta=16'h836c;
545: douta=16'h9d9a;
546: douta=16'h9519;
547: douta=16'h7456;
548: douta=16'h84d8;
549: douta=16'h84f9;
550: douta=16'h8d3a;
551: douta=16'h8519;
552: douta=16'h7cb9;
553: douta=16'h8d7b;
554: douta=16'h853a;
555: douta=16'h959c;
556: douta=16'h8d7a;
557: douta=16'h8519;
558: douta=16'h851a;
559: douta=16'h853a;
560: douta=16'h74fa;
561: douta=16'h7d7b;
562: douta=16'h8dbd;
563: douta=16'h95bc;
564: douta=16'h7d3a;
565: douta=16'h74fa;
566: douta=16'h6499;
567: douta=16'h74d9;
568: douta=16'h5c16;
569: douta=16'h6cb9;
570: douta=16'h29a8;
571: douta=16'h53d4;
572: douta=16'h5c16;
573: douta=16'h5392;
574: douta=16'h7456;
575: douta=16'h84d7;
576: douta=16'h5c57;
577: douta=16'h5bd5;
578: douta=16'h9d59;
579: douta=16'h5b70;
580: douta=16'hce39;
581: douta=16'had35;
582: douta=16'hde77;
583: douta=16'h6b4d;
584: douta=16'hde76;
585: douta=16'h52ed;
586: douta=16'hbdd3;
587: douta=16'hd636;
588: douta=16'hc614;
589: douta=16'h83ac;
590: douta=16'h62a9;
591: douta=16'h2167;
592: douta=16'h10e5;
593: douta=16'h18e5;
594: douta=16'h39a8;
595: douta=16'h63d2;
596: douta=16'h1927;
597: douta=16'h8430;
598: douta=16'h8474;
599: douta=16'h5370;
600: douta=16'h5393;
601: douta=16'h10e3;
602: douta=16'h428d;
603: douta=16'h4374;
604: douta=16'h3b11;
605: douta=16'h53b4;
606: douta=16'h6498;
607: douta=16'hacaf;
608: douta=16'h6478;
609: douta=16'h957a;
610: douta=16'h5bb5;
611: douta=16'h7c76;
612: douta=16'h6c36;
613: douta=16'h8d1a;
614: douta=16'h959b;
615: douta=16'h7cb8;
616: douta=16'h6c56;
617: douta=16'h851a;
618: douta=16'h8d7a;
619: douta=16'h7cd9;
620: douta=16'h8d5a;
621: douta=16'h8d3a;
622: douta=16'h8d3a;
623: douta=16'h8d5b;
624: douta=16'h851a;
625: douta=16'h855a;
626: douta=16'h8e1e;
627: douta=16'h6cfa;
628: douta=16'h857c;
629: douta=16'h857b;
630: douta=16'h74fa;
631: douta=16'h6458;
632: douta=16'h8d5b;
633: douta=16'h6cfa;
634: douta=16'h74fa;
635: douta=16'h1906;
636: douta=16'h5353;
637: douta=16'h19cc;
638: douta=16'h4b51;
639: douta=16'h42d0;
640: douta=16'h4333;
641: douta=16'h322e;
642: douta=16'h84b7;
643: douta=16'h7c35;
644: douta=16'hd69b;
645: douta=16'hbd95;
646: douta=16'hde97;
647: douta=16'h5aed;
648: douta=16'hbd94;
649: douta=16'h8c4f;
650: douta=16'hb530;
651: douta=16'hbd93;
652: douta=16'h8bcc;
653: douta=16'h9c0d;
654: douta=16'h6aea;
655: douta=16'h2987;
656: douta=16'h1926;
657: douta=16'h18e5;
658: douta=16'hacd0;
659: douta=16'h5b90;
660: douta=16'h634d;
661: douta=16'h29a9;
662: douta=16'h1106;
663: douta=16'h29cb;
664: douta=16'h3b10;
665: douta=16'h42f1;
666: douta=16'h4acd;
667: douta=16'h0820;
668: douta=16'h3a8f;
669: douta=16'h5c36;
670: douta=16'hd550;
671: douta=16'h5375;
672: douta=16'h853a;
673: douta=16'hae1c;
674: douta=16'h853a;
675: douta=16'ha5db;
676: douta=16'h7cb8;
677: douta=16'h9dbb;
678: douta=16'h7cd9;
679: douta=16'h9ddb;
680: douta=16'h957a;
681: douta=16'h7cd8;
682: douta=16'h74b8;
683: douta=16'h7cb8;
684: douta=16'h6c36;
685: douta=16'h8d5b;
686: douta=16'h95bc;
687: douta=16'h959c;
688: douta=16'h959b;
689: douta=16'h8d7b;
690: douta=16'h857b;
691: douta=16'h95bd;
692: douta=16'h857b;
693: douta=16'h751b;
694: douta=16'h751b;
695: douta=16'h6cb9;
696: douta=16'h7d5a;
697: douta=16'h8d7b;
698: douta=16'h857b;
699: douta=16'h74fa;
700: douta=16'h2189;
701: douta=16'h8cf5;
702: douta=16'h63b2;
703: douta=16'h8453;
704: douta=16'h4b95;
705: douta=16'h2a2e;
706: douta=16'h7c76;
707: douta=16'h8cb5;
708: douta=16'h9c93;
709: douta=16'h39eb;
710: douta=16'h9470;
711: douta=16'h9450;
712: douta=16'ha4d0;
713: douta=16'hb572;
714: douta=16'hce34;
715: douta=16'h8bac;
716: douta=16'h9c0c;
717: douta=16'hb4ad;
718: douta=16'hac6d;
719: douta=16'h6b0a;
720: douta=16'h18e5;
721: douta=16'h1905;
722: douta=16'h0883;
723: douta=16'h84b6;
724: douta=16'h4229;
725: douta=16'h632d;
726: douta=16'h428c;
727: douta=16'h6b6f;
728: douta=16'h1927;
729: douta=16'h6bd2;
730: douta=16'h328f;
731: douta=16'h3a4b;
732: douta=16'h18c3;
733: douta=16'h0860;
734: douta=16'h9579;
735: douta=16'h7cd7;
736: douta=16'h8d5a;
737: douta=16'h84f9;
738: douta=16'h7cd9;
739: douta=16'h8519;
740: douta=16'h84b8;
741: douta=16'ha5fc;
742: douta=16'h957a;
743: douta=16'h84f9;
744: douta=16'h8d5a;
745: douta=16'h8d3a;
746: douta=16'h7477;
747: douta=16'h8d5a;
748: douta=16'h6c15;
749: douta=16'h8d3a;
750: douta=16'h853a;
751: douta=16'h7cf9;
752: douta=16'h957b;
753: douta=16'h851a;
754: douta=16'h7d3a;
755: douta=16'h7d1b;
756: douta=16'h7d1a;
757: douta=16'h7cfa;
758: douta=16'h53b5;
759: douta=16'h8dfd;
760: douta=16'h6cba;
761: douta=16'h859c;
762: douta=16'h8dbc;
763: douta=16'h7d1a;
764: douta=16'h5b72;
765: douta=16'h8496;
766: douta=16'h6c13;
767: douta=16'h5331;
768: douta=16'h4312;
769: douta=16'h7477;
770: douta=16'h6bf3;
771: douta=16'h8cb5;
772: douta=16'hb535;
773: douta=16'h7b90;
774: douta=16'ha4f2;
775: douta=16'h944f;
776: douta=16'hbd92;
777: douta=16'hb531;
778: douta=16'h7309;
779: douta=16'h9c0d;
780: douta=16'hb4cd;
781: douta=16'hd570;
782: douta=16'hac4d;
783: douta=16'h5a68;
784: douta=16'h2967;
785: douta=16'h08a4;
786: douta=16'h10e4;
787: douta=16'h0000;
788: douta=16'h428b;
789: douta=16'h6b4d;
790: douta=16'h29ea;
791: douta=16'h73ae;
792: douta=16'h42ce;
793: douta=16'h29c9;
794: douta=16'h32ae;
795: douta=16'h3a4c;
796: douta=16'h5371;
797: douta=16'hb48d;
798: douta=16'h84d8;
799: douta=16'h7477;
800: douta=16'h7477;
801: douta=16'h8cf8;
802: douta=16'h8d3a;
803: douta=16'h7cb7;
804: douta=16'h84f8;
805: douta=16'h957b;
806: douta=16'h7d19;
807: douta=16'h95db;
808: douta=16'h7cd9;
809: douta=16'h8d7a;
810: douta=16'h8d39;
811: douta=16'h8d5a;
812: douta=16'h853a;
813: douta=16'h7477;
814: douta=16'h8d3a;
815: douta=16'h851a;
816: douta=16'h74b8;
817: douta=16'h6c77;
818: douta=16'h6436;
819: douta=16'h855b;
820: douta=16'h7d1a;
821: douta=16'h95dc;
822: douta=16'h7cfa;
823: douta=16'h857c;
824: douta=16'h8d9c;
825: douta=16'h7d3b;
826: douta=16'h7d5a;
827: douta=16'h7cf9;
828: douta=16'h7d3a;
829: douta=16'hb5d9;
830: douta=16'h8474;
831: douta=16'h73b0;
832: douta=16'h2a2e;
833: douta=16'h84b8;
834: douta=16'h7c75;
835: douta=16'h9d16;
836: douta=16'h7bf1;
837: douta=16'hc5f5;
838: douta=16'h8bee;
839: douta=16'heef8;
840: douta=16'hb531;
841: douta=16'h6ae9;
842: douta=16'h93eb;
843: douta=16'hb48d;
844: douta=16'hddf3;
845: douta=16'he634;
846: douta=16'hcd6f;
847: douta=16'h3165;
848: douta=16'h39e9;
849: douta=16'h29a8;
850: douta=16'h10a3;
851: douta=16'h2145;
852: douta=16'h1106;
853: douta=16'h10e5;
854: douta=16'h4208;
855: douta=16'h630d;
856: douta=16'h1948;
857: douta=16'h4aab;
858: douta=16'h3a09;
859: douta=16'h29ca;
860: douta=16'h530f;
861: douta=16'ha598;
862: douta=16'h9dbb;
863: douta=16'h8519;
864: douta=16'h7cd8;
865: douta=16'ha5dc;
866: douta=16'h9dbb;
867: douta=16'h9559;
868: douta=16'h8d3a;
869: douta=16'h853a;
870: douta=16'h959a;
871: douta=16'h7cd9;
872: douta=16'h6417;
873: douta=16'h959b;
874: douta=16'h955a;
875: douta=16'h853a;
876: douta=16'h7d3b;
877: douta=16'h7d1a;
878: douta=16'h6c57;
879: douta=16'h6c77;
880: douta=16'h6436;
881: douta=16'h6c15;
882: douta=16'h6415;
883: douta=16'h6c78;
884: douta=16'h6c78;
885: douta=16'h855c;
886: douta=16'h859c;
887: douta=16'h7cfa;
888: douta=16'h857b;
889: douta=16'h7d1a;
890: douta=16'h857c;
891: douta=16'h7d3a;
892: douta=16'h8dbc;
893: douta=16'h52cd;
894: douta=16'h63b2;
895: douta=16'h73d2;
896: douta=16'h2a90;
897: douta=16'h5352;
898: douta=16'h3a4e;
899: douta=16'h7c33;
900: douta=16'h94d3;
901: douta=16'hbd74;
902: douta=16'ha4b1;
903: douta=16'ha4d1;
904: douta=16'h8c0e;
905: douta=16'h836a;
906: douta=16'hb4ad;
907: douta=16'hcd90;
908: douta=16'he654;
909: douta=16'hd5b1;
910: douta=16'hb48e;
911: douta=16'hbd30;
912: douta=16'h6aec;
913: douta=16'h422a;
914: douta=16'h1926;
915: douta=16'h1905;
916: douta=16'h10c4;
917: douta=16'h1106;
918: douta=16'h29a7;
919: douta=16'h734c;
920: douta=16'h5aec;
921: douta=16'h1147;
922: douta=16'h426c;
923: douta=16'h0044;
924: douta=16'h2167;
925: douta=16'h8d39;
926: douta=16'h9d9a;
927: douta=16'hadfc;
928: douta=16'h6435;
929: douta=16'h957a;
930: douta=16'h957b;
931: douta=16'h8d5a;
932: douta=16'h959b;
933: douta=16'h7cd9;
934: douta=16'h6c77;
935: douta=16'hbe9e;
936: douta=16'h6c56;
937: douta=16'h6436;
938: douta=16'h6416;
939: douta=16'h6cb9;
940: douta=16'h6457;
941: douta=16'h4b53;
942: douta=16'h7497;
943: douta=16'h7c77;
944: douta=16'h7c96;
945: douta=16'h6c35;
946: douta=16'h5373;
947: douta=16'h3b13;
948: douta=16'h5c58;
949: douta=16'h6458;
950: douta=16'h74da;
951: douta=16'h74d9;
952: douta=16'h7d3a;
953: douta=16'h7d3b;
954: douta=16'h7499;
955: douta=16'h7cd9;
956: douta=16'h7d1a;
957: douta=16'h1906;
958: douta=16'h63d3;
959: douta=16'h6bb1;
960: douta=16'h3333;
961: douta=16'h53d4;
962: douta=16'h5331;
963: douta=16'h8c54;
964: douta=16'had56;
965: douta=16'h8c50;
966: douta=16'hd657;
967: douta=16'h8c71;
968: douta=16'h8bab;
969: douta=16'hac6b;
970: douta=16'hd56f;
971: douta=16'he675;
972: douta=16'hddf3;
973: douta=16'hbcae;
974: douta=16'hb4ae;
975: douta=16'hd5d2;
976: douta=16'hb4d0;
977: douta=16'h736e;
978: douta=16'h428c;
979: douta=16'h1906;
980: douta=16'h18a4;
981: douta=16'h08a4;
982: douta=16'h2988;
983: douta=16'h0001;
984: douta=16'h62aa;
985: douta=16'h6b4c;
986: douta=16'hb532;
987: douta=16'h636f;
988: douta=16'h7bef;
989: douta=16'h84b7;
990: douta=16'h9579;
991: douta=16'h8d39;
992: douta=16'ha5ba;
993: douta=16'h9d9a;
994: douta=16'h8d39;
995: douta=16'h9dbb;
996: douta=16'h95bb;
997: douta=16'h6c58;
998: douta=16'ha5fc;
999: douta=16'h8518;
1000: douta=16'h1925;
1001: douta=16'h4b32;
1002: douta=16'h7497;
1003: douta=16'h7cb7;
1004: douta=16'h6415;
1005: douta=16'h5b73;
1006: douta=16'h6c77;
1007: douta=16'h5bb3;
1008: douta=16'h9d9a;
1009: douta=16'h2967;
1010: douta=16'h7cd9;
1011: douta=16'h6cb9;
1012: douta=16'h6479;
1013: douta=16'h5c37;
1014: douta=16'h74f9;
1015: douta=16'h7d3a;
1016: douta=16'h6416;
1017: douta=16'h8d9c;
1018: douta=16'h7d1a;
1019: douta=16'h7cd9;
1020: douta=16'h853a;
1021: douta=16'h39ea;
1022: douta=16'h7413;
1023: douta=16'h9517;
1024: douta=16'h4b54;
1025: douta=16'h6458;
1026: douta=16'h63d4;
1027: douta=16'h5b92;
1028: douta=16'hb576;
1029: douta=16'hb534;
1030: douta=16'hce36;
1031: douta=16'h93cb;
1032: douta=16'hbc8b;
1033: douta=16'hd5b0;
1034: douta=16'hee75;
1035: douta=16'he674;
1036: douta=16'hc551;
1037: douta=16'h93ec;
1038: douta=16'hde13;
1039: douta=16'hddf3;
1040: douta=16'hcd50;
1041: douta=16'h8c10;
1042: douta=16'h6b70;
1043: douta=16'h42af;
1044: douta=16'h2988;
1045: douta=16'h10e4;
1046: douta=16'h10a4;
1047: douta=16'h3acf;
1048: douta=16'h2167;
1049: douta=16'h39a6;
1050: douta=16'h4228;
1051: douta=16'h942f;
1052: douta=16'h1105;
1053: douta=16'h5bb4;
1054: douta=16'h9579;
1055: douta=16'h8d18;
1056: douta=16'h8d18;
1057: douta=16'h957a;
1058: douta=16'h9d9a;
1059: douta=16'h9559;
1060: douta=16'ha5db;
1061: douta=16'h9d9a;
1062: douta=16'h9ddc;
1063: douta=16'h84f8;
1064: douta=16'h838b;
1065: douta=16'h8cf8;
1066: douta=16'h9d7a;
1067: douta=16'h8d39;
1068: douta=16'h8d39;
1069: douta=16'h8539;
1070: douta=16'h957a;
1071: douta=16'h63d3;
1072: douta=16'h8518;
1073: douta=16'h2146;
1074: douta=16'h5c16;
1075: douta=16'h6cb9;
1076: douta=16'h74da;
1077: douta=16'h74d9;
1078: douta=16'h74b9;
1079: douta=16'h7d1a;
1080: douta=16'h8d5b;
1081: douta=16'h851a;
1082: douta=16'h853b;
1083: douta=16'h8519;
1084: douta=16'h851a;
1085: douta=16'hdefd;
1086: douta=16'ha558;
1087: douta=16'h3a2a;
1088: douta=16'h3af2;
1089: douta=16'h3b12;
1090: douta=16'h5bb4;
1091: douta=16'h6392;
1092: douta=16'ha536;
1093: douta=16'h8411;
1094: douta=16'h834a;
1095: douta=16'hb4ac;
1096: douta=16'hd5b0;
1097: douta=16'hee75;
1098: douta=16'he634;
1099: douta=16'hbcf0;
1100: douta=16'hb4ce;
1101: douta=16'hc54f;
1102: douta=16'he634;
1103: douta=16'hde13;
1104: douta=16'hcd50;
1105: douta=16'ha471;
1106: douta=16'h8411;
1107: douta=16'h5b50;
1108: douta=16'h6372;
1109: douta=16'h2146;
1110: douta=16'h10e4;
1111: douta=16'h10a3;
1112: douta=16'h0042;
1113: douta=16'h840d;
1114: douta=16'h39a7;
1115: douta=16'h630c;
1116: douta=16'h2187;
1117: douta=16'h7c95;
1118: douta=16'h84f8;
1119: douta=16'h7c97;
1120: douta=16'h7456;
1121: douta=16'ha5ba;
1122: douta=16'h9579;
1123: douta=16'ha5da;
1124: douta=16'h9d9a;
1125: douta=16'ha5db;
1126: douta=16'ha5fb;
1127: douta=16'h959a;
1128: douta=16'h94f6;
1129: douta=16'h0042;
1130: douta=16'h8d39;
1131: douta=16'h957a;
1132: douta=16'h9d9a;
1133: douta=16'h9d99;
1134: douta=16'h8c75;
1135: douta=16'h7455;
1136: douta=16'h7cd8;
1137: douta=16'h10e5;
1138: douta=16'h6478;
1139: douta=16'h3b34;
1140: douta=16'h53f6;
1141: douta=16'h857b;
1142: douta=16'h7498;
1143: douta=16'h7cf9;
1144: douta=16'h7cd9;
1145: douta=16'h8d5a;
1146: douta=16'h853a;
1147: douta=16'h853a;
1148: douta=16'h8d7b;
1149: douta=16'hbe3a;
1150: douta=16'h9d16;
1151: douta=16'h5310;
1152: douta=16'h21ed;
1153: douta=16'h32f2;
1154: douta=16'h74b8;
1155: douta=16'h8497;
1156: douta=16'h5b30;
1157: douta=16'h8bcb;
1158: douta=16'hbcad;
1159: douta=16'hcd6f;
1160: douta=16'hee96;
1161: douta=16'heeb6;
1162: douta=16'hc50e;
1163: douta=16'h8b8a;
1164: douta=16'hc54f;
1165: douta=16'hde13;
1166: douta=16'hde14;
1167: douta=16'he613;
1168: douta=16'hbcf1;
1169: douta=16'h8c12;
1170: douta=16'h8c33;
1171: douta=16'h5b2f;
1172: douta=16'h9c2e;
1173: douta=16'h31ea;
1174: douta=16'h1906;
1175: douta=16'h10e4;
1176: douta=16'h10e4;
1177: douta=16'h0000;
1178: douta=16'h940d;
1179: douta=16'h0861;
1180: douta=16'h8c0d;
1181: douta=16'h8bef;
1182: douta=16'h8d39;
1183: douta=16'h8d38;
1184: douta=16'h7c96;
1185: douta=16'h9538;
1186: douta=16'h8d58;
1187: douta=16'h9579;
1188: douta=16'ha5ba;
1189: douta=16'h7cb7;
1190: douta=16'h959a;
1191: douta=16'ha5ba;
1192: douta=16'h9579;
1193: douta=16'h2926;
1194: douta=16'h9559;
1195: douta=16'h6c35;
1196: douta=16'h84d7;
1197: douta=16'h7c13;
1198: douta=16'h8cb6;
1199: douta=16'h7497;
1200: douta=16'h7476;
1201: douta=16'h31c8;
1202: douta=16'h7d3a;
1203: douta=16'h6457;
1204: douta=16'h7cd9;
1205: douta=16'h7cd9;
1206: douta=16'h74fa;
1207: douta=16'h853a;
1208: douta=16'h6c36;
1209: douta=16'h8d7a;
1210: douta=16'h6c77;
1211: douta=16'h7cb8;
1212: douta=16'h6391;
1213: douta=16'h9d58;
1214: douta=16'h73f3;
1215: douta=16'h5351;
1216: douta=16'h2250;
1217: douta=16'h32d1;
1218: douta=16'h5bb4;
1219: douta=16'h7435;
1220: douta=16'h94b5;
1221: douta=16'ha42c;
1222: douta=16'hd570;
1223: douta=16'heed7;
1224: douta=16'hddd2;
1225: douta=16'hc52f;
1226: douta=16'h8b69;
1227: douta=16'hb4ed;
1228: douta=16'he655;
1229: douta=16'heeb6;
1230: douta=16'he654;
1231: douta=16'hbd10;
1232: douta=16'h9c72;
1233: douta=16'h73d1;
1234: douta=16'h4a6b;
1235: douta=16'hcd2e;
1236: douta=16'hb48d;
1237: douta=16'h630e;
1238: douta=16'h322c;
1239: douta=16'h1906;
1240: douta=16'h10a3;
1241: douta=16'h10a4;
1242: douta=16'h29a8;
1243: douta=16'h1926;
1244: douta=16'h8c2e;
1245: douta=16'h31a6;
1246: douta=16'h7cb7;
1247: douta=16'h9559;
1248: douta=16'h8d38;
1249: douta=16'h8d18;
1250: douta=16'h8d58;
1251: douta=16'h9559;
1252: douta=16'h9559;
1253: douta=16'h8518;
1254: douta=16'h9d9a;
1255: douta=16'h8d39;
1256: douta=16'h9d9a;
1257: douta=16'had34;
1258: douta=16'h1106;
1259: douta=16'h9d79;
1260: douta=16'h9d58;
1261: douta=16'h9d16;
1262: douta=16'h6cb8;
1263: douta=16'h7d5c;
1264: douta=16'h322c;
1265: douta=16'h7d3a;
1266: douta=16'h8d5a;
1267: douta=16'h7498;
1268: douta=16'h853a;
1269: douta=16'h8d5a;
1270: douta=16'h855a;
1271: douta=16'h853b;
1272: douta=16'h855a;
1273: douta=16'h7cd9;
1274: douta=16'h7498;
1275: douta=16'h6cda;
1276: douta=16'h7414;
1277: douta=16'h7cb7;
1278: douta=16'h5330;
1279: douta=16'h7c95;
1280: douta=16'h328f;
1281: douta=16'h4374;
1282: douta=16'h84d8;
1283: douta=16'h5b51;
1284: douta=16'h9bca;
1285: douta=16'hc4ed;
1286: douta=16'he633;
1287: douta=16'heeb6;
1288: douta=16'hd5b1;
1289: douta=16'h8308;
1290: douta=16'hbccd;
1291: douta=16'hde12;
1292: douta=16'hee95;
1293: douta=16'he613;
1294: douta=16'hc530;
1295: douta=16'h9431;
1296: douta=16'h630e;
1297: douta=16'h49e8;
1298: douta=16'h9bcb;
1299: douta=16'he654;
1300: douta=16'hc4ee;
1301: douta=16'h7b4d;
1302: douta=16'h6b71;
1303: douta=16'h3a8e;
1304: douta=16'h2168;
1305: douta=16'h10e4;
1306: douta=16'h10a4;
1307: douta=16'h1905;
1308: douta=16'h6b90;
1309: douta=16'h5269;
1310: douta=16'h6b2b;
1311: douta=16'h8d38;
1312: douta=16'h84b7;
1313: douta=16'h8d39;
1314: douta=16'h9558;
1315: douta=16'h7496;
1316: douta=16'h84d7;
1317: douta=16'h8d39;
1318: douta=16'h8d18;
1319: douta=16'h8d18;
1320: douta=16'h84f8;
1321: douta=16'h9559;
1322: douta=16'h9db9;
1323: douta=16'h1989;
1324: douta=16'h10e5;
1325: douta=16'h1905;
1326: douta=16'h834c;
1327: douta=16'h63f4;
1328: douta=16'h853b;
1329: douta=16'h6c37;
1330: douta=16'h7cb8;
1331: douta=16'h8d5a;
1332: douta=16'h8d5b;
1333: douta=16'h95bc;
1334: douta=16'h74b8;
1335: douta=16'h8d7b;
1336: douta=16'h5bf5;
1337: douta=16'h851a;
1338: douta=16'h857b;
1339: douta=16'h63d4;
1340: douta=16'h3965;
1341: douta=16'h6c56;
1342: douta=16'h84b6;
1343: douta=16'h1083;
1344: douta=16'h31ca;
1345: douta=16'h4bb5;
1346: douta=16'h63d4;
1347: douta=16'h6392;
1348: douta=16'hc4ed;
1349: douta=16'hde13;
1350: douta=16'hee95;
1351: douta=16'hd5b0;
1352: douta=16'hbcee;
1353: douta=16'hb4cd;
1354: douta=16'hde33;
1355: douta=16'he675;
1356: douta=16'hee75;
1357: douta=16'hd590;
1358: douta=16'h83d0;
1359: douta=16'h734f;
1360: douta=16'h2925;
1361: douta=16'hcd2f;
1362: douta=16'hee95;
1363: douta=16'hee54;
1364: douta=16'hc4cf;
1365: douta=16'h93ce;
1366: douta=16'h7bf2;
1367: douta=16'h5b91;
1368: douta=16'h29cb;
1369: douta=16'h31eb;
1370: douta=16'h1905;
1371: douta=16'h2147;
1372: douta=16'h18e5;
1373: douta=16'h10e4;
1374: douta=16'h6b6d;
1375: douta=16'h8bed;
1376: douta=16'h7cb7;
1377: douta=16'h84f8;
1378: douta=16'h63f4;
1379: douta=16'h8d38;
1380: douta=16'h8d18;
1381: douta=16'hbe7c;
1382: douta=16'h8d39;
1383: douta=16'h9559;
1384: douta=16'h8d39;
1385: douta=16'h8d18;
1386: douta=16'h957a;
1387: douta=16'h9d9a;
1388: douta=16'h853a;
1389: douta=16'h2188;
1390: douta=16'h8d59;
1391: douta=16'h959a;
1392: douta=16'h8539;
1393: douta=16'h7cf8;
1394: douta=16'h9dbb;
1395: douta=16'h959a;
1396: douta=16'h8d3a;
1397: douta=16'h855a;
1398: douta=16'h7498;
1399: douta=16'h853a;
1400: douta=16'h95bc;
1401: douta=16'h74b8;
1402: douta=16'h32ae;
1403: douta=16'hae1c;
1404: douta=16'h4b33;
1405: douta=16'h0000;
1406: douta=16'h61e4;
1407: douta=16'h0882;
1408: douta=16'h1083;
1409: douta=16'h32b1;
1410: douta=16'h7456;
1411: douta=16'h6372;
1412: douta=16'hbcef;
1413: douta=16'hee76;
1414: douta=16'he613;
1415: douta=16'h7b07;
1416: douta=16'hbcee;
1417: douta=16'hd5d3;
1418: douta=16'hddf3;
1419: douta=16'hee95;
1420: douta=16'hde12;
1421: douta=16'ha46f;
1422: douta=16'h6b2c;
1423: douta=16'h3145;
1424: douta=16'hc4cc;
1425: douta=16'hde33;
1426: douta=16'heeb6;
1427: douta=16'hd572;
1428: douta=16'hac50;
1429: douta=16'h8c31;
1430: douta=16'h8412;
1431: douta=16'h736f;
1432: douta=16'h6a8a;
1433: douta=16'h4ace;
1434: douta=16'h2147;
1435: douta=16'h5b0e;
1436: douta=16'h10e5;
1437: douta=16'h18c4;
1438: douta=16'h0883;
1439: douta=16'h9492;
1440: douta=16'h634d;
1441: douta=16'h8d18;
1442: douta=16'h9579;
1443: douta=16'h9579;
1444: douta=16'h8d18;
1445: douta=16'h84d7;
1446: douta=16'h7c96;
1447: douta=16'h5352;
1448: douta=16'h9dbb;
1449: douta=16'h8518;
1450: douta=16'h8539;
1451: douta=16'h7cf8;
1452: douta=16'h8518;
1453: douta=16'h18a2;
1454: douta=16'h8538;
1455: douta=16'h8518;
1456: douta=16'h9ddb;
1457: douta=16'h95ba;
1458: douta=16'h8d9a;
1459: douta=16'ha5db;
1460: douta=16'h957a;
1461: douta=16'h7cd9;
1462: douta=16'h7497;
1463: douta=16'h957b;
1464: douta=16'h84f9;
1465: douta=16'h10a2;
1466: douta=16'h4060;
1467: douta=16'h84f9;
1468: douta=16'h42f1;
1469: douta=16'h8d7a;
1470: douta=16'h8497;
1471: douta=16'h0020;
1472: douta=16'h3146;
1473: douta=16'h32b0;
1474: douta=16'h3aaf;
1475: douta=16'h42af;
1476: douta=16'ha557;
1477: douta=16'hee75;
1478: douta=16'hc50e;
1479: douta=16'hbd0f;
1480: douta=16'he634;
1481: douta=16'heeb7;
1482: douta=16'hee75;
1483: douta=16'hac2d;
1484: douta=16'hac70;
1485: douta=16'h6b4d;
1486: douta=16'h6206;
1487: douta=16'hcd2e;
1488: douta=16'he654;
1489: douta=16'hde13;
1490: douta=16'hcd52;
1491: douta=16'hb4f2;
1492: douta=16'h9473;
1493: douta=16'h736f;
1494: douta=16'h6b0e;
1495: douta=16'hc46c;
1496: douta=16'hde12;
1497: douta=16'h8c10;
1498: douta=16'h5b91;
1499: douta=16'h324d;
1500: douta=16'h08a4;
1501: douta=16'h18e5;
1502: douta=16'h10e4;
1503: douta=16'h1906;
1504: douta=16'h31ea;
1505: douta=16'h4a6a;
1506: douta=16'h2169;
1507: douta=16'h8d18;
1508: douta=16'h7c96;
1509: douta=16'h84d7;
1510: douta=16'h7c76;
1511: douta=16'h8d18;
1512: douta=16'h8d39;
1513: douta=16'h7cb7;
1514: douta=16'h63b2;
1515: douta=16'h8d7a;
1516: douta=16'h8519;
1517: douta=16'h95bc;
1518: douta=16'h74b8;
1519: douta=16'h957a;
1520: douta=16'h8d19;
1521: douta=16'h957a;
1522: douta=16'ha5db;
1523: douta=16'ha5db;
1524: douta=16'h959a;
1525: douta=16'h959a;
1526: douta=16'ha5dc;
1527: douta=16'h5c38;
1528: douta=16'h5373;
1529: douta=16'h6245;
1530: douta=16'h5331;
1531: douta=16'h10a5;
1532: douta=16'h7c32;
1533: douta=16'h5352;
1534: douta=16'h84d8;
1535: douta=16'h4acd;
1536: douta=16'h3145;
1537: douta=16'h4333;
1538: douta=16'h5bb4;
1539: douta=16'h6c35;
1540: douta=16'h8433;
1541: douta=16'hb5b8;
1542: douta=16'hc530;
1543: douta=16'hde15;
1544: douta=16'heeb6;
1545: douta=16'hd591;
1546: douta=16'hd5b2;
1547: douta=16'h9450;
1548: douta=16'h838e;
1549: douta=16'h3945;
1550: douta=16'hd570;
1551: douta=16'hee74;
1552: douta=16'hf6b6;
1553: douta=16'hcd71;
1554: douta=16'ha491;
1555: douta=16'ha4b4;
1556: douta=16'h7bd1;
1557: douta=16'h4a4a;
1558: douta=16'hc4cc;
1559: douta=16'he654;
1560: douta=16'hddd3;
1561: douta=16'ha491;
1562: douta=16'h7c13;
1563: douta=16'h5bb2;
1564: douta=16'h3a6d;
1565: douta=16'h3aae;
1566: douta=16'h10e5;
1567: douta=16'h10c4;
1568: douta=16'h18e5;
1569: douta=16'h0883;
1570: douta=16'h7412;
1571: douta=16'h52cb;
1572: douta=16'h6391;
1573: douta=16'h8497;
1574: douta=16'h8d18;
1575: douta=16'h8cf7;
1576: douta=16'h84b7;
1577: douta=16'h84d7;
1578: douta=16'h8d39;
1579: douta=16'ha5db;
1580: douta=16'h7c96;
1581: douta=16'h7476;
1582: douta=16'h8519;
1583: douta=16'h8d5a;
1584: douta=16'h8519;
1585: douta=16'h959b;
1586: douta=16'h74b8;
1587: douta=16'h959b;
1588: douta=16'h8d9c;
1589: douta=16'h3b12;
1590: douta=16'h74b9;
1591: douta=16'h3b13;
1592: douta=16'h4395;
1593: douta=16'h732c;
1594: douta=16'h0882;
1595: douta=16'h6436;
1596: douta=16'h5c57;
1597: douta=16'h63b1;
1598: douta=16'hadd7;
1599: douta=16'h1840;
1600: douta=16'h3965;
1601: douta=16'h2a4e;
1602: douta=16'h3ad1;
1603: douta=16'h6c15;
1604: douta=16'h73f3;
1605: douta=16'had77;
1606: douta=16'hee95;
1607: douta=16'heed8;
1608: douta=16'hee96;
1609: douta=16'hde13;
1610: douta=16'h8c10;
1611: douta=16'h7390;
1612: douta=16'h4985;
1613: douta=16'hd570;
1614: douta=16'he633;
1615: douta=16'hde13;
1616: douta=16'hc530;
1617: douta=16'ha4b2;
1618: douta=16'h9472;
1619: douta=16'h7bb0;
1620: douta=16'h7a87;
1621: douta=16'hddd1;
1622: douta=16'hee74;
1623: douta=16'he632;
1624: douta=16'hbd0f;
1625: douta=16'h9451;
1626: douta=16'h8c94;
1627: douta=16'h8475;
1628: douta=16'h63b2;
1629: douta=16'h7b2d;
1630: douta=16'h3a8d;
1631: douta=16'h4acf;
1632: douta=16'h18e5;
1633: douta=16'h10c4;
1634: douta=16'h1926;
1635: douta=16'h1905;
1636: douta=16'h1926;
1637: douta=16'had11;
1638: douta=16'h62eb;
1639: douta=16'h4208;
1640: douta=16'h7476;
1641: douta=16'h8d18;
1642: douta=16'h9559;
1643: douta=16'h8d39;
1644: douta=16'h6c76;
1645: douta=16'h8d39;
1646: douta=16'h84f8;
1647: douta=16'h5371;
1648: douta=16'h8539;
1649: douta=16'h7496;
1650: douta=16'h4310;
1651: douta=16'h62ed;
1652: douta=16'h6248;
1653: douta=16'h4395;
1654: douta=16'h3b33;
1655: douta=16'h4374;
1656: douta=16'h53d6;
1657: douta=16'h5c37;
1658: douta=16'h51c4;
1659: douta=16'h08e5;
1660: douta=16'had10;
1661: douta=16'h3944;
1662: douta=16'h41a5;
1663: douta=16'h49c7;
1664: douta=16'h3945;
1665: douta=16'h4acf;
1666: douta=16'h3ad1;
1667: douta=16'h5373;
1668: douta=16'h4aef;
1669: douta=16'h8411;
1670: douta=16'hb5b7;
1671: douta=16'hee96;
1672: douta=16'he675;
1673: douta=16'hc531;
1674: douta=16'h7b70;
1675: douta=16'h2904;
1676: douta=16'hd570;
1677: douta=16'he655;
1678: douta=16'hee75;
1679: douta=16'ha491;
1680: douta=16'h9432;
1681: douta=16'h7bd1;
1682: douta=16'h736f;
1683: douta=16'ha40a;
1684: douta=16'hee75;
1685: douta=16'hf6b6;
1686: douta=16'hddd2;
1687: douta=16'hb4d1;
1688: douta=16'h9c72;
1689: douta=16'h83f1;
1690: douta=16'h7bb0;
1691: douta=16'h62cd;
1692: douta=16'hddb0;
1693: douta=16'hddb2;
1694: douta=16'h6bd2;
1695: douta=16'h3a8e;
1696: douta=16'h2168;
1697: douta=16'h2168;
1698: douta=16'h18e6;
1699: douta=16'h1084;
1700: douta=16'h1926;
1701: douta=16'h0000;
1702: douta=16'h2126;
1703: douta=16'h7bef;
1704: douta=16'hde77;
1705: douta=16'h2986;
1706: douta=16'ha4d2;
1707: douta=16'h52cb;
1708: douta=16'h5acb;
1709: douta=16'h39c7;
1710: douta=16'h9348;
1711: douta=16'h31c9;
1712: douta=16'h42ae;
1713: douta=16'h42ae;
1714: douta=16'h6370;
1715: douta=16'h5b91;
1716: douta=16'h5b71;
1717: douta=16'h5a48;
1718: douta=16'h4a8d;
1719: douta=16'h3334;
1720: douta=16'h4bd5;
1721: douta=16'h3af1;
1722: douta=16'hb573;
1723: douta=16'h4985;
1724: douta=16'h41a6;
1725: douta=16'h49e7;
1726: douta=16'h41c7;
1727: douta=16'h41a7;
1728: douta=16'h3103;
1729: douta=16'h31a9;
1730: douta=16'h3a2c;
1731: douta=16'h9cb4;
1732: douta=16'hadb9;
1733: douta=16'h94d5;
1734: douta=16'h8431;
1735: douta=16'hde79;
1736: douta=16'hd5f3;
1737: douta=16'h8c11;
1738: douta=16'h28e3;
1739: douta=16'hd5b0;
1740: douta=16'hee75;
1741: douta=16'he654;
1742: douta=16'hc550;
1743: douta=16'h9c92;
1744: douta=16'h632f;
1745: douta=16'h4aae;
1746: douta=16'he590;
1747: douta=16'hee96;
1748: douta=16'heeb6;
1749: douta=16'hcdb3;
1750: douta=16'h9452;
1751: douta=16'h8432;
1752: douta=16'h736e;
1753: douta=16'h732d;
1754: douta=16'hb44b;
1755: douta=16'hcd0e;
1756: douta=16'hcd92;
1757: douta=16'ha492;
1758: douta=16'h7413;
1759: douta=16'h7413;
1760: douta=16'h5bd4;
1761: douta=16'h29cb;
1762: douta=16'h08c5;
1763: douta=16'h1106;
1764: douta=16'h10e5;
1765: douta=16'h10e5;
1766: douta=16'h1927;
1767: douta=16'h1927;
1768: douta=16'h0062;
1769: douta=16'h10e5;
1770: douta=16'h6c14;
1771: douta=16'h1905;
1772: douta=16'hd50d;
1773: douta=16'h4a4a;
1774: douta=16'h2168;
1775: douta=16'h4a8c;
1776: douta=16'h320b;
1777: douta=16'h4b10;
1778: douta=16'h4b0f;
1779: douta=16'h530f;
1780: douta=16'h5372;
1781: douta=16'h42f0;
1782: douta=16'h3a6c;
1783: douta=16'h49c7;
1784: douta=16'h32f2;
1785: douta=16'h4185;
1786: douta=16'h49a6;
1787: douta=16'h4186;
1788: douta=16'h49c7;
1789: douta=16'h39a6;
1790: douta=16'h49e8;
1791: douta=16'h49e7;
1792: douta=16'h5b2e;
1793: douta=16'h2904;
1794: douta=16'h29c9;
1795: douta=16'ha3ed;
1796: douta=16'h9bed;
1797: douta=16'h52cd;
1798: douta=16'h6baf;
1799: douta=16'h6bb0;
1800: douta=16'h636f;
1801: douta=16'hbc8d;
1802: douta=16'hde53;
1803: douta=16'heeb6;
1804: douta=16'he674;
1805: douta=16'hbd11;
1806: douta=16'h9c92;
1807: douta=16'h7b70;
1808: douta=16'h5a6a;
1809: douta=16'he5d0;
1810: douta=16'hf6f7;
1811: douta=16'he613;
1812: douta=16'hacb2;
1813: douta=16'h9452;
1814: douta=16'h83d0;
1815: douta=16'h732d;
1816: douta=16'h51a5;
1817: douta=16'hd58f;
1818: douta=16'he675;
1819: douta=16'hddd2;
1820: douta=16'hb4d2;
1821: douta=16'h9452;
1822: douta=16'h6b4f;
1823: douta=16'h6b91;
1824: douta=16'h5b10;
1825: douta=16'h5aee;
1826: douta=16'h3a4d;
1827: douta=16'h3aae;
1828: douta=16'h29cb;
1829: douta=16'h322d;
1830: douta=16'h1907;
1831: douta=16'h1927;
1832: douta=16'h10e5;
1833: douta=16'h1105;
1834: douta=16'h10e5;
1835: douta=16'h1926;
1836: douta=16'h2988;
1837: douta=16'h0000;
1838: douta=16'h5373;
1839: douta=16'h6b90;
1840: douta=16'h5b0e;
1841: douta=16'h5b70;
1842: douta=16'h5b50;
1843: douta=16'h5330;
1844: douta=16'h29a8;
1845: douta=16'h6268;
1846: douta=16'h4aaf;
1847: douta=16'h6a66;
1848: douta=16'h51e6;
1849: douta=16'h49c8;
1850: douta=16'h49e8;
1851: douta=16'h41a7;
1852: douta=16'h49c7;
1853: douta=16'h49c7;
1854: douta=16'h49e8;
1855: douta=16'h41c7;
1856: douta=16'h4a09;
1857: douta=16'h3124;
1858: douta=16'h29a9;
1859: douta=16'h7b4c;
1860: douta=16'hac4e;
1861: douta=16'h5aed;
1862: douta=16'h636e;
1863: douta=16'h73d0;
1864: douta=16'h636f;
1865: douta=16'h6baf;
1866: douta=16'hf6f6;
1867: douta=16'hde34;
1868: douta=16'hb4d1;
1869: douta=16'h9431;
1870: douta=16'h6b4f;
1871: douta=16'h51e5;
1872: douta=16'hd591;
1873: douta=16'hee95;
1874: douta=16'hd5d3;
1875: douta=16'h9c93;
1876: douta=16'h8c54;
1877: douta=16'h7bf2;
1878: douta=16'h5aef;
1879: douta=16'hcd0e;
1880: douta=16'hd570;
1881: douta=16'hddf3;
1882: douta=16'hcd50;
1883: douta=16'h9411;
1884: douta=16'h838f;
1885: douta=16'h730d;
1886: douta=16'h62cd;
1887: douta=16'h734d;
1888: douta=16'heeb7;
1889: douta=16'ha4b2;
1890: douta=16'h5b50;
1891: douta=16'h5b72;
1892: douta=16'h4acf;
1893: douta=16'h42af;
1894: douta=16'h21aa;
1895: douta=16'h10a5;
1896: douta=16'h29ca;
1897: douta=16'h10e5;
1898: douta=16'h18e5;
1899: douta=16'h1905;
1900: douta=16'h1906;
1901: douta=16'h1905;
1902: douta=16'h18e5;
1903: douta=16'h0884;
1904: douta=16'h3a8d;
1905: douta=16'h5b0e;
1906: douta=16'h4a4a;
1907: douta=16'h7aa8;
1908: douta=16'h29a9;
1909: douta=16'h5b51;
1910: douta=16'h322d;
1911: douta=16'h6a68;
1912: douta=16'h5a49;
1913: douta=16'h5249;
1914: douta=16'h49c7;
1915: douta=16'h41a7;
1916: douta=16'h49e8;
1917: douta=16'h49e7;
1918: douta=16'h41a7;
1919: douta=16'h41a7;
1920: douta=16'h3944;
1921: douta=16'h3124;
1922: douta=16'h29a8;
1923: douta=16'h4a4a;
1924: douta=16'h5aac;
1925: douta=16'h52cd;
1926: douta=16'h636f;
1927: douta=16'h6bd0;
1928: douta=16'h6bcf;
1929: douta=16'h638f;
1930: douta=16'h6bd0;
1931: douta=16'hc531;
1932: douta=16'h8bcf;
1933: douta=16'h7b6f;
1934: douta=16'h9b6a;
1935: douta=16'hee96;
1936: douta=16'heeb7;
1937: douta=16'hd5b3;
1938: douta=16'h9474;
1939: douta=16'h7bd1;
1940: douta=16'h6b2e;
1941: douta=16'h49a7;
1942: douta=16'hee75;
1943: douta=16'hf6d7;
1944: douta=16'he674;
1945: douta=16'ha471;
1946: douta=16'h7baf;
1947: douta=16'h7b6e;
1948: douta=16'h5249;
1949: douta=16'hbc8f;
1950: douta=16'hd5d4;
1951: douta=16'hcdd5;
1952: douta=16'hb535;
1953: douta=16'h9494;
1954: douta=16'h73d1;
1955: douta=16'h5b30;
1956: douta=16'h4ace;
1957: douta=16'hddd3;
1958: douta=16'h5350;
1959: douta=16'h4af0;
1960: douta=16'h29ca;
1961: douta=16'h1927;
1962: douta=16'h42d0;
1963: douta=16'h2147;
1964: douta=16'h2169;
1965: douta=16'h29aa;
1966: douta=16'h10e5;
1967: douta=16'h10e5;
1968: douta=16'h10c4;
1969: douta=16'h10e5;
1970: douta=16'h3a4d;
1971: douta=16'h428e;
1972: douta=16'h7c13;
1973: douta=16'h5330;
1974: douta=16'h73f4;
1975: douta=16'had34;
1976: douta=16'h5249;
1977: douta=16'h49c7;
1978: douta=16'h49c7;
1979: douta=16'h39a6;
1980: douta=16'h4186;
1981: douta=16'h3986;
1982: douta=16'h41a7;
1983: douta=16'h49e8;
1984: douta=16'h3965;
1985: douta=16'h3124;
1986: douta=16'h2187;
1987: douta=16'h3a0a;
1988: douta=16'h422a;
1989: douta=16'h4aac;
1990: douta=16'h6390;
1991: douta=16'h6bd0;
1992: douta=16'h5b2e;
1993: douta=16'h5b6e;
1994: douta=16'h638e;
1995: douta=16'h530c;
1996: douta=16'h4acb;
1997: douta=16'h4a8c;
1998: douta=16'heeb6;
1999: douta=16'heed7;
2000: douta=16'hc573;
2001: douta=16'had14;
2002: douta=16'h8412;
2003: douta=16'h6b2e;
2004: douta=16'h72ca;
2005: douta=16'hddf2;
2006: douta=16'h83d0;
2007: douta=16'h9c91;
2008: douta=16'h83d1;
2009: douta=16'h7b8f;
2010: douta=16'h62ed;
2011: douta=16'h9bec;
2012: douta=16'hf6d7;
2013: douta=16'hde13;
2014: douta=16'h9453;
2015: douta=16'h9452;
2016: douta=16'h9472;
2017: douta=16'h8432;
2018: douta=16'h736e;
2019: douta=16'heeb5;
2020: douta=16'hacd4;
2021: douta=16'h8433;
2022: douta=16'h630e;
2023: douta=16'h4a8d;
2024: douta=16'h29a9;
2025: douta=16'h7bd2;
2026: douta=16'h5b50;
2027: douta=16'h3a4c;
2028: douta=16'h21cb;
2029: douta=16'h3a4d;
2030: douta=16'h320c;
2031: douta=16'h10e5;
2032: douta=16'h10c4;
2033: douta=16'h10e5;
2034: douta=16'h0884;
2035: douta=16'h6bb1;
2036: douta=16'h5b72;
2037: douta=16'h5b72;
2038: douta=16'h4b31;
2039: douta=16'h6c56;
2040: douta=16'hadda;
2041: douta=16'h5227;
2042: douta=16'h49c7;
2043: douta=16'h41a7;
2044: douta=16'h41a7;
2045: douta=16'h4a08;
2046: douta=16'h49e8;
2047: douta=16'h5208;
2048: douta=16'h41c5;
2049: douta=16'h3124;
2050: douta=16'h2168;
2051: douta=16'h29a9;
2052: douta=16'h320b;
2053: douta=16'h3a4b;
2054: douta=16'h5b2f;
2055: douta=16'h4aed;
2056: douta=16'h532e;
2057: douta=16'h5b4e;
2058: douta=16'h638f;
2059: douta=16'h4acc;
2060: douta=16'h530d;
2061: douta=16'h530c;
2062: douta=16'hacb1;
2063: douta=16'hd5f4;
2064: douta=16'ha4d4;
2065: douta=16'h9cd4;
2066: douta=16'h734e;
2067: douta=16'he5d1;
2068: douta=16'heed7;
2069: douta=16'he635;
2070: douta=16'h9cb3;
2071: douta=16'h6bd3;
2072: douta=16'h6b0d;
2073: douta=16'h5a8b;
2074: douta=16'he612;
2075: douta=16'hee96;
2076: douta=16'hb514;
2077: douta=16'hacd4;
2078: douta=16'h8412;
2079: douta=16'h7baf;
2080: douta=16'h93ee;
2081: douta=16'hc553;
2082: douta=16'h9c53;
2083: douta=16'ha4d4;
2084: douta=16'h8432;
2085: douta=16'h734e;
2086: douta=16'h62ac;
2087: douta=16'ha493;
2088: douta=16'h83d1;
2089: douta=16'h630e;
2090: douta=16'h52ad;
2091: douta=16'hacd4;
2092: douta=16'h8452;
2093: douta=16'h4a8d;
2094: douta=16'h3a4d;
2095: douta=16'h5b72;
2096: douta=16'h530f;
2097: douta=16'h29aa;
2098: douta=16'h08c4;
2099: douta=16'h10e6;
2100: douta=16'h6bf3;
2101: douta=16'h7435;
2102: douta=16'h6c56;
2103: douta=16'h7497;
2104: douta=16'h5bd4;
2105: douta=16'h74b8;
2106: douta=16'h959c;
2107: douta=16'h49e7;
2108: douta=16'h5208;
2109: douta=16'h5208;
2110: douta=16'h5208;
2111: douta=16'h5228;
2112: douta=16'hedec;
2113: douta=16'h7bd1;
2114: douta=16'h10a3;
2115: douta=16'h2146;
2116: douta=16'h29ea;
2117: douta=16'h29ea;
2118: douta=16'h4ace;
2119: douta=16'h530e;
2120: douta=16'h3a6b;
2121: douta=16'h530e;
2122: douta=16'h4aed;
2123: douta=16'h4acc;
2124: douta=16'h4aac;
2125: douta=16'h636f;
2126: douta=16'h63d0;
2127: douta=16'h63d0;
2128: douta=16'h7bd0;
2129: douta=16'h6b2d;
2130: douta=16'hbcae;
2131: douta=16'hf759;
2132: douta=16'he675;
2133: douta=16'h9c93;
2134: douta=16'h7bd1;
2135: douta=16'h6b2d;
2136: douta=16'h4a4b;
2137: douta=16'he674;
2138: douta=16'hbd54;
2139: douta=16'h8c94;
2140: douta=16'h632f;
2141: douta=16'h838f;
2142: douta=16'h5a6c;
2143: douta=16'he655;
2144: douta=16'h8453;
2145: douta=16'h6b91;
2146: douta=16'h9430;
2147: douta=16'h6aec;
2148: douta=16'h8c11;
2149: douta=16'h8412;
2150: douta=16'h736f;
2151: douta=16'h7b8f;
2152: douta=16'h6b4e;
2153: douta=16'hcdd4;
2154: douta=16'h8c53;
2155: douta=16'h8c52;
2156: douta=16'h7390;
2157: douta=16'h632e;
2158: douta=16'hd5d5;
2159: douta=16'h9cf5;
2160: douta=16'h6bb2;
2161: douta=16'h3a2c;
2162: douta=16'h2168;
2163: douta=16'h2126;
2164: douta=16'h1905;
2165: douta=16'h8cf6;
2166: douta=16'h8cf8;
2167: douta=16'h7c75;
2168: douta=16'h5bf5;
2169: douta=16'h1926;
2170: douta=16'h21a9;
2171: douta=16'h29c9;
2172: douta=16'h49c7;
2173: douta=16'h5229;
2174: douta=16'h49e8;
2175: douta=16'h49e8;
2176: douta=16'hdd4b;
2177: douta=16'h5164;
2178: douta=16'h83f2;
2179: douta=16'ha410;
2180: douta=16'h21ca;
2181: douta=16'h2189;
2182: douta=16'h3a6d;
2183: douta=16'h42ae;
2184: douta=16'h324b;
2185: douta=16'h3a6b;
2186: douta=16'h3a6b;
2187: douta=16'h4b0e;
2188: douta=16'h4a8c;
2189: douta=16'h530e;
2190: douta=16'h5b6f;
2191: douta=16'h5b6f;
2192: douta=16'h6390;
2193: douta=16'h5b70;
2194: douta=16'hc510;
2195: douta=16'hacb2;
2196: douta=16'h8432;
2197: douta=16'h83d0;
2198: douta=16'h6b0d;
2199: douta=16'h8b29;
2200: douta=16'hde35;
2201: douta=16'h8c74;
2202: douta=16'h8c94;
2203: douta=16'h734e;
2204: douta=16'h8390;
2205: douta=16'hd5b3;
2206: douta=16'hbd55;
2207: douta=16'h8434;
2208: douta=16'h736f;
2209: douta=16'h420a;
2210: douta=16'h7bb0;
2211: douta=16'h732e;
2212: douta=16'h732d;
2213: douta=16'h31c9;
2214: douta=16'hcdb4;
2215: douta=16'h9cb5;
2216: douta=16'h7bd1;
2217: douta=16'h6b0e;
2218: douta=16'h5aed;
2219: douta=16'h62ac;
2220: douta=16'he697;
2221: douta=16'hc5b6;
2222: douta=16'had15;
2223: douta=16'h6b91;
2224: douta=16'h6b91;
2225: douta=16'h4ace;
2226: douta=16'hc574;
2227: douta=16'h18c5;
2228: douta=16'h10c4;
2229: douta=16'h0083;
2230: douta=16'h9d58;
2231: douta=16'h9d58;
2232: douta=16'h5330;
2233: douta=16'h6c14;
2234: douta=16'h6bf3;
2235: douta=16'h6247;
2236: douta=16'h61e4;
2237: douta=16'h5a28;
2238: douta=16'h41a7;
2239: douta=16'h41c7;
2240: douta=16'he56c;
2241: douta=16'h7aa8;
2242: douta=16'hac92;
2243: douta=16'he676;
2244: douta=16'h7c55;
2245: douta=16'h1927;
2246: douta=16'h326d;
2247: douta=16'h3a8d;
2248: douta=16'h3a4c;
2249: douta=16'h3a6c;
2250: douta=16'h3a8c;
2251: douta=16'h3a6b;
2252: douta=16'h636f;
2253: douta=16'h634f;
2254: douta=16'h532e;
2255: douta=16'h534f;
2256: douta=16'h5b4f;
2257: douta=16'h5b6f;
2258: douta=16'h638f;
2259: douta=16'h6bd0;
2260: douta=16'h736e;
2261: douta=16'h72cb;
2262: douta=16'hde55;
2263: douta=16'hc574;
2264: douta=16'h9d17;
2265: douta=16'h7bf2;
2266: douta=16'h7bf1;
2267: douta=16'h4a6c;
2268: douta=16'hd593;
2269: douta=16'h9cd5;
2270: douta=16'h6b90;
2271: douta=16'h3a2b;
2272: douta=16'h93f0;
2273: douta=16'h424c;
2274: douta=16'h6b0c;
2275: douta=16'h522a;
2276: douta=16'hc511;
2277: douta=16'h73d2;
2278: douta=16'h7bf2;
2279: douta=16'h3a6d;
2280: douta=16'h6b4e;
2281: douta=16'hd5d4;
2282: douta=16'hde15;
2283: douta=16'h8c51;
2284: douta=16'h9c93;
2285: douta=16'h9474;
2286: douta=16'h83f2;
2287: douta=16'h6b90;
2288: douta=16'h6aeb;
2289: douta=16'hde34;
2290: douta=16'h7c13;
2291: douta=16'h4aef;
2292: douta=16'h29ca;
2293: douta=16'h2988;
2294: douta=16'h9d59;
2295: douta=16'h2904;
2296: douta=16'h7a44;
2297: douta=16'h7245;
2298: douta=16'h6a24;
2299: douta=16'h6205;
2300: douta=16'h61e5;
2301: douta=16'h51c6;
2302: douta=16'h5208;
2303: douta=16'h41c8;
2304: douta=16'he54b;
2305: douta=16'h92c8;
2306: douta=16'hcd92;
2307: douta=16'hddf6;
2308: douta=16'h84b7;
2309: douta=16'h8496;
2310: douta=16'h326d;
2311: douta=16'h3aae;
2312: douta=16'h3a8d;
2313: douta=16'h29ea;
2314: douta=16'h10a3;
2315: douta=16'h2967;
2316: douta=16'h422a;
2317: douta=16'h39ea;
2318: douta=16'h2146;
2319: douta=16'h10e5;
2320: douta=16'h42ee;
2321: douta=16'h52ed;
2322: douta=16'h5b0e;
2323: douta=16'h638f;
2324: douta=16'h6bb0;
2325: douta=16'h6bb0;
2326: douta=16'h638f;
2327: douta=16'h9cb3;
2328: douta=16'h9493;
2329: douta=16'h7bf1;
2330: douta=16'h93ee;
2331: douta=16'hacf5;
2332: douta=16'h8c95;
2333: douta=16'h7b90;
2334: douta=16'h62cc;
2335: douta=16'hacd3;
2336: douta=16'h6b4f;
2337: douta=16'h2988;
2338: douta=16'h2968;
2339: douta=16'hbd13;
2340: douta=16'h6370;
2341: douta=16'h6b2f;
2342: douta=16'h736f;
2343: douta=16'hd5f4;
2344: douta=16'hcdf7;
2345: douta=16'hc5b6;
2346: douta=16'ha515;
2347: douta=16'h9472;
2348: douta=16'h8432;
2349: douta=16'h62ee;
2350: douta=16'ha46f;
2351: douta=16'he634;
2352: douta=16'hde34;
2353: douta=16'had14;
2354: douta=16'h7c34;
2355: douta=16'h63f4;
2356: douta=16'h42ae;
2357: douta=16'h7c54;
2358: douta=16'h18e5;
2359: douta=16'h7aa5;
2360: douta=16'h7a65;
2361: douta=16'h7224;
2362: douta=16'h61c4;
2363: douta=16'h59e5;
2364: douta=16'h8c51;
2365: douta=16'h9d13;
2366: douta=16'h7b8d;
2367: douta=16'h4a27;
2368: douta=16'hd484;
2369: douta=16'hff3a;
2370: douta=16'hff3a;
2371: douta=16'h8433;
2372: douta=16'h6b2f;
2373: douta=16'h9518;
2374: douta=16'h21ca;
2375: douta=16'h3a6d;
2376: douta=16'h42af;
2377: douta=16'h1947;
2378: douta=16'h1927;
2379: douta=16'h31c9;
2380: douta=16'h426c;
2381: douta=16'h4a8c;
2382: douta=16'h424c;
2383: douta=16'h31c9;
2384: douta=16'h29a8;
2385: douta=16'h320a;
2386: douta=16'h52cd;
2387: douta=16'h5b2e;
2388: douta=16'h5b2e;
2389: douta=16'h636f;
2390: douta=16'h73f0;
2391: douta=16'h634d;
2392: douta=16'h6b6e;
2393: douta=16'h7baf;
2394: douta=16'h736d;
2395: douta=16'h8bcf;
2396: douta=16'h736d;
2397: douta=16'h836d;
2398: douta=16'h8c32;
2399: douta=16'h732d;
2400: douta=16'h6acb;
2401: douta=16'hc574;
2402: douta=16'h9495;
2403: douta=16'h7bf1;
2404: douta=16'h734f;
2405: douta=16'hb535;
2406: douta=16'hd5f6;
2407: douta=16'had56;
2408: douta=16'h7bf1;
2409: douta=16'h7bf2;
2410: douta=16'h7c12;
2411: douta=16'h524a;
2412: douta=16'hddf4;
2413: douta=16'hde35;
2414: douta=16'hacd1;
2415: douta=16'hacb4;
2416: douta=16'h9cb4;
2417: douta=16'h8453;
2418: douta=16'h73b2;
2419: douta=16'h5b51;
2420: douta=16'h6b2d;
2421: douta=16'h52cc;
2422: douta=16'h1926;
2423: douta=16'h83cc;
2424: douta=16'h82c7;
2425: douta=16'h61c4;
2426: douta=16'h61e5;
2427: douta=16'h59e5;
2428: douta=16'h51a5;
2429: douta=16'h4985;
2430: douta=16'h49a5;
2431: douta=16'h4186;
2432: douta=16'hf6b7;
2433: douta=16'hff3a;
2434: douta=16'hf718;
2435: douta=16'h8c94;
2436: douta=16'h8c74;
2437: douta=16'h31e9;
2438: douta=16'h18e5;
2439: douta=16'h1926;
2440: douta=16'h1967;
2441: douta=16'h1148;
2442: douta=16'h1906;
2443: douta=16'h18e5;
2444: douta=16'h2148;
2445: douta=16'h5b30;
2446: douta=16'h2988;
2447: douta=16'h31a9;
2448: douta=16'h31c9;
2449: douta=16'h29ea;
2450: douta=16'h4aad;
2451: douta=16'h52ed;
2452: douta=16'h634e;
2453: douta=16'h5b2d;
2454: douta=16'h52ab;
2455: douta=16'h528a;
2456: douta=16'h5acb;
2457: douta=16'h630c;
2458: douta=16'h62cb;
2459: douta=16'h734d;
2460: douta=16'h7baf;
2461: douta=16'h83cf;
2462: douta=16'h8431;
2463: douta=16'hb533;
2464: douta=16'hccaa;
2465: douta=16'hc468;
2466: douta=16'h7b6f;
2467: douta=16'h7b4d;
2468: douta=16'he697;
2469: douta=16'hbd96;
2470: douta=16'h94d5;
2471: douta=16'h736f;
2472: douta=16'h6b2e;
2473: douta=16'h8bee;
2474: douta=16'he656;
2475: douta=16'hddf5;
2476: douta=16'hbd95;
2477: douta=16'h8c74;
2478: douta=16'h7bd1;
2479: douta=16'h6b4f;
2480: douta=16'h5acc;
2481: douta=16'h5a8a;
2482: douta=16'h942e;
2483: douta=16'hd5d3;
2484: douta=16'hacf4;
2485: douta=16'h5b30;
2486: douta=16'h31ea;
2487: douta=16'h1906;
2488: douta=16'h8286;
2489: douta=16'h6a04;
2490: douta=16'h61e4;
2491: douta=16'h59c5;
2492: douta=16'h51c5;
2493: douta=16'h51c5;
2494: douta=16'h49a6;
2495: douta=16'h41a6;
2496: douta=16'hf6f9;
2497: douta=16'hf6f9;
2498: douta=16'hc5b6;
2499: douta=16'h94b5;
2500: douta=16'ha517;
2501: douta=16'h7435;
2502: douta=16'h8497;
2503: douta=16'h1105;
2504: douta=16'h1947;
2505: douta=16'h1927;
2506: douta=16'h1926;
2507: douta=16'h1082;
2508: douta=16'h2168;
2509: douta=16'h18e4;
2510: douta=16'h18a1;
2511: douta=16'h0821;
2512: douta=16'h1905;
2513: douta=16'h3a0a;
2514: douta=16'h31e9;
2515: douta=16'h39c8;
2516: douta=16'h3a09;
2517: douta=16'h4a4a;
2518: douta=16'h638e;
2519: douta=16'h8473;
2520: douta=16'h6b8f;
2521: douta=16'hcd70;
2522: douta=16'hcbe3;
2523: douta=16'hc3e2;
2524: douta=16'hcc25;
2525: douta=16'hcc45;
2526: douta=16'hcc45;
2527: douta=16'hcc46;
2528: douta=16'hcc46;
2529: douta=16'hd466;
2530: douta=16'hd466;
2531: douta=16'hd486;
2532: douta=16'h9c51;
2533: douta=16'ha4f5;
2534: douta=16'h73d0;
2535: douta=16'h732e;
2536: douta=16'hbd52;
2537: douta=16'hde15;
2538: douta=16'hb535;
2539: douta=16'h8412;
2540: douta=16'h9494;
2541: douta=16'h630e;
2542: douta=16'h632f;
2543: douta=16'h5228;
2544: douta=16'hc550;
2545: douta=16'he676;
2546: douta=16'he656;
2547: douta=16'hcdb5;
2548: douta=16'h94d5;
2549: douta=16'h6bf3;
2550: douta=16'h4b10;
2551: douta=16'h1106;
2552: douta=16'h10c6;
2553: douta=16'h6a24;
2554: douta=16'h6205;
2555: douta=16'h59c5;
2556: douta=16'h51c6;
2557: douta=16'h49c6;
2558: douta=16'h4985;
2559: douta=16'h4165;
2560: douta=16'hff19;
2561: douta=16'hff19;
2562: douta=16'ha4d5;
2563: douta=16'ha4f5;
2564: douta=16'h9cd5;
2565: douta=16'h7434;
2566: douta=16'h7c76;
2567: douta=16'h73f3;
2568: douta=16'h10c5;
2569: douta=16'h10e5;
2570: douta=16'h10e5;
2571: douta=16'h1906;
2572: douta=16'h18e5;
2573: douta=16'h10e4;
2574: douta=16'h2125;
2575: douta=16'h31ea;
2576: douta=16'h3a2c;
2577: douta=16'h42ce;
2578: douta=16'h51a5;
2579: douta=16'h69e3;
2580: douta=16'h8aa4;
2581: douta=16'h92e4;
2582: douta=16'ha345;
2583: douta=16'hab85;
2584: douta=16'hb384;
2585: douta=16'hbbc5;
2586: douta=16'hc3e5;
2587: douta=16'hc426;
2588: douta=16'hcc25;
2589: douta=16'hcc25;
2590: douta=16'hc3e2;
2591: douta=16'hcca8;
2592: douta=16'heed7;
2593: douta=16'hf7bb;
2594: douta=16'hddaf;
2595: douta=16'hcc22;
2596: douta=16'hd466;
2597: douta=16'hd466;
2598: douta=16'hd5d5;
2599: douta=16'hde35;
2600: douta=16'hbd98;
2601: douta=16'h7bf2;
2602: douta=16'h7b90;
2603: douta=16'h630e;
2604: douta=16'h4a49;
2605: douta=16'hc571;
2606: douta=16'hde56;
2607: douta=16'hde55;
2608: douta=16'hde56;
2609: douta=16'hbd14;
2610: douta=16'h8c93;
2611: douta=16'h7c32;
2612: douta=16'h7c33;
2613: douta=16'h6bf2;
2614: douta=16'h6b91;
2615: douta=16'h428d;
2616: douta=16'h10e5;
2617: douta=16'h7245;
2618: douta=16'h6205;
2619: douta=16'h5a05;
2620: douta=16'h51c6;
2621: douta=16'h49a6;
2622: douta=16'h4185;
2623: douta=16'h4166;
2624: douta=16'hff7b;
2625: douta=16'heeb9;
2626: douta=16'ha4d5;
2627: douta=16'hb514;
2628: douta=16'h73f3;
2629: douta=16'h7c55;
2630: douta=16'h8476;
2631: douta=16'h322a;
2632: douta=16'h0883;
2633: douta=16'h10a5;
2634: douta=16'h2188;
2635: douta=16'h29ca;
2636: douta=16'h20e4;
2637: douta=16'h28a1;
2638: douta=16'h4143;
2639: douta=16'h3102;
2640: douta=16'h59c4;
2641: douta=16'h61e4;
2642: douta=16'h7224;
2643: douta=16'h7a64;
2644: douta=16'h8aa4;
2645: douta=16'h9b05;
2646: douta=16'ha345;
2647: douta=16'hab22;
2648: douta=16'hbc48;
2649: douta=16'hef18;
2650: douta=16'hef17;
2651: douta=16'hcce9;
2652: douta=16'hc3e2;
2653: douta=16'hcc25;
2654: douta=16'hcc66;
2655: douta=16'hcc45;
2656: douta=16'hcc66;
2657: douta=16'hd466;
2658: douta=16'hd466;
2659: douta=16'hd466;
2660: douta=16'hd467;
2661: douta=16'hd467;
2662: douta=16'hd465;
2663: douta=16'h9453;
2664: douta=16'h83f1;
2665: douta=16'h7391;
2666: douta=16'h49e7;
2667: douta=16'hc592;
2668: douta=16'he6b7;
2669: douta=16'he656;
2670: douta=16'hcd95;
2671: douta=16'h9cd5;
2672: douta=16'h8c53;
2673: douta=16'h7bf1;
2674: douta=16'h8411;
2675: douta=16'h630c;
2676: douta=16'h940d;
2677: douta=16'ha46e;
2678: douta=16'hb4d1;
2679: douta=16'h31a8;
2680: douta=16'h10e6;
2681: douta=16'h18e5;
2682: douta=16'h6205;
2683: douta=16'h59e6;
2684: douta=16'h49a5;
2685: douta=16'h49a6;
2686: douta=16'h4185;
2687: douta=16'h4166;
2688: douta=16'hffbc;
2689: douta=16'hd5b3;
2690: douta=16'hb556;
2691: douta=16'hb555;
2692: douta=16'h8454;
2693: douta=16'h7c34;
2694: douta=16'h8454;
2695: douta=16'h18c3;
2696: douta=16'h1861;
2697: douta=16'h1883;
2698: douta=16'h20a2;
2699: douta=16'h28c3;
2700: douta=16'h2904;
2701: douta=16'h3903;
2702: douta=16'h4964;
2703: douta=16'h5984;
2704: douta=16'h5983;
2705: douta=16'h8329;
2706: douta=16'hbd91;
2707: douta=16'hb4ee;
2708: douta=16'h9306;
2709: douta=16'h9282;
2710: douta=16'hab85;
2711: douta=16'hb3a5;
2712: douta=16'hc405;
2713: douta=16'hc405;
2714: douta=16'hc425;
2715: douta=16'hc425;
2716: douta=16'hcc25;
2717: douta=16'hcc26;
2718: douta=16'hcc46;
2719: douta=16'hcc46;
2720: douta=16'hcc66;
2721: douta=16'hcc66;
2722: douta=16'hcc66;
2723: douta=16'hd467;
2724: douta=16'hd466;
2725: douta=16'hd467;
2726: douta=16'hd467;
2727: douta=16'hd487;
2728: douta=16'h9c4e;
2729: douta=16'hc573;
2730: douta=16'hde16;
2731: douta=16'hcdd5;
2732: douta=16'ha4d3;
2733: douta=16'h9494;
2734: douta=16'h7bf2;
2735: douta=16'h73d1;
2736: douta=16'h4a28;
2737: douta=16'h83cd;
2738: douta=16'hb4f1;
2739: douta=16'h83ac;
2740: douta=16'hd5d4;
2741: douta=16'h9c6f;
2742: douta=16'hacd2;
2743: douta=16'h4ace;
2744: douta=16'h18e5;
2745: douta=16'h1926;
2746: douta=16'h59e6;
2747: douta=16'h51c5;
2748: douta=16'h49a5;
2749: douta=16'h4986;
2750: douta=16'h4186;
2751: douta=16'h3986;
2752: douta=16'hfffe;
2753: douta=16'hb555;
2754: douta=16'hbd75;
2755: douta=16'ha516;
2756: douta=16'h8c75;
2757: douta=16'h8475;
2758: douta=16'h324b;
2759: douta=16'h18a2;
2760: douta=16'h1040;
2761: douta=16'h20c3;
2762: douta=16'h39a6;
2763: douta=16'h5269;
2764: douta=16'h2967;
2765: douta=16'h3902;
2766: douta=16'h4963;
2767: douta=16'h6aea;
2768: douta=16'h61e4;
2769: douta=16'h7224;
2770: douta=16'h7244;
2771: douta=16'h7a63;
2772: douta=16'h8ac5;
2773: douta=16'h9b05;
2774: douta=16'hab65;
2775: douta=16'hb3a5;
2776: douta=16'hbbc5;
2777: douta=16'hc405;
2778: douta=16'hc405;
2779: douta=16'hc405;
2780: douta=16'hc425;
2781: douta=16'hcc26;
2782: douta=16'hcc46;
2783: douta=16'hcc46;
2784: douta=16'hd467;
2785: douta=16'hd466;
2786: douta=16'hd466;
2787: douta=16'hd466;
2788: douta=16'hd467;
2789: douta=16'hd467;
2790: douta=16'hd467;
2791: douta=16'hd487;
2792: douta=16'h942f;
2793: douta=16'ha4d3;
2794: douta=16'h94b5;
2795: douta=16'h7bf2;
2796: douta=16'h6bb1;
2797: douta=16'h5acb;
2798: douta=16'h5a8a;
2799: douta=16'hb4d0;
2800: douta=16'hbd10;
2801: douta=16'hbd52;
2802: douta=16'hd635;
2803: douta=16'hde35;
2804: douta=16'hc573;
2805: douta=16'h9cb4;
2806: douta=16'h8c93;
2807: douta=16'h6b6f;
2808: douta=16'h424b;
2809: douta=16'h3189;
2810: douta=16'h1905;
2811: douta=16'h51c5;
2812: douta=16'h49a6;
2813: douta=16'h49a6;
2814: douta=16'h4166;
2815: douta=16'h3986;
2816: douta=16'hde77;
2817: douta=16'ha4b4;
2818: douta=16'hc595;
2819: douta=16'h8c74;
2820: douta=16'h8454;
2821: douta=16'h8454;
2822: douta=16'h18c3;
2823: douta=16'h1082;
2824: douta=16'h1882;
2825: douta=16'h20a2;
2826: douta=16'h20a2;
2827: douta=16'h28e2;
2828: douta=16'h2988;
2829: douta=16'h4143;
2830: douta=16'h51a4;
2831: douta=16'h9d13;
2832: douta=16'h7224;
2833: douta=16'h7244;
2834: douta=16'h7224;
2835: douta=16'h8284;
2836: douta=16'h92c4;
2837: douta=16'ha325;
2838: douta=16'hab85;
2839: douta=16'hb385;
2840: douta=16'hbbe5;
2841: douta=16'hbc06;
2842: douta=16'hc426;
2843: douta=16'hc425;
2844: douta=16'hc425;
2845: douta=16'hcc46;
2846: douta=16'hcc47;
2847: douta=16'hd466;
2848: douta=16'hd467;
2849: douta=16'hd467;
2850: douta=16'hd466;
2851: douta=16'hd467;
2852: douta=16'hd467;
2853: douta=16'hd467;
2854: douta=16'hd467;
2855: douta=16'hd487;
2856: douta=16'hbccd;
2857: douta=16'h9410;
2858: douta=16'h734e;
2859: douta=16'h49e6;
2860: douta=16'hd614;
2861: douta=16'hbd30;
2862: douta=16'hbd52;
2863: douta=16'he676;
2864: douta=16'hde35;
2865: douta=16'ha4d3;
2866: douta=16'hb534;
2867: douta=16'hb514;
2868: douta=16'h8432;
2869: douta=16'h73b1;
2870: douta=16'h5a69;
2871: douta=16'h62ca;
2872: douta=16'h5b50;
2873: douta=16'h736f;
2874: douta=16'h2126;
2875: douta=16'h51e6;
2876: douta=16'h49a6;
2877: douta=16'h4186;
2878: douta=16'h3966;
2879: douta=16'h4166;
2880: douta=16'he698;
2881: douta=16'had15;
2882: douta=16'hbd55;
2883: douta=16'h9494;
2884: douta=16'h8434;
2885: douta=16'h73f2;
2886: douta=16'h20c3;
2887: douta=16'h1882;
2888: douta=16'h18a2;
2889: douta=16'h20a2;
2890: douta=16'h20c2;
2891: douta=16'h28e2;
2892: douta=16'h18e5;
2893: douta=16'h4963;
2894: douta=16'h59a4;
2895: douta=16'h8bec;
2896: douta=16'h59a4;
2897: douta=16'h7a64;
2898: douta=16'h7a44;
2899: douta=16'h82a5;
2900: douta=16'h9304;
2901: douta=16'ha325;
2902: douta=16'hab85;
2903: douta=16'hb3a6;
2904: douta=16'hbbe6;
2905: douta=16'hbc06;
2906: douta=16'hc406;
2907: douta=16'hcc47;
2908: douta=16'hcc46;
2909: douta=16'hcc47;
2910: douta=16'hcc46;
2911: douta=16'hcc46;
2912: douta=16'hd467;
2913: douta=16'hcc67;
2914: douta=16'hd467;
2915: douta=16'hd467;
2916: douta=16'hd467;
2917: douta=16'hd487;
2918: douta=16'hd467;
2919: douta=16'hd487;
2920: douta=16'hbcce;
2921: douta=16'hd486;
2922: douta=16'h9c2e;
2923: douta=16'hbd73;
2924: douta=16'hcdd6;
2925: douta=16'hd5f4;
2926: douta=16'hbd33;
2927: douta=16'hb513;
2928: douta=16'h9cb4;
2929: douta=16'h8c73;
2930: douta=16'h7bb0;
2931: douta=16'h51e6;
2932: douta=16'h5226;
2933: douta=16'h62c9;
2934: douta=16'h83cd;
2935: douta=16'h9c4f;
2936: douta=16'h2967;
2937: douta=16'h0883;
2938: douta=16'h2126;
2939: douta=16'h51c6;
2940: douta=16'h4986;
2941: douta=16'h4185;
2942: douta=16'h4186;
2943: douta=16'h4186;
2944: douta=16'hde37;
2945: douta=16'hb514;
2946: douta=16'h9494;
2947: douta=16'h94b5;
2948: douta=16'h8c95;
2949: douta=16'h20c3;
2950: douta=16'h20c3;
2951: douta=16'h1882;
2952: douta=16'h2082;
2953: douta=16'h2082;
2954: douta=16'h28e2;
2955: douta=16'h30e3;
2956: douta=16'h28e4;
2957: douta=16'h4963;
2958: douta=16'h59a4;
2959: douta=16'h61a3;
2960: douta=16'h51a4;
2961: douta=16'h7a64;
2962: douta=16'h7a84;
2963: douta=16'h8ac5;
2964: douta=16'h9305;
2965: douta=16'ha345;
2966: douta=16'hb3a5;
2967: douta=16'hbbc5;
2968: douta=16'hbbe6;
2969: douta=16'hc406;
2970: douta=16'hc426;
2971: douta=16'hcc26;
2972: douta=16'hcc46;
2973: douta=16'hcc46;
2974: douta=16'hcc46;
2975: douta=16'hcc47;
2976: douta=16'hcc46;
2977: douta=16'hd467;
2978: douta=16'hcc67;
2979: douta=16'hd468;
2980: douta=16'hd467;
2981: douta=16'hd467;
2982: douta=16'hd487;
2983: douta=16'hd488;
2984: douta=16'hb4ce;
2985: douta=16'hd487;
2986: douta=16'ha4b1;
2987: douta=16'hcdf5;
2988: douta=16'hbd96;
2989: douta=16'h9493;
2990: douta=16'h83f1;
2991: douta=16'h83f0;
2992: douta=16'h2903;
2993: douta=16'h62ca;
2994: douta=16'h730a;
2995: douta=16'h8c0e;
2996: douta=16'h9c6f;
2997: douta=16'hc572;
2998: douta=16'hd5d4;
2999: douta=16'hacd2;
3000: douta=16'h632e;
3001: douta=16'h426c;
3002: douta=16'h1905;
3003: douta=16'h10e5;
3004: douta=16'h632c;
3005: douta=16'h5228;
3006: douta=16'h4985;
3007: douta=16'h5185;
3008: douta=16'hb535;
3009: douta=16'hc595;
3010: douta=16'h9474;
3011: douta=16'h9495;
3012: douta=16'h9d59;
3013: douta=16'h20a3;
3014: douta=16'h20c3;
3015: douta=16'h20a2;
3016: douta=16'h20a2;
3017: douta=16'h20c2;
3018: douta=16'h28e3;
3019: douta=16'h3103;
3020: douta=16'h4963;
3021: douta=16'h5184;
3022: douta=16'h61e4;
3023: douta=16'h6a24;
3024: douta=16'h6204;
3025: douta=16'h7a84;
3026: douta=16'h8285;
3027: douta=16'h8ac4;
3028: douta=16'h9325;
3029: douta=16'ha345;
3030: douta=16'hb3a6;
3031: douta=16'hbbc6;
3032: douta=16'hbbe5;
3033: douta=16'hc405;
3034: douta=16'hc426;
3035: douta=16'hcc46;
3036: douta=16'hcc46;
3037: douta=16'hcc47;
3038: douta=16'hcc46;
3039: douta=16'hcc67;
3040: douta=16'hd467;
3041: douta=16'hd467;
3042: douta=16'hd467;
3043: douta=16'hd487;
3044: douta=16'hd467;
3045: douta=16'hd467;
3046: douta=16'hd487;
3047: douta=16'hd488;
3048: douta=16'haccd;
3049: douta=16'hcc68;
3050: douta=16'hc468;
3051: douta=16'h83f1;
3052: douta=16'h738f;
3053: douta=16'h49e6;
3054: douta=16'h5a68;
3055: douta=16'h6b0a;
3056: douta=16'h83cd;
3057: douta=16'h942f;
3058: douta=16'hb4f0;
3059: douta=16'hd5d3;
3060: douta=16'hd615;
3061: douta=16'hd5b3;
3062: douta=16'hb4f3;
3063: douta=16'ha4b3;
3064: douta=16'h8c93;
3065: douta=16'h422a;
3066: douta=16'h1927;
3067: douta=16'h18c5;
3068: douta=16'h59e6;
3069: douta=16'h59e6;
3070: douta=16'h59e6;
3071: douta=16'h59e6;
3072: douta=16'had15;
3073: douta=16'hbd55;
3074: douta=16'ha4f5;
3075: douta=16'h8453;
3076: douta=16'h20c3;
3077: douta=16'h20c3;
3078: douta=16'h20c3;
3079: douta=16'h20a2;
3080: douta=16'h20a2;
3081: douta=16'h28c2;
3082: douta=16'h30e2;
3083: douta=16'h3903;
3084: douta=16'h4964;
3085: douta=16'h59a4;
3086: douta=16'h61c3;
3087: douta=16'h7224;
3088: douta=16'h7a44;
3089: douta=16'h7aa5;
3090: douta=16'h8285;
3091: douta=16'h8ac5;
3092: douta=16'h9b25;
3093: douta=16'hab66;
3094: douta=16'hb3c6;
3095: douta=16'hbbe6;
3096: douta=16'hc405;
3097: douta=16'hc406;
3098: douta=16'hc426;
3099: douta=16'hcc26;
3100: douta=16'hcc47;
3101: douta=16'hcc47;
3102: douta=16'hcc68;
3103: douta=16'hcc67;
3104: douta=16'hcc87;
3105: douta=16'hd468;
3106: douta=16'hcc67;
3107: douta=16'hd487;
3108: douta=16'hcc45;
3109: douta=16'hcc25;
3110: douta=16'hd52e;
3111: douta=16'he6b6;
3112: douta=16'hf79b;
3113: douta=16'hf799;
3114: douta=16'he612;
3115: douta=16'h7b6c;
3116: douta=16'h7b6c;
3117: douta=16'h944f;
3118: douta=16'hacaf;
3119: douta=16'hde35;
3120: douta=16'hd5f4;
3121: douta=16'hc5d4;
3122: douta=16'hd5b4;
3123: douta=16'h9453;
3124: douta=16'h7bf1;
3125: douta=16'h7bd1;
3126: douta=16'h49e7;
3127: douta=16'h3144;
3128: douta=16'h6aea;
3129: douta=16'h52cd;
3130: douta=16'h6b4f;
3131: douta=16'h2127;
3132: douta=16'h6206;
3133: douta=16'h61e6;
3134: douta=16'h59a5;
3135: douta=16'h7b4b;
3136: douta=16'hcdb6;
3137: douta=16'h94b4;
3138: douta=16'h94d5;
3139: douta=16'h9d17;
3140: douta=16'h20e3;
3141: douta=16'h20e3;
3142: douta=16'h20c3;
3143: douta=16'h20a2;
3144: douta=16'h20a2;
3145: douta=16'h28e2;
3146: douta=16'h30e3;
3147: douta=16'h4209;
3148: douta=16'h51a4;
3149: douta=16'h59a4;
3150: douta=16'h6ac9;
3151: douta=16'h7244;
3152: douta=16'h7a64;
3153: douta=16'h8285;
3154: douta=16'h8ac5;
3155: douta=16'h8ac5;
3156: douta=16'ha326;
3157: douta=16'haba6;
3158: douta=16'hb3c6;
3159: douta=16'hbbe6;
3160: douta=16'hbc05;
3161: douta=16'hc426;
3162: douta=16'hc425;
3163: douta=16'hc3e3;
3164: douta=16'hc447;
3165: douta=16'hddb0;
3166: douta=16'hf77b;
3167: douta=16'hffdc;
3168: douta=16'he694;
3169: douta=16'hd52b;
3170: douta=16'hcc45;
3171: douta=16'hcc47;
3172: douta=16'hd467;
3173: douta=16'hd488;
3174: douta=16'hd488;
3175: douta=16'hcc88;
3176: douta=16'hcc88;
3177: douta=16'hcc88;
3178: douta=16'hcc68;
3179: douta=16'h9c70;
3180: douta=16'ha4b0;
3181: douta=16'hcd94;
3182: douta=16'hd5f5;
3183: douta=16'hacf4;
3184: douta=16'h8c74;
3185: douta=16'h8433;
3186: douta=16'h4a6a;
3187: douta=16'h2923;
3188: douta=16'h5227;
3189: douta=16'h6ac9;
3190: douta=16'h7b4b;
3191: douta=16'ha46f;
3192: douta=16'ha46f;
3193: douta=16'h3a2b;
3194: douta=16'h0882;
3195: douta=16'h10e5;
3196: douta=16'h1948;
3197: douta=16'h7286;
3198: douta=16'h7a87;
3199: douta=16'h7a87;
3200: douta=16'hc5b5;
3201: douta=16'ha557;
3202: douta=16'h94d5;
3203: douta=16'h1060;
3204: douta=16'h20e3;
3205: douta=16'h20c3;
3206: douta=16'h1882;
3207: douta=16'h20a2;
3208: douta=16'h20c2;
3209: douta=16'h28e2;
3210: douta=16'h3103;
3211: douta=16'h424a;
3212: douta=16'h51a4;
3213: douta=16'h59c4;
3214: douta=16'hb594;
3215: douta=16'h7244;
3216: douta=16'h7a85;
3217: douta=16'h8244;
3218: douta=16'h82c6;
3219: douta=16'hb4af;
3220: douta=16'hde96;
3221: douta=16'hf779;
3222: douta=16'hde32;
3223: douta=16'hc4ca;
3224: douta=16'hbbe5;
3225: douta=16'hc3e5;
3226: douta=16'hc427;
3227: douta=16'hcc47;
3228: douta=16'hcc47;
3229: douta=16'hcc47;
3230: douta=16'hcc48;
3231: douta=16'hcc68;
3232: douta=16'hcc68;
3233: douta=16'hcc68;
3234: douta=16'hd488;
3235: douta=16'hd488;
3236: douta=16'hd488;
3237: douta=16'hcc88;
3238: douta=16'hd488;
3239: douta=16'hd488;
3240: douta=16'hcc68;
3241: douta=16'hd488;
3242: douta=16'hcc25;
3243: douta=16'hccec;
3244: douta=16'hacd2;
3245: douta=16'h9cb4;
3246: douta=16'h7bf2;
3247: douta=16'h3944;
3248: douta=16'h72e9;
3249: douta=16'h8bcd;
3250: douta=16'h9c6f;
3251: douta=16'h730b;
3252: douta=16'hbd52;
3253: douta=16'hd5b3;
3254: douta=16'hd5b3;
3255: douta=16'hc532;
3256: douta=16'hac91;
3257: douta=16'h8c10;
3258: douta=16'h3a2a;
3259: douta=16'h1906;
3260: douta=16'h1128;
3261: douta=16'h8ac7;
3262: douta=16'h8ac7;
3263: douta=16'h8ae7;
3264: douta=16'hbd95;
3265: douta=16'h9cf5;
3266: douta=16'h8433;
3267: douta=16'h20c3;
3268: douta=16'h426b;
3269: douta=16'h20a2;
3270: douta=16'h20a2;
3271: douta=16'h1861;
3272: douta=16'h2082;
3273: douta=16'h3965;
3274: douta=16'h62c9;
3275: douta=16'h1906;
3276: douta=16'h944e;
3277: douta=16'h7b29;
3278: douta=16'h7224;
3279: douta=16'h7203;
3280: douta=16'h8285;
3281: douta=16'h51a4;
3282: douta=16'h92e5;
3283: douta=16'h9306;
3284: douta=16'ha366;
3285: douta=16'hb3a6;
3286: douta=16'hbbe7;
3287: douta=16'hbbe6;
3288: douta=16'hc407;
3289: douta=16'hc426;
3290: douta=16'hcc47;
3291: douta=16'hcc47;
3292: douta=16'hcc67;
3293: douta=16'hcc48;
3294: douta=16'hcc67;
3295: douta=16'hcc25;
3296: douta=16'hcc68;
3297: douta=16'hdd8f;
3298: douta=16'heef8;
3299: douta=16'hffdc;
3300: douta=16'hf738;
3301: douta=16'hddcf;
3302: douta=16'hcca9;
3303: douta=16'hcc26;
3304: douta=16'had11;
3305: douta=16'hd4a9;
3306: douta=16'hcc88;
3307: douta=16'hcc68;
3308: douta=16'h62aa;
3309: douta=16'h730a;
3310: douta=16'h8c0e;
3311: douta=16'hacaf;
3312: douta=16'hcd73;
3313: douta=16'h8bad;
3314: douta=16'hacb3;
3315: douta=16'h7390;
3316: douta=16'h8c32;
3317: douta=16'h7390;
3318: douta=16'h738f;
3319: douta=16'h6b4f;
3320: douta=16'h73b1;
3321: douta=16'h6b70;
3322: douta=16'h6370;
3323: douta=16'h3a2a;
3324: douta=16'hffff;
3325: douta=16'h9b49;
3326: douta=16'h9328;
3327: douta=16'h9328;
3328: douta=16'h9494;
3329: douta=16'ha4f5;
3330: douta=16'h31c7;
3331: douta=16'h28e3;
3332: douta=16'h20e3;
3333: douta=16'h20e3;
3334: douta=16'h20a2;
3335: douta=16'h20a2;
3336: douta=16'h28e3;
3337: douta=16'h3123;
3338: douta=16'h4144;
3339: douta=16'h18a5;
3340: douta=16'h61e4;
3341: douta=16'h6a04;
3342: douta=16'h7a64;
3343: douta=16'h8286;
3344: douta=16'h82a5;
3345: douta=16'h9326;
3346: douta=16'h9306;
3347: douta=16'h9326;
3348: douta=16'ha326;
3349: douta=16'hab64;
3350: douta=16'hc4ac;
3351: douta=16'hde53;
3352: douta=16'hf77a;
3353: douta=16'hef38;
3354: douta=16'hddf1;
3355: douta=16'hcca8;
3356: douta=16'hcc25;
3357: douta=16'hcc46;
3358: douta=16'hcc67;
3359: douta=16'hcc67;
3360: douta=16'hd488;
3361: douta=16'hcc88;
3362: douta=16'hcc88;
3363: douta=16'hcc88;
3364: douta=16'hcc88;
3365: douta=16'hd4a9;
3366: douta=16'hd4a9;
3367: douta=16'hd488;
3368: douta=16'had31;
3369: douta=16'hcc68;
3370: douta=16'hcc88;
3371: douta=16'hcc68;
3372: douta=16'h8bcd;
3373: douta=16'hbd12;
3374: douta=16'hbd73;
3375: douta=16'hcd92;
3376: douta=16'h8c32;
3377: douta=16'h8c32;
3378: douta=16'h7bb0;
3379: douta=16'h630e;
3380: douta=16'h736f;
3381: douta=16'h5acc;
3382: douta=16'h526a;
3383: douta=16'h8c32;
3384: douta=16'h8432;
3385: douta=16'h634e;
3386: douta=16'h6c94;
3387: douta=16'hddb2;
3388: douta=16'ha368;
3389: douta=16'ha369;
3390: douta=16'h9b48;
3391: douta=16'h9b48;
3392: douta=16'ha515;
3393: douta=16'ha4f5;
3394: douta=16'h3125;
3395: douta=16'h424b;
3396: douta=16'h28c3;
3397: douta=16'h20e3;
3398: douta=16'h20a2;
3399: douta=16'h20a2;
3400: douta=16'h28e2;
3401: douta=16'h3103;
3402: douta=16'h3902;
3403: douta=16'h51c5;
3404: douta=16'h838b;
3405: douta=16'had30;
3406: douta=16'hbd71;
3407: douta=16'ha44c;
3408: douta=16'h8b07;
3409: douta=16'h8285;
3410: douta=16'h92c5;
3411: douta=16'h9306;
3412: douta=16'hab86;
3413: douta=16'hb3c7;
3414: douta=16'hbbe7;
3415: douta=16'hbc06;
3416: douta=16'hc447;
3417: douta=16'hc448;
3418: douta=16'hcc47;
3419: douta=16'hcc67;
3420: douta=16'hcc48;
3421: douta=16'hcc48;
3422: douta=16'hcc68;
3423: douta=16'hcc68;
3424: douta=16'hcc68;
3425: douta=16'hcc68;
3426: douta=16'hd488;
3427: douta=16'hcc88;
3428: douta=16'hd4a9;
3429: douta=16'hd489;
3430: douta=16'hd488;
3431: douta=16'hd4a9;
3432: douta=16'had32;
3433: douta=16'hd488;
3434: douta=16'hcc89;
3435: douta=16'hcc69;
3436: douta=16'h8bef;
3437: douta=16'ha4d4;
3438: douta=16'h9452;
3439: douta=16'h6b90;
3440: douta=16'h630e;
3441: douta=16'h630e;
3442: douta=16'h62ed;
3443: douta=16'h8bf1;
3444: douta=16'h7bb0;
3445: douta=16'h6b0d;
3446: douta=16'hffff;
3447: douta=16'hbb87;
3448: douta=16'haba8;
3449: douta=16'haba8;
3450: douta=16'ha388;
3451: douta=16'hab88;
3452: douta=16'ha388;
3453: douta=16'ha368;
3454: douta=16'ha368;
3455: douta=16'ha368;
3456: douta=16'h9cb4;
3457: douta=16'h8c96;
3458: douta=16'h28e3;
3459: douta=16'h28e3;
3460: douta=16'h20a3;
3461: douta=16'h20c3;
3462: douta=16'h2082;
3463: douta=16'h20c2;
3464: douta=16'h30e2;
3465: douta=16'h4143;
3466: douta=16'h49a6;
3467: douta=16'h59c4;
3468: douta=16'h61e4;
3469: douta=16'h6a04;
3470: douta=16'h7a84;
3471: douta=16'h82a5;
3472: douta=16'h8ac6;
3473: douta=16'h8ac6;
3474: douta=16'h9306;
3475: douta=16'h9326;
3476: douta=16'ha386;
3477: douta=16'hb3c7;
3478: douta=16'hbbe7;
3479: douta=16'hc407;
3480: douta=16'hc427;
3481: douta=16'hc428;
3482: douta=16'hcc47;
3483: douta=16'hcc47;
3484: douta=16'hcc68;
3485: douta=16'hcc48;
3486: douta=16'hcc68;
3487: douta=16'hcc68;
3488: douta=16'hcc69;
3489: douta=16'hcc88;
3490: douta=16'hcc89;
3491: douta=16'hcc88;
3492: douta=16'hd488;
3493: douta=16'hcc89;
3494: douta=16'hcc88;
3495: douta=16'hcc89;
3496: douta=16'had33;
3497: douta=16'hcc89;
3498: douta=16'hcc89;
3499: douta=16'hcc68;
3500: douta=16'hdc86;
3501: douta=16'h7390;
3502: douta=16'h6b4f;
3503: douta=16'h62ee;
3504: douta=16'h7b90;
3505: douta=16'h8431;
3506: douta=16'hffff;
3507: douta=16'hcbc7;
3508: douta=16'hbc08;
3509: douta=16'hb3c9;
3510: douta=16'hbbc9;
3511: douta=16'hb3c8;
3512: douta=16'hb3a8;
3513: douta=16'hb3a8;
3514: douta=16'hb3c8;
3515: douta=16'haba8;
3516: douta=16'hab88;
3517: douta=16'hab88;
3518: douta=16'hab88;
3519: douta=16'ha368;
3520: douta=16'hbd75;
3521: douta=16'h7c53;
3522: douta=16'h28e3;
3523: douta=16'h28e3;
3524: douta=16'h20c3;
3525: douta=16'h20a2;
3526: douta=16'h20c2;
3527: douta=16'h28e3;
3528: douta=16'h3103;
3529: douta=16'h4144;
3530: douta=16'h528b;
3531: douta=16'h59c4;
3532: douta=16'h6204;
3533: douta=16'h7203;
3534: douta=16'h7a84;
3535: douta=16'h8aa6;
3536: douta=16'h8ac6;
3537: douta=16'h9307;
3538: douta=16'h9b47;
3539: douta=16'h9326;
3540: douta=16'hab86;
3541: douta=16'hb3c7;
3542: douta=16'hbbe7;
3543: douta=16'hbc07;
3544: douta=16'hc427;
3545: douta=16'hc448;
3546: douta=16'hc447;
3547: douta=16'hcc67;
3548: douta=16'hcc68;
3549: douta=16'hcc68;
3550: douta=16'hcc68;
3551: douta=16'hcc68;
3552: douta=16'hcc68;
3553: douta=16'hd489;
3554: douta=16'hd489;
3555: douta=16'hd48a;
3556: douta=16'hd489;
3557: douta=16'hcc69;
3558: douta=16'hcc89;
3559: douta=16'hcc89;
3560: douta=16'had33;
3561: douta=16'hcc89;
3562: douta=16'hcc69;
3563: douta=16'hcc69;
3564: douta=16'hcc69;
3565: douta=16'hc449;
3566: douta=16'hd485;
3567: douta=16'hc428;
3568: douta=16'hcc4a;
3569: douta=16'hc448;
3570: douta=16'hc449;
3571: douta=16'hbc08;
3572: douta=16'hbc09;
3573: douta=16'hbc09;
3574: douta=16'hbbe9;
3575: douta=16'hb3e9;
3576: douta=16'hb3c8;
3577: douta=16'hb3c8;
3578: douta=16'hb3c8;
3579: douta=16'hb3a8;
3580: douta=16'haba9;
3581: douta=16'haba8;
3582: douta=16'ha388;
3583: douta=16'ha389;
3584: douta=16'h8c95;
3585: douta=16'h2082;
3586: douta=16'h28e3;
3587: douta=16'h28e3;
3588: douta=16'h20c3;
3589: douta=16'h20c2;
3590: douta=16'h28c3;
3591: douta=16'h28e2;
3592: douta=16'h3103;
3593: douta=16'h4143;
3594: douta=16'h31a7;
3595: douta=16'h59c4;
3596: douta=16'h6204;
3597: douta=16'h6a46;
3598: douta=16'h7a85;
3599: douta=16'h8aa6;
3600: douta=16'h8ac6;
3601: douta=16'h9306;
3602: douta=16'h7265;
3603: douta=16'h7a23;
3604: douta=16'haba6;
3605: douta=16'hb3e7;
3606: douta=16'hbc07;
3607: douta=16'hc428;
3608: douta=16'hc427;
3609: douta=16'hc448;
3610: douta=16'hc448;
3611: douta=16'hcc68;
3612: douta=16'hcc68;
3613: douta=16'hcc68;
3614: douta=16'hcc68;
3615: douta=16'hcc68;
3616: douta=16'hcc89;
3617: douta=16'hcc89;
3618: douta=16'hcc89;
3619: douta=16'hcc89;
3620: douta=16'hcc69;
3621: douta=16'hcc89;
3622: douta=16'hcc69;
3623: douta=16'hcc89;
3624: douta=16'had73;
3625: douta=16'hcc69;
3626: douta=16'hcc69;
3627: douta=16'hcc69;
3628: douta=16'hcc69;
3629: douta=16'hcc69;
3630: douta=16'hcc69;
3631: douta=16'hcc69;
3632: douta=16'hcc49;
3633: douta=16'hc449;
3634: douta=16'hc429;
3635: douta=16'hc429;
3636: douta=16'hbc09;
3637: douta=16'hbc09;
3638: douta=16'hbbe9;
3639: douta=16'hbbe9;
3640: douta=16'hb3e9;
3641: douta=16'hb3c8;
3642: douta=16'hb3c8;
3643: douta=16'haba9;
3644: douta=16'haba9;
3645: douta=16'hab88;
3646: douta=16'ha389;
3647: douta=16'ha368;
3648: douta=16'h94f7;
3649: douta=16'h28e3;
3650: douta=16'h28e3;
3651: douta=16'h28e3;
3652: douta=16'h20e3;
3653: douta=16'h20c2;
3654: douta=16'h28e3;
3655: douta=16'h28e3;
3656: douta=16'h3123;
3657: douta=16'h4963;
3658: douta=16'h0884;
3659: douta=16'h59c4;
3660: douta=16'h6a24;
3661: douta=16'h9cd1;
3662: douta=16'h7a85;
3663: douta=16'h82c6;
3664: douta=16'h8ae6;
3665: douta=16'h9306;
3666: douta=16'h8aa5;
3667: douta=16'h0000;
3668: douta=16'hb3c7;
3669: douta=16'hb3e7;
3670: douta=16'hbc07;
3671: douta=16'hc428;
3672: douta=16'hc428;
3673: douta=16'hc448;
3674: douta=16'hcc49;
3675: douta=16'hcc68;
3676: douta=16'hcc68;
3677: douta=16'hcc68;
3678: douta=16'hcc68;
3679: douta=16'hcc69;
3680: douta=16'hcc89;
3681: douta=16'hcc8a;
3682: douta=16'hcc89;
3683: douta=16'hcc89;
3684: douta=16'hcc8a;
3685: douta=16'hcc89;
3686: douta=16'hcc89;
3687: douta=16'hcc89;
3688: douta=16'hb594;
3689: douta=16'hcc69;
3690: douta=16'hcc69;
3691: douta=16'hcc89;
3692: douta=16'hcc69;
3693: douta=16'hcc69;
3694: douta=16'hcc69;
3695: douta=16'hcc49;
3696: douta=16'hc449;
3697: douta=16'hc429;
3698: douta=16'hc449;
3699: douta=16'hc429;
3700: douta=16'hbc29;
3701: douta=16'hbc09;
3702: douta=16'hbc09;
3703: douta=16'hb3e9;
3704: douta=16'hbc09;
3705: douta=16'hb3e9;
3706: douta=16'hb3c9;
3707: douta=16'haba9;
3708: douta=16'haba9;
3709: douta=16'haba8;
3710: douta=16'haba9;
3711: douta=16'ha389;
3712: douta=16'h9518;
3713: douta=16'h28e3;
3714: douta=16'h28e3;
3715: douta=16'h20e3;
3716: douta=16'h28e3;
3717: douta=16'h20c3;
3718: douta=16'h28e3;
3719: douta=16'h3103;
3720: douta=16'h3923;
3721: douta=16'h4964;
3722: douta=16'h3104;
3723: douta=16'h61e4;
3724: douta=16'h7245;
3725: douta=16'hacf0;
3726: douta=16'h7a85;
3727: douta=16'h82c6;
3728: douta=16'h8ae6;
3729: douta=16'h9b27;
3730: douta=16'hac4b;
3731: douta=16'hb44e;
3732: douta=16'haba7;
3733: douta=16'hbbe8;
3734: douta=16'hbc08;
3735: douta=16'hc407;
3736: douta=16'hc448;
3737: douta=16'hcc49;
3738: douta=16'hc449;
3739: douta=16'hc448;
3740: douta=16'hcc68;
3741: douta=16'hcc68;
3742: douta=16'hcc69;
3743: douta=16'hcc69;
3744: douta=16'hcc69;
3745: douta=16'hcc89;
3746: douta=16'hcc89;
3747: douta=16'hcc89;
3748: douta=16'hcc69;
3749: douta=16'hcc89;
3750: douta=16'hcc69;
3751: douta=16'hcc69;
3752: douta=16'hb594;
3753: douta=16'hcc69;
3754: douta=16'hcc69;
3755: douta=16'hcc69;
3756: douta=16'hcc69;
3757: douta=16'hcc69;
3758: douta=16'hcc69;
3759: douta=16'hc449;
3760: douta=16'hc449;
3761: douta=16'hc429;
3762: douta=16'hc429;
3763: douta=16'hc429;
3764: douta=16'hbc29;
3765: douta=16'hbc09;
3766: douta=16'hbc09;
3767: douta=16'hbc09;
3768: douta=16'hbbe9;
3769: douta=16'hb3e9;
3770: douta=16'hb3c9;
3771: douta=16'haba9;
3772: douta=16'haba9;
3773: douta=16'haba9;
3774: douta=16'haba9;
3775: douta=16'ha389;
3776: douta=16'h1861;
3777: douta=16'h20e3;
3778: douta=16'h2904;
3779: douta=16'h20e3;
3780: douta=16'h20a3;
3781: douta=16'h20c2;
3782: douta=16'h28e3;
3783: douta=16'h3103;
3784: douta=16'h3944;
3785: douta=16'h4964;
3786: douta=16'h6204;
3787: douta=16'h6204;
3788: douta=16'h6a44;
3789: douta=16'h7a85;
3790: douta=16'h82a5;
3791: douta=16'h82c6;
3792: douta=16'h8b07;
3793: douta=16'h9b47;
3794: douta=16'hde77;
3795: douta=16'hde76;
3796: douta=16'habc8;
3797: douta=16'hb3e8;
3798: douta=16'hbc08;
3799: douta=16'hc428;
3800: douta=16'hc448;
3801: douta=16'hc448;
3802: douta=16'hc448;
3803: douta=16'hc448;
3804: douta=16'hcc69;
3805: douta=16'hcc68;
3806: douta=16'hcc89;
3807: douta=16'hcc69;
3808: douta=16'hcc69;
3809: douta=16'hcc69;
3810: douta=16'hcc69;
3811: douta=16'hcc89;
3812: douta=16'hcc89;
3813: douta=16'hcc89;
3814: douta=16'hcc69;
3815: douta=16'hcc89;
3816: douta=16'hb595;
3817: douta=16'hcc6a;
3818: douta=16'hcc6a;
3819: douta=16'hcc69;
3820: douta=16'hcc49;
3821: douta=16'hc449;
3822: douta=16'hcc49;
3823: douta=16'hc449;
3824: douta=16'hc449;
3825: douta=16'hc449;
3826: douta=16'hc429;
3827: douta=16'hc429;
3828: douta=16'hc40a;
3829: douta=16'hbc2a;
3830: douta=16'hbc09;
3831: douta=16'hbc09;
3832: douta=16'hb3e9;
3833: douta=16'hb3e9;
3834: douta=16'hb3c9;
3835: douta=16'habc9;
3836: douta=16'habc9;
3837: douta=16'habc9;
3838: douta=16'haba9;
3839: douta=16'ha389;
3840: douta=16'h2904;
3841: douta=16'h2904;
3842: douta=16'h2904;
3843: douta=16'h20e3;
3844: douta=16'h20c2;
3845: douta=16'h28e3;
3846: douta=16'h2903;
3847: douta=16'h3903;
3848: douta=16'h4144;
3849: douta=16'h4a28;
3850: douta=16'h59c4;
3851: douta=16'h6204;
3852: douta=16'h7245;
3853: douta=16'h7244;
3854: douta=16'h82a6;
3855: douta=16'h8ae6;
3856: douta=16'h9307;
3857: douta=16'h9b47;
3858: douta=16'ha368;
3859: douta=16'ha388;
3860: douta=16'hb3c8;
3861: douta=16'hb3e8;
3862: douta=16'hbc08;
3863: douta=16'hbc28;
3864: douta=16'hc449;
3865: douta=16'hc449;
3866: douta=16'hc468;
3867: douta=16'hcc69;
3868: douta=16'hcc69;
3869: douta=16'hcc69;
3870: douta=16'hcc89;
3871: douta=16'hcc69;
3872: douta=16'hcc89;
3873: douta=16'hcc69;
3874: douta=16'hcc89;
3875: douta=16'hcc69;
3876: douta=16'hcc89;
3877: douta=16'hcc69;
3878: douta=16'hcc69;
3879: douta=16'hc489;
3880: douta=16'hb5d5;
3881: douta=16'hcc69;
3882: douta=16'hcc69;
3883: douta=16'hcc69;
3884: douta=16'hcc6a;
3885: douta=16'hcc6a;
3886: douta=16'hc449;
3887: douta=16'hc449;
3888: douta=16'hc449;
3889: douta=16'hc44a;
3890: douta=16'hc42a;
3891: douta=16'hbc29;
3892: douta=16'hbc0a;
3893: douta=16'hbc2a;
3894: douta=16'hbc09;
3895: douta=16'hbc09;
3896: douta=16'hbc09;
3897: douta=16'hb3e9;
3898: douta=16'hb3c9;
3899: douta=16'haba9;
3900: douta=16'habc9;
3901: douta=16'haba9;
3902: douta=16'ha389;
3903: douta=16'ha389;
3904: douta=16'h3125;
3905: douta=16'h2924;
3906: douta=16'h2904;
3907: douta=16'h2103;
3908: douta=16'h20e3;
3909: douta=16'h2903;
3910: douta=16'h28e3;
3911: douta=16'h3923;
3912: douta=16'h4143;
3913: douta=16'h4a4a;
3914: douta=16'h59e4;
3915: douta=16'h6a25;
3916: douta=16'h7224;
3917: douta=16'h7a85;
3918: douta=16'h82c6;
3919: douta=16'h8ae7;
3920: douta=16'h9327;
3921: douta=16'h9b47;
3922: douta=16'h9b68;
3923: douta=16'ha387;
3924: douta=16'hb3c8;
3925: douta=16'hb408;
3926: douta=16'hbc09;
3927: douta=16'hbc29;
3928: douta=16'hc449;
3929: douta=16'hc449;
3930: douta=16'hc469;
3931: douta=16'hcc8a;
3932: douta=16'hcc6a;
3933: douta=16'hcc69;
3934: douta=16'hcc69;
3935: douta=16'hcc6a;
3936: douta=16'hcc69;
3937: douta=16'hcc89;
3938: douta=16'hcc69;
3939: douta=16'hcc69;
3940: douta=16'hcc69;
3941: douta=16'hcc6a;
3942: douta=16'hcc69;
3943: douta=16'hcc6a;
3944: douta=16'hb5d5;
3945: douta=16'hcc6a;
3946: douta=16'hcc69;
3947: douta=16'hcc69;
3948: douta=16'hc46a;
3949: douta=16'hc469;
3950: douta=16'hc449;
3951: douta=16'hc469;
3952: douta=16'hc44a;
3953: douta=16'hc44a;
3954: douta=16'hc44a;
3955: douta=16'hbc2a;
3956: douta=16'hbc2a;
3957: douta=16'hbc0a;
3958: douta=16'hbc09;
3959: douta=16'hbbe9;
3960: douta=16'hbbe9;
3961: douta=16'hb3e9;
3962: douta=16'hb3c9;
3963: douta=16'habc9;
3964: douta=16'haba9;
3965: douta=16'haba9;
3966: douta=16'ha389;
3967: douta=16'ha389;
3968: douta=16'h2924;
3969: douta=16'h2904;
3970: douta=16'h2904;
3971: douta=16'h2104;
3972: douta=16'h20e3;
3973: douta=16'h28e3;
3974: douta=16'h3103;
3975: douta=16'h3923;
3976: douta=16'h4164;
3977: douta=16'h1906;
3978: douta=16'h59e5;
3979: douta=16'h6a25;
3980: douta=16'h7ae9;
3981: douta=16'h82a6;
3982: douta=16'h82c6;
3983: douta=16'h8ae7;
3984: douta=16'h8b07;
3985: douta=16'h9b28;
3986: douta=16'ha388;
3987: douta=16'ha387;
3988: douta=16'hb3e8;
3989: douta=16'hb409;
3990: douta=16'hbc2a;
3991: douta=16'hbc29;
3992: douta=16'hc449;
3993: douta=16'hc469;
3994: douta=16'hc46a;
3995: douta=16'hc46a;
3996: douta=16'hc48a;
3997: douta=16'hcc89;
3998: douta=16'hcc6a;
3999: douta=16'hc469;
4000: douta=16'hcc89;
4001: douta=16'hcc6a;
4002: douta=16'hcc6a;
4003: douta=16'hcc6a;
4004: douta=16'hcc6a;
4005: douta=16'hcc6a;
4006: douta=16'hcc6a;
4007: douta=16'hcc8a;
4008: douta=16'hbdd6;
4009: douta=16'hcc6a;
4010: douta=16'hc46a;
4011: douta=16'hc449;
4012: douta=16'hc44a;
4013: douta=16'hc469;
4014: douta=16'hc44a;
4015: douta=16'hc44a;
4016: douta=16'hc44a;
4017: douta=16'hc44a;
4018: douta=16'hbc2a;
4019: douta=16'hbc2a;
4020: douta=16'hbc2a;
4021: douta=16'hbc09;
4022: douta=16'hbc09;
4023: douta=16'hb3ea;
4024: douta=16'hb3e9;
4025: douta=16'hb3ca;
4026: douta=16'hb3e9;
4027: douta=16'haba9;
4028: douta=16'haba9;
4029: douta=16'ha389;
4030: douta=16'ha369;
4031: douta=16'ha389;
4032: douta=16'h2924;
4033: douta=16'h2104;
4034: douta=16'h2104;
4035: douta=16'h2924;
4036: douta=16'h20e3;
4037: douta=16'h28e3;
4038: douta=16'h3124;
4039: douta=16'h4144;
4040: douta=16'h4185;
4041: douta=16'h1084;
4042: douta=16'h59e4;
4043: douta=16'h6a25;
4044: douta=16'h94f4;
4045: douta=16'h82a7;
4046: douta=16'h82c6;
4047: douta=16'h8b07;
4048: douta=16'h9328;
4049: douta=16'h9b48;
4050: douta=16'h9b48;
4051: douta=16'ha388;
4052: douta=16'hb3e9;
4053: douta=16'hb409;
4054: douta=16'hbc2a;
4055: douta=16'hbc2a;
4056: douta=16'hc44a;
4057: douta=16'hc44a;
4058: douta=16'hc46a;
4059: douta=16'hc48a;
4060: douta=16'hc46a;
4061: douta=16'hcc8a;
4062: douta=16'hc46a;
4063: douta=16'hcc6a;
4064: douta=16'hcc6a;
4065: douta=16'hcc6a;
4066: douta=16'hc469;
4067: douta=16'hcc6a;
4068: douta=16'hc46a;
4069: douta=16'hcc6a;
4070: douta=16'hcc6a;
4071: douta=16'hc46a;
4072: douta=16'hbe16;
4073: douta=16'hc469;
4074: douta=16'hc469;
4075: douta=16'hc469;
4076: douta=16'hc46a;
4077: douta=16'hc44a;
4078: douta=16'hc44a;
4079: douta=16'hc44a;
4080: douta=16'hc44a;
4081: douta=16'hc42a;
4082: douta=16'hbc2a;
4083: douta=16'hbc2a;
4084: douta=16'hbc0a;
4085: douta=16'hbc09;
4086: douta=16'hb40a;
4087: douta=16'hb3ea;
4088: douta=16'hb3ea;
4089: douta=16'habca;
4090: douta=16'habca;
4091: douta=16'haba9;
4092: douta=16'habaa;
4093: douta=16'hab89;
4094: douta=16'ha389;
4095: douta=16'ha369;

default :douta  =	16'h	0000;
endcase
end


endmodule 
