
module bufferram (
  input [15:0] addra,      
  output reg [15:0] douta 
);

always@(*) begin
  case(addra)
0: douta=16'h74d9;
1: douta=16'h6cba;
2: douta=16'h32b0;
3: douta=16'h4311;
4: douta=16'h6436;
5: douta=16'h6c77;
6: douta=16'h6c14;
7: douta=16'h7414;
8: douta=16'h7c76;
9: douta=16'h6435;
10: douta=16'h31ea;
11: douta=16'h6c15;
12: douta=16'h31c8;
13: douta=16'hb536;
14: douta=16'ha536;
15: douta=16'hb597;
16: douta=16'h6bd3;
17: douta=16'h9516;
18: douta=16'h322d;
19: douta=16'h326f;
20: douta=16'h9d37;
21: douta=16'h9d36;
22: douta=16'hce19;
23: douta=16'h84b6;
24: douta=16'h8c95;
25: douta=16'h5bb2;
26: douta=16'h8494;
27: douta=16'h94f6;
28: douta=16'hc659;
29: douta=16'hd618;
30: douta=16'hffbc;
31: douta=16'h8454;
32: douta=16'h6b50;
33: douta=16'h6bd2;
34: douta=16'h5bd4;
35: douta=16'h94f5;
36: douta=16'he6fb;
37: douta=16'hd6da;
38: douta=16'h5b52;
39: douta=16'h8cb4;
40: douta=16'h63b2;
41: douta=16'had36;
42: douta=16'hd678;
43: douta=16'h94d6;
44: douta=16'hf77b;
45: douta=16'h7c75;
46: douta=16'had97;
47: douta=16'h3ad1;
48: douta=16'h7454;
49: douta=16'had77;
50: douta=16'hb5b8;
51: douta=16'he6b9;
52: douta=16'h94d6;
53: douta=16'had98;
54: douta=16'h9cd4;
55: douta=16'h5392;
56: douta=16'h3b11;
57: douta=16'hb5d8;
58: douta=16'ha576;
59: douta=16'h7415;
60: douta=16'hb5b8;
61: douta=16'h6c58;
62: douta=16'hd6ba;
63: douta=16'h2a90;
64: douta=16'h8cd3;
65: douta=16'h7cb6;
66: douta=16'hd6fa;
67: douta=16'hcebb;
68: douta=16'hae1b;
69: douta=16'h6437;
70: douta=16'h4b73;
71: douta=16'h6435;
72: douta=16'h7454;
73: douta=16'hc67a;
74: douta=16'ha598;
75: douta=16'had98;
76: douta=16'h5bd5;
77: douta=16'h94d6;
78: douta=16'h3b11;
79: douta=16'hb639;
80: douta=16'hbdd8;
81: douta=16'hce9b;
82: douta=16'h7c34;
83: douta=16'h6c76;
84: douta=16'h6c35;
85: douta=16'h7474;
86: douta=16'h9598;
87: douta=16'ha578;
88: douta=16'h7455;
89: douta=16'ha536;
90: douta=16'hadd8;
91: douta=16'h9d15;
92: douta=16'h21ab;
93: douta=16'h5b71;
94: douta=16'h2a2c;
95: douta=16'h7474;
96: douta=16'hbdd8;
97: douta=16'hf77c;
98: douta=16'hce18;
99: douta=16'hbdd7;
100: douta=16'h6b90;
101: douta=16'h8c92;
102: douta=16'h638f;
103: douta=16'he6f9;
104: douta=16'h8472;
105: douta=16'hd636;
106: douta=16'h9c30;
107: douta=16'h5b4f;
108: douta=16'h2169;
109: douta=16'h94d2;
110: douta=16'hce99;
111: douta=16'h6b90;
112: douta=16'hd677;
113: douta=16'h5a6b;
114: douta=16'h736f;
115: douta=16'h08a5;
116: douta=16'h52ee;
117: douta=16'h5b4f;
118: douta=16'h8c72;
119: douta=16'h9d14;
120: douta=16'ha4f2;
121: douta=16'h5b0e;
122: douta=16'h8c10;
123: douta=16'h8430;
124: douta=16'h0908;
125: douta=16'h1149;
126: douta=16'h6b6f;
127: douta=16'h5acc;
128: douta=16'he695;
129: douta=16'h5b30;
130: douta=16'hc5d6;
131: douta=16'h1109;
132: douta=16'h52ac;
133: douta=16'h324c;
134: douta=16'h326d;
135: douta=16'h29c9;
136: douta=16'h7411;
137: douta=16'ha4d3;
138: douta=16'h94b2;
139: douta=16'h94b4;
140: douta=16'h2966;
141: douta=16'h10e5;
142: douta=16'h0043;
143: douta=16'h7bcf;
144: douta=16'h8452;
145: douta=16'h5ace;
146: douta=16'h7c74;
147: douta=16'h42f0;
148: douta=16'h532f;
149: douta=16'h73f2;
150: douta=16'h94f5;
151: douta=16'h8453;
152: douta=16'h7c54;
153: douta=16'h4b31;
154: douta=16'h3ad0;
155: douta=16'h5b71;
156: douta=16'h3ace;
157: douta=16'hb5d7;
158: douta=16'h6bf4;
159: douta=16'ha515;
160: douta=16'h73f4;
161: douta=16'h19ee;
162: douta=16'h63f4;
163: douta=16'h9518;
164: douta=16'ha599;
165: douta=16'h74b8;
166: douta=16'ha558;
167: douta=16'h4373;
168: douta=16'h5bd4;
169: douta=16'h4b11;
170: douta=16'h5371;
171: douta=16'h84d5;
172: douta=16'h6c99;
173: douta=16'h7cb8;
174: douta=16'h7d19;
175: douta=16'h2a6f;
176: douta=16'h5352;
177: douta=16'h5b92;
178: douta=16'ha5bb;
179: douta=16'h74d9;
180: douta=16'h118a;
181: douta=16'h19ed;
182: douta=16'h6c55;
183: douta=16'h7476;
184: douta=16'h8d7c;
185: douta=16'h7cd9;
186: douta=16'h2b35;
187: douta=16'h4b53;
188: douta=16'h6c57;
189: douta=16'h8519;
190: douta=16'h3b54;
191: douta=16'h5c37;
192: douta=16'h5c57;
193: douta=16'h4b52;
194: douta=16'h3b11;
195: douta=16'h4b31;
196: douta=16'h8519;
197: douta=16'h74b8;
198: douta=16'h6c35;
199: douta=16'h5351;
200: douta=16'h63b3;
201: douta=16'h63d4;
202: douta=16'hc61a;
203: douta=16'h9537;
204: douta=16'hb5f9;
205: douta=16'h73f3;
206: douta=16'h6c13;
207: douta=16'h52f0;
208: douta=16'h9517;
209: douta=16'h8495;
210: douta=16'hce39;
211: douta=16'h9d37;
212: douta=16'hd6ba;
213: douta=16'hde99;
214: douta=16'had57;
215: douta=16'h3312;
216: douta=16'h7414;
217: douta=16'hadb8;
218: douta=16'hbdf7;
219: douta=16'hd679;
220: douta=16'h9d99;
221: douta=16'h8c53;
222: douta=16'hcdf8;
223: douta=16'hc618;
224: douta=16'h8c52;
225: douta=16'hbdf7;
226: douta=16'hce59;
227: douta=16'hb5b8;
228: douta=16'hd6bb;
229: douta=16'h7434;
230: douta=16'h3a6f;
231: douta=16'h8c94;
232: douta=16'hc619;
233: douta=16'hc5f8;
234: douta=16'hc5f8;
235: douta=16'h326f;
236: douta=16'h6c54;
237: douta=16'h5b91;
238: douta=16'hb5d8;
239: douta=16'he719;
240: douta=16'h9d37;
241: douta=16'hef3b;
242: douta=16'hce7b;
243: douta=16'hbd97;
244: douta=16'h3ab0;
245: douta=16'h94d4;
246: douta=16'h84b5;
247: douta=16'h9d35;
248: douta=16'ha517;
249: douta=16'hdefb;
250: douta=16'hd679;
251: douta=16'h8475;
252: douta=16'h7455;
253: douta=16'h74d8;
254: douta=16'h8cb6;
255: douta=16'h9516;
256: douta=16'h9d99;
257: douta=16'ha516;
258: douta=16'hc6bd;
259: douta=16'hc618;
260: douta=16'h4b52;
261: douta=16'h3a90;
262: douta=16'h7434;
263: douta=16'hbe39;
264: douta=16'hae1b;
265: douta=16'h9559;
266: douta=16'h5bb5;
267: douta=16'h63b4;
268: douta=16'h2a4e;
269: douta=16'h5bd3;
270: douta=16'h9558;
271: douta=16'had57;
272: douta=16'heefa;
273: douta=16'h6cb8;
274: douta=16'h7435;
275: douta=16'h8cf7;
276: douta=16'h9579;
277: douta=16'hb619;
278: douta=16'hadda;
279: douta=16'hc69b;
280: douta=16'h6351;
281: douta=16'hd67a;
282: douta=16'h4b32;
283: douta=16'h326d;
284: douta=16'h84d4;
285: douta=16'h7412;
286: douta=16'hceba;
287: douta=16'ha577;
288: douta=16'h63d2;
289: douta=16'h6392;
290: douta=16'h4a8c;
291: douta=16'h1948;
292: douta=16'ha535;
293: douta=16'hce78;
294: douta=16'ha492;
295: douta=16'h7390;
296: douta=16'ha491;
297: douta=16'h320a;
298: douta=16'h7411;
299: douta=16'hb595;
300: douta=16'hc5f7;
301: douta=16'h94d4;
302: douta=16'h42ef;
303: douta=16'h4a2a;
304: douta=16'h322a;
305: douta=16'h5b2c;
306: douta=16'h632d;
307: douta=16'hdeb7;
308: douta=16'h9c91;
309: douta=16'hce17;
310: douta=16'h83af;
311: douta=16'h94b4;
312: douta=16'h4a4a;
313: douta=16'h3a4b;
314: douta=16'h9d53;
315: douta=16'h9d34;
316: douta=16'h9d14;
317: douta=16'h8432;
318: douta=16'h8c51;
319: douta=16'h634f;
320: douta=16'h8411;
321: douta=16'h7bf0;
322: douta=16'h322b;
323: douta=16'h636f;
324: douta=16'hce57;
325: douta=16'hce57;
326: douta=16'h4aaf;
327: douta=16'hbdb5;
328: douta=16'h08e8;
329: douta=16'h42ad;
330: douta=16'h322c;
331: douta=16'h63b0;
332: douta=16'h3187;
333: douta=16'h10c5;
334: douta=16'h18e6;
335: douta=16'h4aef;
336: douta=16'h94d3;
337: douta=16'h21a9;
338: douta=16'h1968;
339: douta=16'h5b6e;
340: douta=16'h8433;
341: douta=16'h7c13;
342: douta=16'h42af;
343: douta=16'h29eb;
344: douta=16'h530f;
345: douta=16'h7433;
346: douta=16'hb534;
347: douta=16'hc617;
348: douta=16'h6c15;
349: douta=16'h3aae;
350: douta=16'h7412;
351: douta=16'h2ad1;
352: douta=16'h7454;
353: douta=16'h9516;
354: douta=16'hde9a;
355: douta=16'h7477;
356: douta=16'h4333;
357: douta=16'h4331;
358: douta=16'h4b53;
359: douta=16'h84d5;
360: douta=16'h6c55;
361: douta=16'ha5db;
362: douta=16'h6b71;
363: douta=16'h6436;
364: douta=16'h5330;
365: douta=16'h6416;
366: douta=16'h3b52;
367: douta=16'h9517;
368: douta=16'h6c36;
369: douta=16'h4b53;
370: douta=16'h2a4f;
371: douta=16'h19cc;
372: douta=16'h4311;
373: douta=16'h5c57;
374: douta=16'h7c35;
375: douta=16'h84f8;
376: douta=16'h3b54;
377: douta=16'h6499;
378: douta=16'h2270;
379: douta=16'h7cd9;
380: douta=16'h84f9;
381: douta=16'h4b75;
382: douta=16'h1a2f;
383: douta=16'h5c15;
384: douta=16'h6c97;
385: douta=16'h53b4;
386: douta=16'h6457;
387: douta=16'h4b32;
388: douta=16'h53b4;
389: douta=16'h53f5;
390: douta=16'h5352;
391: douta=16'h7c75;
392: douta=16'h9517;
393: douta=16'h8497;
394: douta=16'h4333;
395: douta=16'h5311;
396: douta=16'h5b51;
397: douta=16'h9cd5;
398: douta=16'had98;
399: douta=16'hde99;
400: douta=16'hadd9;
401: douta=16'h8455;
402: douta=16'h6bd2;
403: douta=16'h63b4;
404: douta=16'h8c95;
405: douta=16'h7454;
406: douta=16'hbdf7;
407: douta=16'h84d7;
408: douta=16'ha578;
409: douta=16'had37;
410: douta=16'hbdd8;
411: douta=16'h5bb4;
412: douta=16'hce7a;
413: douta=16'ha598;
414: douta=16'he71a;
415: douta=16'hd69a;
416: douta=16'hbdb6;
417: douta=16'hce38;
418: douta=16'h63d3;
419: douta=16'h73f2;
420: douta=16'hc638;
421: douta=16'hcebb;
422: douta=16'h73b2;
423: douta=16'hf75b;
424: douta=16'h9d77;
425: douta=16'h4333;
426: douta=16'hb596;
427: douta=16'had36;
428: douta=16'hbe7a;
429: douta=16'h9516;
430: douta=16'hc699;
431: douta=16'h9d36;
432: douta=16'h3b11;
433: douta=16'h8412;
434: douta=16'hd658;
435: douta=16'hef3a;
436: douta=16'hb5b6;
437: douta=16'hd6b9;
438: douta=16'h9d78;
439: douta=16'h7496;
440: douta=16'h3b11;
441: douta=16'h6371;
442: douta=16'h84b6;
443: douta=16'hc5f8;
444: douta=16'hdefb;
445: douta=16'hbe19;
446: douta=16'hc67a;
447: douta=16'h7435;
448: douta=16'h84d5;
449: douta=16'h2af0;
450: douta=16'h4332;
451: douta=16'hdeba;
452: douta=16'h9d58;
453: douta=16'hd679;
454: douta=16'h8496;
455: douta=16'h8c95;
456: douta=16'h2250;
457: douta=16'h4332;
458: douta=16'h84d6;
459: douta=16'he75d;
460: douta=16'h7c77;
461: douta=16'h8538;
462: douta=16'h5bd5;
463: douta=16'h9d58;
464: douta=16'h9599;
465: douta=16'h7c96;
466: douta=16'hc69b;
467: douta=16'hbe39;
468: douta=16'h9dba;
469: douta=16'hd69b;
470: douta=16'h3b32;
471: douta=16'h63d3;
472: douta=16'had55;
473: douta=16'hce59;
474: douta=16'h9cb6;
475: douta=16'h6c13;
476: douta=16'ha536;
477: douta=16'hce59;
478: douta=16'h19cd;
479: douta=16'h21cd;
480: douta=16'hadb8;
481: douta=16'h8433;
482: douta=16'had55;
483: douta=16'h7c32;
484: douta=16'h8c52;
485: douta=16'h2188;
486: douta=16'h530f;
487: douta=16'had54;
488: douta=16'ha555;
489: douta=16'h7c51;
490: douta=16'h9514;
491: douta=16'h5aee;
492: douta=16'h5b0f;
493: douta=16'h8493;
494: douta=16'h9cd3;
495: douta=16'ha4b2;
496: douta=16'h52ac;
497: douta=16'h8c51;
498: douta=16'h4a8c;
499: douta=16'h424c;
500: douta=16'h634e;
501: douta=16'h3a6b;
502: douta=16'heef9;
503: douta=16'hbdb5;
504: douta=16'hd657;
505: douta=16'h41c9;
506: douta=16'h8c71;
507: douta=16'h5b2f;
508: douta=16'h7c12;
509: douta=16'h636f;
510: douta=16'h9cd3;
511: douta=16'h8431;
512: douta=16'h73d0;
513: douta=16'hc5d6;
514: douta=16'h6b4f;
515: douta=16'h6391;
516: douta=16'h2a2d;
517: douta=16'h21c9;
518: douta=16'h2989;
519: douta=16'hd657;
520: douta=16'hcdd4;
521: douta=16'h9cf3;
522: douta=16'hbdb5;
523: douta=16'h5b0d;
524: douta=16'h2105;
525: douta=16'h10c4;
526: douta=16'h10e5;
527: douta=16'h3a4c;
528: douta=16'h5b4f;
529: douta=16'h94b3;
530: douta=16'h52ce;
531: douta=16'h73b0;
532: douta=16'h4ace;
533: douta=16'h7bf1;
534: douta=16'h6bb1;
535: douta=16'h9cb3;
536: douta=16'h9d37;
537: douta=16'h63d3;
538: douta=16'h5bd3;
539: douta=16'h2a2d;
540: douta=16'h6bd2;
541: douta=16'h9c94;
542: douta=16'hbdb7;
543: douta=16'h7434;
544: douta=16'h328f;
545: douta=16'h4b31;
546: douta=16'h3ad0;
547: douta=16'h8cf8;
548: douta=16'h6c34;
549: douta=16'hce5a;
550: douta=16'h6436;
551: douta=16'h19ee;
552: douta=16'h3aaf;
553: douta=16'h11ac;
554: douta=16'h4b31;
555: douta=16'h5bf5;
556: douta=16'h8d19;
557: douta=16'h8d18;
558: douta=16'h6457;
559: douta=16'h9559;
560: douta=16'h21ce;
561: douta=16'h4b72;
562: douta=16'h8517;
563: douta=16'h8d18;
564: douta=16'h4b51;
565: douta=16'h11ed;
566: douta=16'h6435;
567: douta=16'h5bd4;
568: douta=16'h9e1d;
569: douta=16'h5c15;
570: douta=16'h5c38;
571: douta=16'h3ad2;
572: douta=16'h53d5;
573: douta=16'h5bb2;
574: douta=16'h6436;
575: douta=16'h5bf7;
576: douta=16'h2a6f;
577: douta=16'h32d1;
578: douta=16'h4353;
579: douta=16'h4b53;
580: douta=16'h7cf9;
581: douta=16'h7d3b;
582: douta=16'h5352;
583: douta=16'h7c56;
584: douta=16'h7434;
585: douta=16'h7435;
586: douta=16'h8d18;
587: douta=16'h84b7;
588: douta=16'h94d6;
589: douta=16'h428e;
590: douta=16'h6b91;
591: douta=16'ha536;
592: douta=16'h94d6;
593: douta=16'hce38;
594: douta=16'hadb8;
595: douta=16'h7476;
596: douta=16'h7c34;
597: douta=16'h7455;
598: douta=16'h8cd6;
599: douta=16'h84b6;
600: douta=16'h9516;
601: douta=16'hef3c;
602: douta=16'hef5b;
603: douta=16'h9d58;
604: douta=16'h7cd7;
605: douta=16'h6bb3;
606: douta=16'hb5b8;
607: douta=16'hce59;
608: douta=16'hdeba;
609: douta=16'he6da;
610: douta=16'h7475;
611: douta=16'h7c12;
612: douta=16'hc619;
613: douta=16'h8494;
614: douta=16'hde58;
615: douta=16'hded9;
616: douta=16'hd6da;
617: douta=16'h9cf7;
618: douta=16'h8c93;
619: douta=16'h94f5;
620: douta=16'h84b5;
621: douta=16'h8474;
622: douta=16'he71b;
623: douta=16'had98;
624: douta=16'h6c36;
625: douta=16'ha4d4;
626: douta=16'hb5f8;
627: douta=16'ha577;
628: douta=16'ha556;
629: douta=16'hdeb9;
630: douta=16'h9537;
631: douta=16'h63f4;
632: douta=16'h6bf4;
633: douta=16'hb5f9;
634: douta=16'h9599;
635: douta=16'h7bd0;
636: douta=16'hae19;
637: douta=16'h8cf6;
638: douta=16'hbe5b;
639: douta=16'hadb8;
640: douta=16'h9d98;
641: douta=16'h7415;
642: douta=16'h7477;
643: douta=16'hb5d8;
644: douta=16'h7c74;
645: douta=16'hc619;
646: douta=16'hb5f9;
647: douta=16'hbe19;
648: douta=16'h32b1;
649: douta=16'h11ce;
650: douta=16'h4b74;
651: douta=16'ha596;
652: douta=16'hbdd8;
653: douta=16'h9dda;
654: douta=16'h9518;
655: douta=16'hdefc;
656: douta=16'h74f8;
657: douta=16'h4b53;
658: douta=16'h6c55;
659: douta=16'h9538;
660: douta=16'h5bd5;
661: douta=16'he71b;
662: douta=16'h9518;
663: douta=16'h63d2;
664: douta=16'h7c12;
665: douta=16'h9d77;
666: douta=16'h8473;
667: douta=16'h7c74;
668: douta=16'hbdd7;
669: douta=16'hff7c;
670: douta=16'h5bf5;
671: douta=16'h42d0;
672: douta=16'h324e;
673: douta=16'h426d;
674: douta=16'had96;
675: douta=16'h8c94;
676: douta=16'hb596;
677: douta=16'h632e;
678: douta=16'h8474;
679: douta=16'h52ec;
680: douta=16'h5b4e;
681: douta=16'h9cf3;
682: douta=16'h8472;
683: douta=16'hc5d6;
684: douta=16'h7c31;
685: douta=16'h0907;
686: douta=16'h4a6a;
687: douta=16'h9450;
688: douta=16'ha470;
689: douta=16'h9471;
690: douta=16'h3a0b;
691: douta=16'h632e;
692: douta=16'h8c50;
693: douta=16'h3a0a;
694: douta=16'h7c31;
695: douta=16'h7c11;
696: douta=16'hce77;
697: douta=16'hacf3;
698: douta=16'h7c10;
699: douta=16'h634f;
700: douta=16'h4aad;
701: douta=16'h29ea;
702: douta=16'h2187;
703: douta=16'h6b8f;
704: douta=16'h94d4;
705: douta=16'he6d8;
706: douta=16'h630d;
707: douta=16'h9d16;
708: douta=16'h6414;
709: douta=16'h0884;
710: douta=16'h0043;
711: douta=16'h5b2f;
712: douta=16'h8450;
713: douta=16'h9cb2;
714: douta=16'hc5b4;
715: douta=16'h9cd2;
716: douta=16'h18c4;
717: douta=16'h10c5;
718: douta=16'h1926;
719: douta=16'h1949;
720: douta=16'h1149;
721: douta=16'h9d15;
722: douta=16'h73d1;
723: douta=16'h9493;
724: douta=16'h4aae;
725: douta=16'h5b4f;
726: douta=16'h29a9;
727: douta=16'h9d14;
728: douta=16'h6bd1;
729: douta=16'h5b70;
730: douta=16'h7c55;
731: douta=16'h63d3;
732: douta=16'h21cb;
733: douta=16'hce58;
734: douta=16'h9d37;
735: douta=16'hde9a;
736: douta=16'h6415;
737: douta=16'h9d59;
738: douta=16'h4b74;
739: douta=16'h5373;
740: douta=16'h7414;
741: douta=16'h9d37;
742: douta=16'hadda;
743: douta=16'h52d0;
744: douta=16'h84b7;
745: douta=16'h328f;
746: douta=16'h222f;
747: douta=16'h4353;
748: douta=16'ha5ba;
749: douta=16'h9d79;
750: douta=16'h84b7;
751: douta=16'h6c77;
752: douta=16'h3b53;
753: douta=16'h53f7;
754: douta=16'h63d2;
755: douta=16'h84f7;
756: douta=16'hbdfa;
757: douta=16'h63f4;
758: douta=16'h3af1;
759: douta=16'h4311;
760: douta=16'h3b74;
761: douta=16'ha5da;
762: douta=16'h53d6;
763: douta=16'h6479;
764: douta=16'h32f3;
765: douta=16'h4b73;
766: douta=16'h9559;
767: douta=16'h53f6;
768: douta=16'h4b73;
769: douta=16'h5bd4;
770: douta=16'h6458;
771: douta=16'h5373;
772: douta=16'h7477;
773: douta=16'h53b4;
774: douta=16'h116a;
775: douta=16'h7c96;
776: douta=16'h84b6;
777: douta=16'ha579;
778: douta=16'h8495;
779: douta=16'h9517;
780: douta=16'h5b92;
781: douta=16'had56;
782: douta=16'ha576;
783: douta=16'had77;
784: douta=16'h6c36;
785: douta=16'h8cf6;
786: douta=16'h8433;
787: douta=16'h63d3;
788: douta=16'h42d0;
789: douta=16'h9d36;
790: douta=16'hc618;
791: douta=16'hb5d9;
792: douta=16'ha599;
793: douta=16'h9d36;
794: douta=16'hbdd7;
795: douta=16'h222e;
796: douta=16'hadd8;
797: douta=16'h9d17;
798: douta=16'hdeda;
799: douta=16'hce9a;
800: douta=16'hb5b8;
801: douta=16'ha516;
802: douta=16'h5392;
803: douta=16'h8473;
804: douta=16'hb5b7;
805: douta=16'hd6b9;
806: douta=16'ha4f5;
807: douta=16'hf6fb;
808: douta=16'h8d16;
809: douta=16'h2a8f;
810: douta=16'ha576;
811: douta=16'hb576;
812: douta=16'hbe59;
813: douta=16'ha557;
814: douta=16'hbe9a;
815: douta=16'h8c53;
816: douta=16'h5351;
817: douta=16'hce37;
818: douta=16'hc659;
819: douta=16'hf77c;
820: douta=16'h9d15;
821: douta=16'hbe18;
822: douta=16'h8495;
823: douta=16'h32d1;
824: douta=16'h5bb3;
825: douta=16'h8c95;
826: douta=16'ha5d8;
827: douta=16'hd679;
828: douta=16'he6fb;
829: douta=16'hb5b9;
830: douta=16'h8519;
831: douta=16'h83f3;
832: douta=16'h5372;
833: douta=16'h3a8f;
834: douta=16'h84b6;
835: douta=16'hb5f8;
836: douta=16'hef1b;
837: douta=16'hbe9b;
838: douta=16'h7c34;
839: douta=16'h6415;
840: douta=16'h4b0f;
841: douta=16'h9578;
842: douta=16'ha5da;
843: douta=16'h84d6;
844: douta=16'hd6bb;
845: douta=16'h8496;
846: douta=16'hc619;
847: douta=16'ha5fb;
848: douta=16'h5bf5;
849: douta=16'h5353;
850: douta=16'h84d7;
851: douta=16'hbe7b;
852: douta=16'h6c77;
853: douta=16'hb65b;
854: douta=16'h6393;
855: douta=16'h21ab;
856: douta=16'h9d55;
857: douta=16'h84b5;
858: douta=16'hbe18;
859: douta=16'h94b5;
860: douta=16'hce59;
861: douta=16'h5bb2;
862: douta=16'h322d;
863: douta=16'h6bb3;
864: douta=16'h9db8;
865: douta=16'hacd4;
866: douta=16'h8473;
867: douta=16'h5330;
868: douta=16'h322b;
869: douta=16'h632f;
870: douta=16'h4aad;
871: douta=16'h8c72;
872: douta=16'ha555;
873: douta=16'h9cb3;
874: douta=16'h630d;
875: douta=16'h5b0e;
876: douta=16'h73af;
877: douta=16'h736e;
878: douta=16'had12;
879: douta=16'h94b1;
880: douta=16'hcdf5;
881: douta=16'h1969;
882: douta=16'h1107;
883: douta=16'h9cd3;
884: douta=16'hde99;
885: douta=16'h9451;
886: douta=16'h530f;
887: douta=16'h4a8d;
888: douta=16'h6b8f;
889: douta=16'h428b;
890: douta=16'h5b6f;
891: douta=16'h7c31;
892: douta=16'h7c11;
893: douta=16'ha514;
894: douta=16'h5b0d;
895: douta=16'h39eb;
896: douta=16'h9410;
897: douta=16'h3a8e;
898: douta=16'h530e;
899: douta=16'h5b4f;
900: douta=16'h8431;
901: douta=16'h73f1;
902: douta=16'hce36;
903: douta=16'h5b71;
904: douta=16'h5b51;
905: douta=16'h6bb1;
906: douta=16'h320c;
907: douta=16'h8472;
908: douta=16'h18e4;
909: douta=16'h10c4;
910: douta=16'h29c8;
911: douta=16'h94d2;
912: douta=16'h8451;
913: douta=16'h52ce;
914: douta=16'h5b51;
915: douta=16'h1108;
916: douta=16'h6bd1;
917: douta=16'h6b90;
918: douta=16'hd636;
919: douta=16'ha555;
920: douta=16'h52ef;
921: douta=16'h9d15;
922: douta=16'h7411;
923: douta=16'h322c;
924: douta=16'had75;
925: douta=16'h7c55;
926: douta=16'hde9a;
927: douta=16'h5c16;
928: douta=16'h4b31;
929: douta=16'h84b5;
930: douta=16'h7c95;
931: douta=16'had77;
932: douta=16'h9d58;
933: douta=16'h9d58;
934: douta=16'h3a8f;
935: douta=16'h3290;
936: douta=16'h19ee;
937: douta=16'h7c95;
938: douta=16'h9536;
939: douta=16'hadba;
940: douta=16'h6cb9;
941: douta=16'h32b1;
942: douta=16'h6436;
943: douta=16'h3b53;
944: douta=16'h4332;
945: douta=16'h84f8;
946: douta=16'h3b34;
947: douta=16'h7455;
948: douta=16'h222e;
949: douta=16'h2a4f;
950: douta=16'ha5b9;
951: douta=16'hb65c;
952: douta=16'h84b7;
953: douta=16'h5c17;
954: douta=16'h959b;
955: douta=16'h11ac;
956: douta=16'h63f4;
957: douta=16'h6c78;
958: douta=16'h4355;
959: douta=16'h5395;
960: douta=16'h6c98;
961: douta=16'h5c17;
962: douta=16'h4bf6;
963: douta=16'h4b32;
964: douta=16'h63d4;
965: douta=16'h7cd8;
966: douta=16'h6c56;
967: douta=16'h7c35;
968: douta=16'h5351;
969: douta=16'h4b31;
970: douta=16'h7c75;
971: douta=16'had98;
972: douta=16'hce5a;
973: douta=16'h94f5;
974: douta=16'h5bd3;
975: douta=16'h428f;
976: douta=16'h3ad0;
977: douta=16'h6bf1;
978: douta=16'hc639;
979: douta=16'hbe3a;
980: douta=16'h9d78;
981: douta=16'hd6ba;
982: douta=16'ha577;
983: douta=16'h5372;
984: douta=16'h6bd3;
985: douta=16'hc639;
986: douta=16'he6da;
987: douta=16'h9d36;
988: douta=16'hce7a;
989: douta=16'h9495;
990: douta=16'he6bb;
991: douta=16'h7c54;
992: douta=16'had97;
993: douta=16'heed9;
994: douta=16'ha578;
995: douta=16'hbdd8;
996: douta=16'had98;
997: douta=16'h6bd2;
998: douta=16'h7c53;
999: douta=16'ha534;
1000: douta=16'hce58;
1001: douta=16'ha4f5;
1002: douta=16'hf75a;
1003: douta=16'h7bf0;
1004: douta=16'h6415;
1005: douta=16'h4312;
1006: douta=16'hdeba;
1007: douta=16'he73a;
1008: douta=16'ha557;
1009: douta=16'hf77d;
1010: douta=16'h5c36;
1011: douta=16'h9c93;
1012: douta=16'h21ab;
1013: douta=16'h9515;
1014: douta=16'hbdd6;
1015: douta=16'ha578;
1016: douta=16'hce7a;
1017: douta=16'h6c56;
1018: douta=16'h7495;
1019: douta=16'h63f3;
1020: douta=16'h426d;
1021: douta=16'h7474;
1022: douta=16'ha557;
1023: douta=16'he6b9;
1024: douta=16'h6bd3;
1025: douta=16'heed9;
1026: douta=16'h53d5;
1027: douta=16'h5bb4;
1028: douta=16'h84f7;
1029: douta=16'h4b71;
1030: douta=16'had98;
1031: douta=16'h8d38;
1032: douta=16'hd67a;
1033: douta=16'h32b0;
1034: douta=16'h7c14;
1035: douta=16'h7496;
1036: douta=16'h6414;
1037: douta=16'h7454;
1038: douta=16'h84b4;
1039: douta=16'hd6fb;
1040: douta=16'h6c98;
1041: douta=16'hdf1d;
1042: douta=16'h8cf8;
1043: douta=16'h7434;
1044: douta=16'h63b4;
1045: douta=16'h84d7;
1046: douta=16'h9577;
1047: douta=16'h9517;
1048: douta=16'hb5f8;
1049: douta=16'h5331;
1050: douta=16'h63b1;
1051: douta=16'h63b2;
1052: douta=16'h9536;
1053: douta=16'h7412;
1054: douta=16'h9d57;
1055: douta=16'had76;
1056: douta=16'h6c13;
1057: douta=16'h8c93;
1058: douta=16'h3a4c;
1059: douta=16'h3a8e;
1060: douta=16'h5330;
1061: douta=16'hef3a;
1062: douta=16'h3a4c;
1063: douta=16'h4aac;
1064: douta=16'h0885;
1065: douta=16'h6b8e;
1066: douta=16'hce78;
1067: douta=16'h738f;
1068: douta=16'hcdf6;
1069: douta=16'h944e;
1070: douta=16'hce14;
1071: douta=16'h31ea;
1072: douta=16'h638f;
1073: douta=16'ha512;
1074: douta=16'he6b7;
1075: douta=16'hb575;
1076: douta=16'h31ec;
1077: douta=16'h7bd0;
1078: douta=16'ha4d3;
1079: douta=16'had75;
1080: douta=16'h73af;
1081: douta=16'hd698;
1082: douta=16'h8433;
1083: douta=16'ha516;
1084: douta=16'h08a4;
1085: douta=16'h0063;
1086: douta=16'h73f1;
1087: douta=16'h8c52;
1088: douta=16'ha575;
1089: douta=16'h5b70;
1090: douta=16'h8453;
1091: douta=16'h21cb;
1092: douta=16'h322c;
1093: douta=16'h5350;
1094: douta=16'h63f2;
1095: douta=16'h8454;
1096: douta=16'h8c72;
1097: douta=16'h8473;
1098: douta=16'h5b2f;
1099: douta=16'h94f5;
1100: douta=16'h18a3;
1101: douta=16'h08c4;
1102: douta=16'h1906;
1103: douta=16'h2189;
1104: douta=16'h6bb0;
1105: douta=16'hb555;
1106: douta=16'h7c12;
1107: douta=16'h8453;
1108: douta=16'h39e9;
1109: douta=16'h52cd;
1110: douta=16'h29ca;
1111: douta=16'h530f;
1112: douta=16'hff58;
1113: douta=16'hc5f6;
1114: douta=16'ha515;
1115: douta=16'h3a4c;
1116: douta=16'h5331;
1117: douta=16'hb5d7;
1118: douta=16'h9d57;
1119: douta=16'h63b2;
1120: douta=16'h5373;
1121: douta=16'h9539;
1122: douta=16'h32d2;
1123: douta=16'h224e;
1124: douta=16'h3aaf;
1125: douta=16'h84b4;
1126: douta=16'hbe59;
1127: douta=16'h5bf5;
1128: douta=16'h2a2e;
1129: douta=16'h012b;
1130: douta=16'h3af0;
1131: douta=16'h4312;
1132: douta=16'h6c56;
1133: douta=16'hc639;
1134: douta=16'h9518;
1135: douta=16'h5c16;
1136: douta=16'h32d2;
1137: douta=16'h222e;
1138: douta=16'h7c75;
1139: douta=16'h8d19;
1140: douta=16'h9538;
1141: douta=16'h53f6;
1142: douta=16'h63f5;
1143: douta=16'h11ac;
1144: douta=16'h2270;
1145: douta=16'h7497;
1146: douta=16'h8519;
1147: douta=16'h857c;
1148: douta=16'h5438;
1149: douta=16'h3312;
1150: douta=16'h3ad0;
1151: douta=16'ha5da;
1152: douta=16'h6c78;
1153: douta=16'h74d9;
1154: douta=16'h43b5;
1155: douta=16'h4311;
1156: douta=16'h5bb3;
1157: douta=16'h5b94;
1158: douta=16'h5393;
1159: douta=16'h9518;
1160: douta=16'h7c75;
1161: douta=16'h6bf4;
1162: douta=16'h6b92;
1163: douta=16'h84b7;
1164: douta=16'h94d6;
1165: douta=16'hce59;
1166: douta=16'h9d57;
1167: douta=16'h9d16;
1168: douta=16'h63b2;
1169: douta=16'h5330;
1170: douta=16'h6bf3;
1171: douta=16'h7cb6;
1172: douta=16'h8cd5;
1173: douta=16'hbdd8;
1174: douta=16'hce18;
1175: douta=16'h7cb6;
1176: douta=16'h6bd2;
1177: douta=16'h94f6;
1178: douta=16'h94d5;
1179: douta=16'ha576;
1180: douta=16'hc679;
1181: douta=16'hde59;
1182: douta=16'hff9b;
1183: douta=16'h6bd3;
1184: douta=16'h8c95;
1185: douta=16'hd679;
1186: douta=16'h9d15;
1187: douta=16'hde98;
1188: douta=16'hd6ba;
1189: douta=16'hbe58;
1190: douta=16'h6bb2;
1191: douta=16'h9493;
1192: douta=16'h84b4;
1193: douta=16'h8c53;
1194: douta=16'hc657;
1195: douta=16'had55;
1196: douta=16'h959a;
1197: douta=16'h4313;
1198: douta=16'h9516;
1199: douta=16'ha534;
1200: douta=16'h9d16;
1201: douta=16'hf7bd;
1202: douta=16'h7496;
1203: douta=16'hfefa;
1204: douta=16'h2a2d;
1205: douta=16'h8433;
1206: douta=16'h9cd5;
1207: douta=16'h9d58;
1208: douta=16'hce59;
1209: douta=16'hadd9;
1210: douta=16'h9558;
1211: douta=16'h42d0;
1212: douta=16'h9494;
1213: douta=16'h3a6f;
1214: douta=16'h6414;
1215: douta=16'hdef9;
1216: douta=16'hc619;
1217: douta=16'hffbb;
1218: douta=16'h63b4;
1219: douta=16'h6c76;
1220: douta=16'h9558;
1221: douta=16'h5bb3;
1222: douta=16'h4b11;
1223: douta=16'h84f7;
1224: douta=16'h94d5;
1225: douta=16'h7476;
1226: douta=16'hb5b9;
1227: douta=16'h853a;
1228: douta=16'h84f7;
1229: douta=16'h9d37;
1230: douta=16'h6c34;
1231: douta=16'ha5fa;
1232: douta=16'h9559;
1233: douta=16'h9558;
1234: douta=16'hbe39;
1235: douta=16'h9538;
1236: douta=16'h7415;
1237: douta=16'h5351;
1238: douta=16'h53d3;
1239: douta=16'h7413;
1240: douta=16'hbe18;
1241: douta=16'had56;
1242: douta=16'h7c75;
1243: douta=16'h8c73;
1244: douta=16'h3aae;
1245: douta=16'h1128;
1246: douta=16'h7455;
1247: douta=16'h9d57;
1248: douta=16'h4312;
1249: douta=16'hb596;
1250: douta=16'h3a2c;
1251: douta=16'h29eb;
1252: douta=16'h3a2c;
1253: douta=16'h9d35;
1254: douta=16'h6b8f;
1255: douta=16'h632e;
1256: douta=16'h83d0;
1257: douta=16'h6b6e;
1258: douta=16'h3aab;
1259: douta=16'h4aab;
1260: douta=16'h8c90;
1261: douta=16'hbd72;
1262: douta=16'hd614;
1263: douta=16'h7411;
1264: douta=16'h426d;
1265: douta=16'h634f;
1266: douta=16'h9513;
1267: douta=16'hded9;
1268: douta=16'h634f;
1269: douta=16'ha514;
1270: douta=16'h6b8f;
1271: douta=16'h63af;
1272: douta=16'h6b8f;
1273: douta=16'ha555;
1274: douta=16'h8c53;
1275: douta=16'h8c73;
1276: douta=16'h39e9;
1277: douta=16'h4a6b;
1278: douta=16'h1128;
1279: douta=16'h6370;
1280: douta=16'h7c32;
1281: douta=16'h6370;
1282: douta=16'h94d4;
1283: douta=16'h52ee;
1284: douta=16'h734f;
1285: douta=16'h5b51;
1286: douta=16'h2a0d;
1287: douta=16'h6390;
1288: douta=16'hc638;
1289: douta=16'h6b90;
1290: douta=16'h6bb1;
1291: douta=16'had35;
1292: douta=16'h18c3;
1293: douta=16'h10e4;
1294: douta=16'h2168;
1295: douta=16'h1106;
1296: douta=16'h218a;
1297: douta=16'ha534;
1298: douta=16'h7c33;
1299: douta=16'h8c94;
1300: douta=16'h7bf0;
1301: douta=16'h634f;
1302: douta=16'h00e6;
1303: douta=16'h21ca;
1304: douta=16'h6c10;
1305: douta=16'h73f1;
1306: douta=16'hbdb6;
1307: douta=16'hb534;
1308: douta=16'h8c94;
1309: douta=16'h6c13;
1310: douta=16'h6bf4;
1311: douta=16'h42cf;
1312: douta=16'ha577;
1313: douta=16'h84b7;
1314: douta=16'h5b93;
1315: douta=16'h2a91;
1316: douta=16'h5372;
1317: douta=16'h114a;
1318: douta=16'h8cf6;
1319: douta=16'h7454;
1320: douta=16'h8c95;
1321: douta=16'h6391;
1322: douta=16'h6458;
1323: douta=16'h5bd5;
1324: douta=16'h32f1;
1325: douta=16'h63f4;
1326: douta=16'h9538;
1327: douta=16'h6499;
1328: douta=16'h2290;
1329: douta=16'h3aaf;
1330: douta=16'h4333;
1331: douta=16'h4352;
1332: douta=16'hce9a;
1333: douta=16'h5bb3;
1334: douta=16'h957b;
1335: douta=16'h4353;
1336: douta=16'h3af2;
1337: douta=16'h32d1;
1338: douta=16'h5c36;
1339: douta=16'h7cd8;
1340: douta=16'h6c36;
1341: douta=16'h5c58;
1342: douta=16'h4b32;
1343: douta=16'h5bd5;
1344: douta=16'h6c78;
1345: douta=16'h53d6;
1346: douta=16'h6478;
1347: douta=16'h4b53;
1348: douta=16'h5b93;
1349: douta=16'h7cb7;
1350: douta=16'h5393;
1351: douta=16'h5311;
1352: douta=16'h63f4;
1353: douta=16'h4af1;
1354: douta=16'h8cb5;
1355: douta=16'h7c96;
1356: douta=16'hc639;
1357: douta=16'hbdd9;
1358: douta=16'h9d16;
1359: douta=16'h7413;
1360: douta=16'h6bf4;
1361: douta=16'h94b4;
1362: douta=16'hc5f8;
1363: douta=16'h9d58;
1364: douta=16'hbdd7;
1365: douta=16'h9d16;
1366: douta=16'had76;
1367: douta=16'h7c34;
1368: douta=16'h9cd4;
1369: douta=16'hbdb6;
1370: douta=16'hc618;
1371: douta=16'hc639;
1372: douta=16'hce5a;
1373: douta=16'hc619;
1374: douta=16'h9d58;
1375: douta=16'h73f1;
1376: douta=16'hadb8;
1377: douta=16'hff9b;
1378: douta=16'hbdf8;
1379: douta=16'he6b9;
1380: douta=16'hb5d8;
1381: douta=16'h5bb2;
1382: douta=16'h6b91;
1383: douta=16'h9d35;
1384: douta=16'hce59;
1385: douta=16'had35;
1386: douta=16'hffdb;
1387: douta=16'h9cb3;
1388: douta=16'h3acf;
1389: douta=16'h52ef;
1390: douta=16'ha555;
1391: douta=16'hde78;
1392: douta=16'had77;
1393: douta=16'hbe39;
1394: douta=16'h6371;
1395: douta=16'h9d16;
1396: douta=16'h6bb2;
1397: douta=16'hc618;
1398: douta=16'hb596;
1399: douta=16'hbe3a;
1400: douta=16'hbdf8;
1401: douta=16'h6c56;
1402: douta=16'h8517;
1403: douta=16'h4b31;
1404: douta=16'h5b70;
1405: douta=16'hbdf7;
1406: douta=16'h9d18;
1407: douta=16'hf77b;
1408: douta=16'hc5d8;
1409: douta=16'hd71c;
1410: douta=16'h63b4;
1411: douta=16'h5372;
1412: douta=16'h8495;
1413: douta=16'h6c55;
1414: douta=16'he6fa;
1415: douta=16'h74b8;
1416: douta=16'h9d98;
1417: douta=16'h3291;
1418: douta=16'h9cb4;
1419: douta=16'h6456;
1420: douta=16'h3af1;
1421: douta=16'h6bd3;
1422: douta=16'h5bb3;
1423: douta=16'h9599;
1424: douta=16'h6457;
1425: douta=16'hd69b;
1426: douta=16'h9d79;
1427: douta=16'h8cf6;
1428: douta=16'h9517;
1429: douta=16'h63b3;
1430: douta=16'h84d6;
1431: douta=16'h9d77;
1432: douta=16'h9d57;
1433: douta=16'h5b10;
1434: douta=16'h5370;
1435: douta=16'ha5d7;
1436: douta=16'h52ee;
1437: douta=16'h94d5;
1438: douta=16'ha557;
1439: douta=16'ha557;
1440: douta=16'h5b2f;
1441: douta=16'h5b0f;
1442: douta=16'h6b90;
1443: douta=16'h532f;
1444: douta=16'h8495;
1445: douta=16'h8cb5;
1446: douta=16'hc658;
1447: douta=16'h8c31;
1448: douta=16'h738e;
1449: douta=16'h0000;
1450: douta=16'h18e3;
1451: douta=16'h0861;
1452: douta=16'h10e3;
1453: douta=16'h5351;
1454: douta=16'h426d;
1455: douta=16'h3a2b;
1456: douta=16'h636f;
1457: douta=16'h3a0a;
1458: douta=16'h7c12;
1459: douta=16'h532f;
1460: douta=16'hb596;
1461: douta=16'h630e;
1462: douta=16'h636f;
1463: douta=16'h3a2a;
1464: douta=16'hc617;
1465: douta=16'hbdb7;
1466: douta=16'h5b51;
1467: douta=16'h73f2;
1468: douta=16'h29a9;
1469: douta=16'h29a8;
1470: douta=16'h532e;
1471: douta=16'hb5b6;
1472: douta=16'h8474;
1473: douta=16'h7bd0;
1474: douta=16'h5b2f;
1475: douta=16'h6bf1;
1476: douta=16'h5bb1;
1477: douta=16'h8c94;
1478: douta=16'h7bf2;
1479: douta=16'h8473;
1480: douta=16'h7454;
1481: douta=16'h2168;
1482: douta=16'h6b8f;
1483: douta=16'h4af0;
1484: douta=16'h2124;
1485: douta=16'h10e4;
1486: douta=16'h39e9;
1487: douta=16'h9494;
1488: douta=16'h738f;
1489: douta=16'h3ab0;
1490: douta=16'h7c33;
1491: douta=16'h3a6e;
1492: douta=16'h4aee;
1493: douta=16'h4acd;
1494: douta=16'hc617;
1495: douta=16'hd615;
1496: douta=16'h5352;
1497: douta=16'h6bb2;
1498: douta=16'h1969;
1499: douta=16'h63d2;
1500: douta=16'h8cb5;
1501: douta=16'h6bd2;
1502: douta=16'h4aee;
1503: douta=16'hc63a;
1504: douta=16'h6c16;
1505: douta=16'h19ac;
1506: douta=16'h29ec;
1507: douta=16'h9516;
1508: douta=16'h9517;
1509: douta=16'hd69a;
1510: douta=16'h84d7;
1511: douta=16'h6416;
1512: douta=16'h4b54;
1513: douta=16'h4394;
1514: douta=16'h5bb3;
1515: douta=16'h4bd5;
1516: douta=16'hb65c;
1517: douta=16'h959a;
1518: douta=16'h7477;
1519: douta=16'h21ac;
1520: douta=16'h2a6f;
1521: douta=16'h222d;
1522: douta=16'h9518;
1523: douta=16'h9518;
1524: douta=16'h5b94;
1525: douta=16'h2a4f;
1526: douta=16'h42f0;
1527: douta=16'h42f0;
1528: douta=16'h9517;
1529: douta=16'h7499;
1530: douta=16'h74b8;
1531: douta=16'h4375;
1532: douta=16'h3313;
1533: douta=16'h1a0d;
1534: douta=16'h9d78;
1535: douta=16'h74d9;
1536: douta=16'h19ee;
1537: douta=16'h32d1;
1538: douta=16'h53f6;
1539: douta=16'h7498;
1540: douta=16'h63f5;
1541: douta=16'h6436;
1542: douta=16'h74b8;
1543: douta=16'h5b50;
1544: douta=16'h7414;
1545: douta=16'ha537;
1546: douta=16'hc61a;
1547: douta=16'hadfb;
1548: douta=16'h7c13;
1549: douta=16'h63b2;
1550: douta=16'h8452;
1551: douta=16'h7c14;
1552: douta=16'h8c95;
1553: douta=16'hce59;
1554: douta=16'h194a;
1555: douta=16'h8cd5;
1556: douta=16'h5352;
1557: douta=16'h9cf5;
1558: douta=16'he6d9;
1559: douta=16'had56;
1560: douta=16'hce18;
1561: douta=16'hb597;
1562: douta=16'h8474;
1563: douta=16'h5b30;
1564: douta=16'hb5d8;
1565: douta=16'hb598;
1566: douta=16'hbdd7;
1567: douta=16'hd65a;
1568: douta=16'h7413;
1569: douta=16'h8c94;
1570: douta=16'h3aaf;
1571: douta=16'h83f2;
1572: douta=16'h9d35;
1573: douta=16'hc5f7;
1574: douta=16'he6ba;
1575: douta=16'hf77b;
1576: douta=16'h7413;
1577: douta=16'h4aee;
1578: douta=16'h83f0;
1579: douta=16'hb596;
1580: douta=16'hbd95;
1581: douta=16'heed8;
1582: douta=16'h9473;
1583: douta=16'had75;
1584: douta=16'h426d;
1585: douta=16'h6bf2;
1586: douta=16'h6370;
1587: douta=16'hf79a;
1588: douta=16'hde79;
1589: douta=16'hb5b7;
1590: douta=16'he71b;
1591: douta=16'hbe19;
1592: douta=16'hbe18;
1593: douta=16'h8cb4;
1594: douta=16'had77;
1595: douta=16'hbdf9;
1596: douta=16'hef1b;
1597: douta=16'hbdf9;
1598: douta=16'h1a0e;
1599: douta=16'h7c33;
1600: douta=16'hbe18;
1601: douta=16'ha5b9;
1602: douta=16'hbe5a;
1603: douta=16'h7476;
1604: douta=16'h95ba;
1605: douta=16'h3b33;
1606: douta=16'h63f3;
1607: douta=16'h4b51;
1608: douta=16'h8495;
1609: douta=16'h8d38;
1610: douta=16'had97;
1611: douta=16'hbe1a;
1612: douta=16'h94d6;
1613: douta=16'h6c96;
1614: douta=16'h6b93;
1615: douta=16'h5b72;
1616: douta=16'h9d78;
1617: douta=16'h5bf5;
1618: douta=16'h9538;
1619: douta=16'hb619;
1620: douta=16'hd6ba;
1621: douta=16'h9d78;
1622: douta=16'h4b74;
1623: douta=16'h8c95;
1624: douta=16'h8c94;
1625: douta=16'h9d36;
1626: douta=16'h9cd6;
1627: douta=16'hb596;
1628: douta=16'h6bd1;
1629: douta=16'h5b10;
1630: douta=16'h7c53;
1631: douta=16'h7c53;
1632: douta=16'ha535;
1633: douta=16'ha576;
1634: douta=16'hb5b8;
1635: douta=16'h7c33;
1636: douta=16'h42ef;
1637: douta=16'h530e;
1638: douta=16'h1106;
1639: douta=16'h426b;
1640: douta=16'h424a;
1641: douta=16'ha536;
1642: douta=16'h2103;
1643: douta=16'h18e3;
1644: douta=16'h10a2;
1645: douta=16'h29a9;
1646: douta=16'h29a8;
1647: douta=16'h73d0;
1648: douta=16'h6b6f;
1649: douta=16'ha4f4;
1650: douta=16'h634f;
1651: douta=16'h632e;
1652: douta=16'h320b;
1653: douta=16'h5b0d;
1654: douta=16'h526a;
1655: douta=16'hbd33;
1656: douta=16'h73b0;
1657: douta=16'h532f;
1658: douta=16'h7c31;
1659: douta=16'h4a8c;
1660: douta=16'ha4f4;
1661: douta=16'hce37;
1662: douta=16'h5b0e;
1663: douta=16'h4ace;
1664: douta=16'h3a2c;
1665: douta=16'h9d14;
1666: douta=16'h9472;
1667: douta=16'ha536;
1668: douta=16'h8c52;
1669: douta=16'h4ace;
1670: douta=16'h5b70;
1671: douta=16'h8c72;
1672: douta=16'h6bd2;
1673: douta=16'hbdd7;
1674: douta=16'h9cf4;
1675: douta=16'h9cf5;
1676: douta=16'h1083;
1677: douta=16'h10e5;
1678: douta=16'h29a9;
1679: douta=16'h7413;
1680: douta=16'h532f;
1681: douta=16'h9cd5;
1682: douta=16'h73f3;
1683: douta=16'h5b70;
1684: douta=16'h5b50;
1685: douta=16'h5350;
1686: douta=16'h0065;
1687: douta=16'h7c31;
1688: douta=16'h94d4;
1689: douta=16'had75;
1690: douta=16'h94d4;
1691: douta=16'h328f;
1692: douta=16'h326d;
1693: douta=16'h6bf3;
1694: douta=16'h42ad;
1695: douta=16'h6b90;
1696: douta=16'h63d3;
1697: douta=16'h9517;
1698: douta=16'hb61a;
1699: douta=16'h3a8f;
1700: douta=16'h6392;
1701: douta=16'h53b4;
1702: douta=16'h4b52;
1703: douta=16'h7436;
1704: douta=16'h84b6;
1705: douta=16'h6c36;
1706: douta=16'h7cda;
1707: douta=16'h8455;
1708: douta=16'h00e9;
1709: douta=16'h2a2d;
1710: douta=16'h5415;
1711: douta=16'hb61a;
1712: douta=16'h84f9;
1713: douta=16'h9539;
1714: douta=16'h6c35;
1715: douta=16'h5b93;
1716: douta=16'h9d38;
1717: douta=16'h5310;
1718: douta=16'h5b52;
1719: douta=16'h2a6f;
1720: douta=16'h2ad2;
1721: douta=16'h118b;
1722: douta=16'h6415;
1723: douta=16'h6459;
1724: douta=16'h5bb5;
1725: douta=16'h853b;
1726: douta=16'h5c36;
1727: douta=16'h3b33;
1728: douta=16'h4b73;
1729: douta=16'h53f6;
1730: douta=16'h4bd5;
1731: douta=16'h32b0;
1732: douta=16'h5b93;
1733: douta=16'h6bf5;
1734: douta=16'h7497;
1735: douta=16'h42cf;
1736: douta=16'h5393;
1737: douta=16'h4b31;
1738: douta=16'had97;
1739: douta=16'ha599;
1740: douta=16'hc5d8;
1741: douta=16'h9d16;
1742: douta=16'h8454;
1743: douta=16'h63b2;
1744: douta=16'h5b6f;
1745: douta=16'hbe19;
1746: douta=16'h73f3;
1747: douta=16'hb5d9;
1748: douta=16'h9d37;
1749: douta=16'h9cf6;
1750: douta=16'hbdd7;
1751: douta=16'hbe17;
1752: douta=16'hbdd8;
1753: douta=16'hc638;
1754: douta=16'hded9;
1755: douta=16'h9d16;
1756: douta=16'h9d37;
1757: douta=16'h9495;
1758: douta=16'h7c53;
1759: douta=16'hb5b7;
1760: douta=16'hb597;
1761: douta=16'he699;
1762: douta=16'h7c13;
1763: douta=16'had35;
1764: douta=16'h94d4;
1765: douta=16'h7c52;
1766: douta=16'hce38;
1767: douta=16'hce78;
1768: douta=16'ha556;
1769: douta=16'h8474;
1770: douta=16'hb575;
1771: douta=16'h7c11;
1772: douta=16'h8432;
1773: douta=16'hc5f6;
1774: douta=16'had33;
1775: douta=16'he6d9;
1776: douta=16'hcdf7;
1777: douta=16'h6bd2;
1778: douta=16'h0908;
1779: douta=16'had75;
1780: douta=16'hce37;
1781: douta=16'hc5f9;
1782: douta=16'heefa;
1783: douta=16'hbdb9;
1784: douta=16'hce7a;
1785: douta=16'h5b71;
1786: douta=16'h63b3;
1787: douta=16'hb5d8;
1788: douta=16'hd6ba;
1789: douta=16'hef3b;
1790: douta=16'h7c56;
1791: douta=16'hce38;
1792: douta=16'h84b7;
1793: douta=16'h7476;
1794: douta=16'h9579;
1795: douta=16'h8454;
1796: douta=16'h959a;
1797: douta=16'h7cb8;
1798: douta=16'hc67a;
1799: douta=16'h5395;
1800: douta=16'h4b10;
1801: douta=16'h5b52;
1802: douta=16'h5351;
1803: douta=16'h63d2;
1804: douta=16'hc65a;
1805: douta=16'ha599;
1806: douta=16'h94b6;
1807: douta=16'h7c56;
1808: douta=16'h8496;
1809: douta=16'h6434;
1810: douta=16'h3ad1;
1811: douta=16'h9517;
1812: douta=16'hb5f9;
1813: douta=16'hadb8;
1814: douta=16'h7456;
1815: douta=16'hdeba;
1816: douta=16'h4a8d;
1817: douta=16'h636f;
1818: douta=16'h42ae;
1819: douta=16'had76;
1820: douta=16'had98;
1821: douta=16'h7c13;
1822: douta=16'h8413;
1823: douta=16'h4aef;
1824: douta=16'h52ce;
1825: douta=16'ha598;
1826: douta=16'h8cb5;
1827: douta=16'h7c95;
1828: douta=16'h7455;
1829: douta=16'hb575;
1830: douta=16'h2a4d;
1831: douta=16'h3a4a;
1832: douta=16'h10e5;
1833: douta=16'h8472;
1834: douta=16'h2924;
1835: douta=16'h1903;
1836: douta=16'h0020;
1837: douta=16'h4a6a;
1838: douta=16'h424a;
1839: douta=16'h29a9;
1840: douta=16'h4aad;
1841: douta=16'had75;
1842: douta=16'h8c94;
1843: douta=16'ha4f3;
1844: douta=16'h62cc;
1845: douta=16'h2188;
1846: douta=16'h7bf0;
1847: douta=16'h94d3;
1848: douta=16'had55;
1849: douta=16'h42ae;
1850: douta=16'h3a2b;
1851: douta=16'h5acd;
1852: douta=16'h42ee;
1853: douta=16'h8472;
1854: douta=16'ha514;
1855: douta=16'h73d1;
1856: douta=16'h7bd0;
1857: douta=16'h4acf;
1858: douta=16'h8431;
1859: douta=16'h73b0;
1860: douta=16'hc5f6;
1861: douta=16'h7bf1;
1862: douta=16'h8433;
1863: douta=16'h5b2f;
1864: douta=16'h6bd1;
1865: douta=16'hb596;
1866: douta=16'h8c94;
1867: douta=16'hbdd7;
1868: douta=16'h0883;
1869: douta=16'h08c4;
1870: douta=16'h1127;
1871: douta=16'h3a6c;
1872: douta=16'h5330;
1873: douta=16'h4b0f;
1874: douta=16'h7c11;
1875: douta=16'h9492;
1876: douta=16'h7bf2;
1877: douta=16'h73f2;
1878: douta=16'h31ec;
1879: douta=16'h21aa;
1880: douta=16'h19ab;
1881: douta=16'h4b51;
1882: douta=16'hce58;
1883: douta=16'h73d2;
1884: douta=16'h63d3;
1885: douta=16'h63b1;
1886: douta=16'h322c;
1887: douta=16'h6390;
1888: douta=16'h2a4e;
1889: douta=16'h9d78;
1890: douta=16'h84f7;
1891: douta=16'h94f7;
1892: douta=16'hc67b;
1893: douta=16'h6436;
1894: douta=16'h32d1;
1895: douta=16'h63f5;
1896: douta=16'h2a8f;
1897: douta=16'h7cf8;
1898: douta=16'h6c56;
1899: douta=16'hb61b;
1900: douta=16'h5b93;
1901: douta=16'h63f4;
1902: douta=16'h2270;
1903: douta=16'h4332;
1904: douta=16'h8d17;
1905: douta=16'h84d8;
1906: douta=16'h7456;
1907: douta=16'h4b52;
1908: douta=16'h5bd3;
1909: douta=16'h73f3;
1910: douta=16'h8495;
1911: douta=16'h7bd2;
1912: douta=16'h3b33;
1913: douta=16'h19cc;
1914: douta=16'h222e;
1915: douta=16'h3b96;
1916: douta=16'h8cd6;
1917: douta=16'h74b7;
1918: douta=16'h7d3b;
1919: douta=16'h6478;
1920: douta=16'h2a90;
1921: douta=16'h5c16;
1922: douta=16'h4332;
1923: douta=16'h3ad1;
1924: douta=16'h6c36;
1925: douta=16'h6c36;
1926: douta=16'h74b9;
1927: douta=16'h63b3;
1928: douta=16'h116a;
1929: douta=16'h5b30;
1930: douta=16'hb577;
1931: douta=16'hce7b;
1932: douta=16'h9d37;
1933: douta=16'h7414;
1934: douta=16'h29eb;
1935: douta=16'h428d;
1936: douta=16'h9d17;
1937: douta=16'hce79;
1938: douta=16'had97;
1939: douta=16'hb5d8;
1940: douta=16'h7414;
1941: douta=16'ha516;
1942: douta=16'h73f1;
1943: douta=16'hbdd7;
1944: douta=16'hbdb6;
1945: douta=16'ha536;
1946: douta=16'hbdf7;
1947: douta=16'h9493;
1948: douta=16'h8cf6;
1949: douta=16'hbd95;
1950: douta=16'hc639;
1951: douta=16'hce59;
1952: douta=16'hce38;
1953: douta=16'hacf5;
1954: douta=16'h6bf1;
1955: douta=16'hde99;
1956: douta=16'h9cd5;
1957: douta=16'h8cd4;
1958: douta=16'hffbc;
1959: douta=16'hef5b;
1960: douta=16'h63b1;
1961: douta=16'h9c73;
1962: douta=16'h9492;
1963: douta=16'h7bef;
1964: douta=16'h9cb3;
1965: douta=16'hde77;
1966: douta=16'ha4f3;
1967: douta=16'h7c12;
1968: douta=16'h9452;
1969: douta=16'h5b91;
1970: douta=16'h5b2f;
1971: douta=16'hce78;
1972: douta=16'hce18;
1973: douta=16'ha5b8;
1974: douta=16'h9473;
1975: douta=16'h7433;
1976: douta=16'ha577;
1977: douta=16'h8c52;
1978: douta=16'hd659;
1979: douta=16'he75c;
1980: douta=16'hae1b;
1981: douta=16'ha599;
1982: douta=16'h6414;
1983: douta=16'h84b5;
1984: douta=16'hd6da;
1985: douta=16'hbe5b;
1986: douta=16'he6fb;
1987: douta=16'hbe1a;
1988: douta=16'h6435;
1989: douta=16'h5bb4;
1990: douta=16'h8473;
1991: douta=16'h3ab0;
1992: douta=16'h2a0e;
1993: douta=16'ha5b8;
1994: douta=16'h84f8;
1995: douta=16'hdeba;
1996: douta=16'hb5d9;
1997: douta=16'h5bf5;
1998: douta=16'h5374;
1999: douta=16'h9d98;
2000: douta=16'h5bb4;
2001: douta=16'h4b10;
2002: douta=16'h8497;
2003: douta=16'hc639;
2004: douta=16'h8d39;
2005: douta=16'h8d18;
2006: douta=16'h42cf;
2007: douta=16'h7454;
2008: douta=16'h422a;
2009: douta=16'h4aad;
2010: douta=16'h8454;
2011: douta=16'hb5b8;
2012: douta=16'h5371;
2013: douta=16'h6330;
2014: douta=16'h8495;
2015: douta=16'h52ee;
2016: douta=16'h8452;
2017: douta=16'hbdf8;
2018: douta=16'h8c73;
2019: douta=16'hb575;
2020: douta=16'h322d;
2021: douta=16'h3a2b;
2022: douta=16'h3a4c;
2023: douta=16'h8cb5;
2024: douta=16'h9d15;
2025: douta=16'h8452;
2026: douta=16'h2925;
2027: douta=16'h2124;
2028: douta=16'h2104;
2029: douta=16'h6b8f;
2030: douta=16'h424a;
2031: douta=16'h5acc;
2032: douta=16'hde37;
2033: douta=16'h7370;
2034: douta=16'h52cd;
2035: douta=16'h39ca;
2036: douta=16'h1948;
2037: douta=16'h73f0;
2038: douta=16'h94b3;
2039: douta=16'h8c11;
2040: douta=16'h6b70;
2041: douta=16'h31a9;
2042: douta=16'h31cb;
2043: douta=16'h00c6;
2044: douta=16'h73f1;
2045: douta=16'hc617;
2046: douta=16'h6c13;
2047: douta=16'h7453;
2048: douta=16'h32ae;
2049: douta=16'h5b90;
2050: douta=16'h19a8;
2051: douta=16'h1147;
2052: douta=16'h0084;
2053: douta=16'h0002;
2054: douta=16'h0002;
2055: douta=16'h0022;
2056: douta=16'h0042;
2057: douta=16'h0042;
2058: douta=16'h0022;
2059: douta=16'h0001;
2060: douta=16'h0063;
2061: douta=16'h0062;
2062: douta=16'h0022;
2063: douta=16'h0002;
2064: douta=16'h0043;
2065: douta=16'h2188;
2066: douta=16'h08e6;
2067: douta=16'h322b;
2068: douta=16'h5371;
2069: douta=16'h7434;
2070: douta=16'hc637;
2071: douta=16'hc596;
2072: douta=16'h5b30;
2073: douta=16'h426d;
2074: douta=16'h19cb;
2075: douta=16'h19cd;
2076: douta=16'h6c34;
2077: douta=16'had97;
2078: douta=16'h9d36;
2079: douta=16'h8494;
2080: douta=16'ha557;
2081: douta=16'h63f4;
2082: douta=16'h7435;
2083: douta=16'h3ab0;
2084: douta=16'h11ac;
2085: douta=16'h32b0;
2086: douta=16'h4bb4;
2087: douta=16'h9d9a;
2088: douta=16'h8cd7;
2089: douta=16'h3af1;
2090: douta=16'h7455;
2091: douta=16'h3b32;
2092: douta=16'h6414;
2093: douta=16'h63f5;
2094: douta=16'hb5d8;
2095: douta=16'h8cf6;
2096: douta=16'h3ad1;
2097: douta=16'h6c35;
2098: douta=16'h3a90;
2099: douta=16'h7456;
2100: douta=16'h7c55;
2101: douta=16'h5b93;
2102: douta=16'h53b4;
2103: douta=16'h1a2e;
2104: douta=16'h4b53;
2105: douta=16'h7c76;
2106: douta=16'h7498;
2107: douta=16'h6c57;
2108: douta=16'h53f6;
2109: douta=16'h4bf7;
2110: douta=16'h3b53;
2111: douta=16'h6cb8;
2112: douta=16'h32b0;
2113: douta=16'h6c77;
2114: douta=16'h6498;
2115: douta=16'h6478;
2116: douta=16'h2a6e;
2117: douta=16'h4352;
2118: douta=16'h4311;
2119: douta=16'h94f6;
2120: douta=16'h8518;
2121: douta=16'h9d58;
2122: douta=16'h42ef;
2123: douta=16'h426e;
2124: douta=16'h42ef;
2125: douta=16'hbdd8;
2126: douta=16'hc5d7;
2127: douta=16'hce5a;
2128: douta=16'h7c54;
2129: douta=16'h8cb4;
2130: douta=16'h8c74;
2131: douta=16'h7bf3;
2132: douta=16'h6bd2;
2133: douta=16'h94b5;
2134: douta=16'had37;
2135: douta=16'hbe38;
2136: douta=16'had57;
2137: douta=16'h7454;
2138: douta=16'h5b30;
2139: douta=16'h9cf5;
2140: douta=16'hadb8;
2141: douta=16'hf75a;
2142: douta=16'he6db;
2143: douta=16'h9d15;
2144: douta=16'h9493;
2145: douta=16'hc617;
2146: douta=16'hbd75;
2147: douta=16'hdeb9;
2148: douta=16'hce59;
2149: douta=16'h7476;
2150: douta=16'h8c11;
2151: douta=16'h94d2;
2152: douta=16'ha534;
2153: douta=16'h8c30;
2154: douta=16'hff7b;
2155: douta=16'hf75b;
2156: douta=16'h83f2;
2157: douta=16'h94b3;
2158: douta=16'h8c92;
2159: douta=16'h8451;
2160: douta=16'hb596;
2161: douta=16'hb576;
2162: douta=16'hd657;
2163: douta=16'h8493;
2164: douta=16'h73b0;
2165: douta=16'h4350;
2166: douta=16'h84b5;
2167: douta=16'hff9c;
2168: douta=16'h9d98;
2169: douta=16'hbd75;
2170: douta=16'h328f;
2171: douta=16'h9517;
2172: douta=16'h6c76;
2173: douta=16'ha5d9;
2174: douta=16'hd67a;
2175: douta=16'h9578;
2176: douta=16'h6cd9;
2177: douta=16'h32f3;
2178: douta=16'hce9a;
2179: douta=16'h9537;
2180: douta=16'h84d7;
2181: douta=16'h84b6;
2182: douta=16'hd6dc;
2183: douta=16'hce7b;
2184: douta=16'h5373;
2185: douta=16'hb5f9;
2186: douta=16'h6c77;
2187: douta=16'h5b72;
2188: douta=16'h8cb5;
2189: douta=16'h8495;
2190: douta=16'hdefa;
2191: douta=16'hd679;
2192: douta=16'hbe9c;
2193: douta=16'h8d39;
2194: douta=16'ha557;
2195: douta=16'hbe5b;
2196: douta=16'ha5da;
2197: douta=16'h5373;
2198: douta=16'hc639;
2199: douta=16'h7455;
2200: douta=16'hb5d7;
2201: douta=16'h6bd2;
2202: douta=16'had34;
2203: douta=16'h42ae;
2204: douta=16'h6391;
2205: douta=16'h8d17;
2206: douta=16'h5b30;
2207: douta=16'hd5f8;
2208: douta=16'h4aae;
2209: douta=16'h630e;
2210: douta=16'h8473;
2211: douta=16'hb619;
2212: douta=16'hd658;
2213: douta=16'h5b70;
2214: douta=16'h9c72;
2215: douta=16'h2167;
2216: douta=16'h1926;
2217: douta=16'h1926;
2218: douta=16'h5acb;
2219: douta=16'h2124;
2220: douta=16'h20e4;
2221: douta=16'had75;
2222: douta=16'h5b0e;
2223: douta=16'hb554;
2224: douta=16'h5b0e;
2225: douta=16'h634e;
2226: douta=16'h5b4e;
2227: douta=16'ha534;
2228: douta=16'h9492;
2229: douta=16'h9430;
2230: douta=16'h634f;
2231: douta=16'h8cb3;
2232: douta=16'h4aad;
2233: douta=16'hb5f6;
2234: douta=16'h6370;
2235: douta=16'h73f2;
2236: douta=16'h428c;
2237: douta=16'h1127;
2238: douta=16'h0083;
2239: douta=16'h0842;
2240: douta=16'h0863;
2241: douta=16'h0063;
2242: douta=16'h08a4;
2243: douta=16'h08a4;
2244: douta=16'h08a4;
2245: douta=16'h0884;
2246: douta=16'h10c4;
2247: douta=16'h08a4;
2248: douta=16'h08c4;
2249: douta=16'h0884;
2250: douta=16'h0884;
2251: douta=16'h08a4;
2252: douta=16'h0883;
2253: douta=16'h0883;
2254: douta=16'h0063;
2255: douta=16'h0863;
2256: douta=16'h0863;
2257: douta=16'h0883;
2258: douta=16'h0062;
2259: douta=16'h0062;
2260: douta=16'h0021;
2261: douta=16'h0001;
2262: douta=16'h0022;
2263: douta=16'h1167;
2264: douta=16'h42ad;
2265: douta=16'h9d34;
2266: douta=16'hc63a;
2267: douta=16'h6436;
2268: douta=16'h6371;
2269: douta=16'h322d;
2270: douta=16'h2a2d;
2271: douta=16'h9d36;
2272: douta=16'h7c74;
2273: douta=16'hd67a;
2274: douta=16'h7c55;
2275: douta=16'h7498;
2276: douta=16'h3af2;
2277: douta=16'h2a4f;
2278: douta=16'h32af;
2279: douta=16'h222e;
2280: douta=16'h4b53;
2281: douta=16'h63f4;
2282: douta=16'h7476;
2283: douta=16'hb5ba;
2284: douta=16'h5351;
2285: douta=16'h5351;
2286: douta=16'h326e;
2287: douta=16'h5352;
2288: douta=16'h9517;
2289: douta=16'ha578;
2290: douta=16'h7498;
2291: douta=16'h32f1;
2292: douta=16'h4b31;
2293: douta=16'h8cd6;
2294: douta=16'h6416;
2295: douta=16'h6c14;
2296: douta=16'h5bf6;
2297: douta=16'h3b13;
2298: douta=16'h3b32;
2299: douta=16'h8518;
2300: douta=16'h959c;
2301: douta=16'h5c38;
2302: douta=16'h74da;
2303: douta=16'h2ad2;
2304: douta=16'h1a0d;
2305: douta=16'h7478;
2306: douta=16'h53f5;
2307: douta=16'h74d9;
2308: douta=16'h5b93;
2309: douta=16'h328f;
2310: douta=16'h6c56;
2311: douta=16'h6bb2;
2312: douta=16'h7c34;
2313: douta=16'h8c94;
2314: douta=16'h94d5;
2315: douta=16'ha557;
2316: douta=16'h5bd3;
2317: douta=16'h5351;
2318: douta=16'h73d1;
2319: douta=16'h7413;
2320: douta=16'hadd9;
2321: douta=16'hd679;
2322: douta=16'hb597;
2323: douta=16'had97;
2324: douta=16'ha577;
2325: douta=16'h8453;
2326: douta=16'h6b91;
2327: douta=16'had96;
2328: douta=16'hb5b8;
2329: douta=16'hb5b8;
2330: douta=16'ha516;
2331: douta=16'h73d2;
2332: douta=16'h8cb6;
2333: douta=16'hce38;
2334: douta=16'hdeb9;
2335: douta=16'hc639;
2336: douta=16'hc617;
2337: douta=16'hb555;
2338: douta=16'h7c12;
2339: douta=16'hb5b6;
2340: douta=16'hd6b9;
2341: douta=16'h8cd5;
2342: douta=16'he6d9;
2343: douta=16'hc637;
2344: douta=16'h5350;
2345: douta=16'h42ad;
2346: douta=16'hb594;
2347: douta=16'hbdd6;
2348: douta=16'hd658;
2349: douta=16'hbd96;
2350: douta=16'h7390;
2351: douta=16'h8cd4;
2352: douta=16'h6b0e;
2353: douta=16'hb533;
2354: douta=16'hffba;
2355: douta=16'h9cd4;
2356: douta=16'hbdd6;
2357: douta=16'h42cf;
2358: douta=16'h6b50;
2359: douta=16'h9d56;
2360: douta=16'h9516;
2361: douta=16'he6d8;
2362: douta=16'h8cb5;
2363: douta=16'hd71c;
2364: douta=16'h859a;
2365: douta=16'h6c55;
2366: douta=16'h63d3;
2367: douta=16'h94d5;
2368: douta=16'h9518;
2369: douta=16'h9538;
2370: douta=16'hce9b;
2371: douta=16'h9d38;
2372: douta=16'h6c35;
2373: douta=16'h84d6;
2374: douta=16'h84b6;
2375: douta=16'h7c75;
2376: douta=16'h8d18;
2377: douta=16'hbe5a;
2378: douta=16'h6477;
2379: douta=16'h84b6;
2380: douta=16'h6bf2;
2381: douta=16'h7413;
2382: douta=16'h8517;
2383: douta=16'hbe5a;
2384: douta=16'h957a;
2385: douta=16'hbe3b;
2386: douta=16'h7c56;
2387: douta=16'h8d59;
2388: douta=16'h6bf5;
2389: douta=16'h32b0;
2390: douta=16'h63d2;
2391: douta=16'h63d2;
2392: douta=16'h8cb4;
2393: douta=16'h8cb5;
2394: douta=16'hde98;
2395: douta=16'h84d6;
2396: douta=16'h3a0c;
2397: douta=16'h530f;
2398: douta=16'h6391;
2399: douta=16'h94d4;
2400: douta=16'h9d15;
2401: douta=16'had54;
2402: douta=16'h6b90;
2403: douta=16'h6bf2;
2404: douta=16'h94d4;
2405: douta=16'h7454;
2406: douta=16'hf73b;
2407: douta=16'h63d2;
2408: douta=16'h8453;
2409: douta=16'h3189;
2410: douta=16'h3167;
2411: douta=16'h2924;
2412: douta=16'h20e3;
2413: douta=16'h6b8f;
2414: douta=16'h7bd0;
2415: douta=16'hbdd6;
2416: douta=16'ha533;
2417: douta=16'h2988;
2418: douta=16'h632e;
2419: douta=16'h31c8;
2420: douta=16'h8c92;
2421: douta=16'hb574;
2422: douta=16'ha556;
2423: douta=16'ha577;
2424: douta=16'h3a4c;
2425: douta=16'h3acc;
2426: douta=16'h2168;
2427: douta=16'h1126;
2428: douta=16'h0002;
2429: douta=16'h0042;
2430: douta=16'h0883;
2431: douta=16'h08a4;
2432: douta=16'h08a4;
2433: douta=16'h10c5;
2434: douta=16'h0884;
2435: douta=16'h08a4;
2436: douta=16'h08c4;
2437: douta=16'h08a4;
2438: douta=16'h08a4;
2439: douta=16'h0884;
2440: douta=16'h08a4;
2441: douta=16'h08a4;
2442: douta=16'h08a4;
2443: douta=16'h0884;
2444: douta=16'h0884;
2445: douta=16'h0884;
2446: douta=16'h0883;
2447: douta=16'h0883;
2448: douta=16'h0883;
2449: douta=16'h0883;
2450: douta=16'h0883;
2451: douta=16'h0883;
2452: douta=16'h0883;
2453: douta=16'h08a4;
2454: douta=16'h0843;
2455: douta=16'h0001;
2456: douta=16'h0002;
2457: douta=16'h0063;
2458: douta=16'h63f1;
2459: douta=16'h53b5;
2460: douta=16'had98;
2461: douta=16'h7414;
2462: douta=16'h4b31;
2463: douta=16'h3a8e;
2464: douta=16'h3a8e;
2465: douta=16'h7474;
2466: douta=16'h7cb7;
2467: douta=16'h84b8;
2468: douta=16'h6415;
2469: douta=16'h4394;
2470: douta=16'h7cf9;
2471: douta=16'h3ab0;
2472: douta=16'h4311;
2473: douta=16'h3ad0;
2474: douta=16'h3ad0;
2475: douta=16'h6c35;
2476: douta=16'h8cb6;
2477: douta=16'h9559;
2478: douta=16'h7414;
2479: douta=16'h6bf4;
2480: douta=16'h5bb3;
2481: douta=16'h7cb6;
2482: douta=16'h5bd4;
2483: douta=16'h7c96;
2484: douta=16'h5bd3;
2485: douta=16'h5bb4;
2486: douta=16'h114a;
2487: douta=16'h4310;
2488: douta=16'h9579;
2489: douta=16'h5417;
2490: douta=16'h63f5;
2491: douta=16'h0a0e;
2492: douta=16'h3b53;
2493: douta=16'h3b54;
2494: douta=16'h74da;
2495: douta=16'h853a;
2496: douta=16'h32f2;
2497: douta=16'h6436;
2498: douta=16'h6437;
2499: douta=16'h6c98;
2500: douta=16'h21ac;
2501: douta=16'h5393;
2502: douta=16'h4b32;
2503: douta=16'h4aef;
2504: douta=16'h9d58;
2505: douta=16'h7c75;
2506: douta=16'h5b72;
2507: douta=16'h6bd2;
2508: douta=16'h5393;
2509: douta=16'h8476;
2510: douta=16'hb5b8;
2511: douta=16'ha577;
2512: douta=16'hbe3a;
2513: douta=16'had77;
2514: douta=16'h5b2f;
2515: douta=16'h73f2;
2516: douta=16'h7c74;
2517: douta=16'ha536;
2518: douta=16'ha536;
2519: douta=16'hbdf7;
2520: douta=16'hc5f7;
2521: douta=16'ha577;
2522: douta=16'h7c33;
2523: douta=16'h5b51;
2524: douta=16'h9d57;
2525: douta=16'heefa;
2526: douta=16'hdeb9;
2527: douta=16'h94f5;
2528: douta=16'ha514;
2529: douta=16'ha4f4;
2530: douta=16'h9cb4;
2531: douta=16'he719;
2532: douta=16'hb576;
2533: douta=16'h5b71;
2534: douta=16'hcdf5;
2535: douta=16'hbdd7;
2536: douta=16'h7c52;
2537: douta=16'ha4d3;
2538: douta=16'hef19;
2539: douta=16'hce77;
2540: douta=16'hc5d6;
2541: douta=16'hce77;
2542: douta=16'h0085;
2543: douta=16'h532e;
2544: douta=16'hbdd5;
2545: douta=16'hcdb5;
2546: douta=16'hff19;
2547: douta=16'h4b0f;
2548: douta=16'hb556;
2549: douta=16'h39ea;
2550: douta=16'had13;
2551: douta=16'hd6b9;
2552: douta=16'h9536;
2553: douta=16'hff9b;
2554: douta=16'h6371;
2555: douta=16'h7c95;
2556: douta=16'h42d0;
2557: douta=16'h5351;
2558: douta=16'hb5b7;
2559: douta=16'hc659;
2560: douta=16'h5394;
2561: douta=16'h5b93;
2562: douta=16'h6c14;
2563: douta=16'h4331;
2564: douta=16'h8495;
2565: douta=16'h84f7;
2566: douta=16'h9d99;
2567: douta=16'h7cd7;
2568: douta=16'h8d17;
2569: douta=16'h64d9;
2570: douta=16'h3a2f;
2571: douta=16'h5bd3;
2572: douta=16'h6bf3;
2573: douta=16'hbe1a;
2574: douta=16'h8d18;
2575: douta=16'hcedc;
2576: douta=16'h9579;
2577: douta=16'h74b8;
2578: douta=16'hce59;
2579: douta=16'h8d18;
2580: douta=16'h4310;
2581: douta=16'h5332;
2582: douta=16'ha576;
2583: douta=16'h94b5;
2584: douta=16'h7414;
2585: douta=16'h9452;
2586: douta=16'h9537;
2587: douta=16'h42cf;
2588: douta=16'h5b2f;
2589: douta=16'h6b90;
2590: douta=16'ha576;
2591: douta=16'h73f3;
2592: douta=16'h8cb4;
2593: douta=16'h5b2f;
2594: douta=16'h94d5;
2595: douta=16'h532f;
2596: douta=16'hb5f7;
2597: douta=16'hde99;
2598: douta=16'h6391;
2599: douta=16'h6371;
2600: douta=16'h29ea;
2601: douta=16'h6370;
2602: douta=16'h5b2f;
2603: douta=16'h3986;
2604: douta=16'h18e3;
2605: douta=16'h528c;
2606: douta=16'ha4d4;
2607: douta=16'h422b;
2608: douta=16'h3a4b;
2609: douta=16'h4aac;
2610: douta=16'h7c72;
2611: douta=16'h8cb2;
2612: douta=16'h29c8;
2613: douta=16'h0083;
2614: douta=16'h08a4;
2615: douta=16'h10a4;
2616: douta=16'h10a4;
2617: douta=16'h10e4;
2618: douta=16'h10c5;
2619: douta=16'h10a5;
2620: douta=16'h08a4;
2621: douta=16'h08a4;
2622: douta=16'h0883;
2623: douta=16'h0062;
2624: douta=16'h0042;
2625: douta=16'h10a4;
2626: douta=16'h2168;
2627: douta=16'h29a9;
2628: douta=16'h31ca;
2629: douta=16'h3a4c;
2630: douta=16'h3a6c;
2631: douta=16'h4aef;
2632: douta=16'h4aaf;
2633: douta=16'h428f;
2634: douta=16'h428f;
2635: douta=16'h42ae;
2636: douta=16'h426d;
2637: douta=16'h3a2c;
2638: douta=16'h3a2b;
2639: douta=16'h320b;
2640: douta=16'h31ca;
2641: douta=16'h29a9;
2642: douta=16'h1926;
2643: douta=16'h10e5;
2644: douta=16'h0062;
2645: douta=16'h0041;
2646: douta=16'h0882;
2647: douta=16'h0884;
2648: douta=16'h08c3;
2649: douta=16'h08a3;
2650: douta=16'h08a4;
2651: douta=16'h08a4;
2652: douta=16'h0883;
2653: douta=16'h0000;
2654: douta=16'h0000;
2655: douta=16'h21ea;
2656: douta=16'h8518;
2657: douta=16'h4b30;
2658: douta=16'h94f6;
2659: douta=16'h19ac;
2660: douta=16'h19cd;
2661: douta=16'h2a90;
2662: douta=16'h7475;
2663: douta=16'h3b11;
2664: douta=16'h6c14;
2665: douta=16'h5352;
2666: douta=16'h63f4;
2667: douta=16'h324e;
2668: douta=16'h3a6e;
2669: douta=16'h4b2f;
2670: douta=16'h21ec;
2671: douta=16'h6c34;
2672: douta=16'h9d79;
2673: douta=16'h9d79;
2674: douta=16'h3ad0;
2675: douta=16'h224f;
2676: douta=16'h4b32;
2677: douta=16'h63d3;
2678: douta=16'h4b53;
2679: douta=16'h4b73;
2680: douta=16'h2250;
2681: douta=16'h3312;
2682: douta=16'h6c56;
2683: douta=16'h6cdb;
2684: douta=16'h6c57;
2685: douta=16'h6cdb;
2686: douta=16'h5c58;
2687: douta=16'h1a0e;
2688: douta=16'h7d5c;
2689: douta=16'h6c57;
2690: douta=16'h3af1;
2691: douta=16'h4332;
2692: douta=16'h6c35;
2693: douta=16'h84f9;
2694: douta=16'h74b7;
2695: douta=16'h8495;
2696: douta=16'h5331;
2697: douta=16'h4b30;
2698: douta=16'h5330;
2699: douta=16'h6350;
2700: douta=16'h9d37;
2701: douta=16'h84d7;
2702: douta=16'ha555;
2703: douta=16'h94d5;
2704: douta=16'h8454;
2705: douta=16'h7413;
2706: douta=16'h8c73;
2707: douta=16'hb597;
2708: douta=16'ha576;
2709: douta=16'hde99;
2710: douta=16'h9cf5;
2711: douta=16'h9516;
2712: douta=16'h6bb2;
2713: douta=16'ha4f4;
2714: douta=16'h9cf3;
2715: douta=16'hbdd8;
2716: douta=16'h94d5;
2717: douta=16'hd699;
2718: douta=16'h94f4;
2719: douta=16'hb5d7;
2720: douta=16'ha514;
2721: douta=16'hb595;
2722: douta=16'hce38;
2723: douta=16'hded9;
2724: douta=16'had55;
2725: douta=16'h4ace;
2726: douta=16'hce16;
2727: douta=16'hc5f6;
2728: douta=16'h9d15;
2729: douta=16'h8411;
2730: douta=16'hbdb5;
2731: douta=16'h3aae;
2732: douta=16'hc5d4;
2733: douta=16'he6d8;
2734: douta=16'hd617;
2735: douta=16'h8431;
2736: douta=16'heeb8;
2737: douta=16'h9471;
2738: douta=16'h94b2;
2739: douta=16'h5b0b;
2740: douta=16'hf77a;
2741: douta=16'hbd75;
2742: douta=16'hfffc;
2743: douta=16'ha514;
2744: douta=16'h4b50;
2745: douta=16'h8452;
2746: douta=16'hbdf8;
2747: douta=16'ha5b8;
2748: douta=16'h8475;
2749: douta=16'h7474;
2750: douta=16'hb577;
2751: douta=16'h52ce;
2752: douta=16'h9537;
2753: douta=16'hb63b;
2754: douta=16'h9579;
2755: douta=16'hae1a;
2756: douta=16'h7497;
2757: douta=16'h94f6;
2758: douta=16'h3a8f;
2759: douta=16'h32b0;
2760: douta=16'h6c14;
2761: douta=16'h63f4;
2762: douta=16'h9578;
2763: douta=16'h6c56;
2764: douta=16'h7476;
2765: douta=16'ha61b;
2766: douta=16'h53d4;
2767: douta=16'h5b93;
2768: douta=16'h7c96;
2769: douta=16'h2a6f;
2770: douta=16'hc65a;
2771: douta=16'h8518;
2772: douta=16'h957a;
2773: douta=16'h9cd6;
2774: douta=16'hadfa;
2775: douta=16'ha556;
2776: douta=16'h3a4c;
2777: douta=16'h9cd3;
2778: douta=16'h5350;
2779: douta=16'h42f0;
2780: douta=16'h8d37;
2781: douta=16'h9d16;
2782: douta=16'hbdd8;
2783: douta=16'h5330;
2784: douta=16'h73b0;
2785: douta=16'h7413;
2786: douta=16'h8d77;
2787: douta=16'h84d6;
2788: douta=16'h7413;
2789: douta=16'h7cb5;
2790: douta=16'h6bf2;
2791: douta=16'h9d56;
2792: douta=16'h5b72;
2793: douta=16'hbe5b;
2794: douta=16'h6bd1;
2795: douta=16'h6b4d;
2796: douta=16'h20e4;
2797: douta=16'h2145;
2798: douta=16'h5b0d;
2799: douta=16'h9d34;
2800: douta=16'h7411;
2801: douta=16'h4aac;
2802: douta=16'h10c5;
2803: douta=16'h0884;
2804: douta=16'h10e4;
2805: douta=16'h10c4;
2806: douta=16'h10c5;
2807: douta=16'h10e5;
2808: douta=16'h10e4;
2809: douta=16'h0063;
2810: douta=16'h0862;
2811: douta=16'h1084;
2812: douta=16'h29c9;
2813: douta=16'h3a2b;
2814: douta=16'h4a8e;
2815: douta=16'h4ace;
2816: douta=16'h5b72;
2817: douta=16'h4b51;
2818: douta=16'h6415;
2819: douta=16'h63f6;
2820: douta=16'h6c56;
2821: douta=16'h6415;
2822: douta=16'h6c57;
2823: douta=16'h6c57;
2824: douta=16'h74d9;
2825: douta=16'h6c98;
2826: douta=16'h7d1a;
2827: douta=16'h7d1a;
2828: douta=16'h7cf9;
2829: douta=16'h853a;
2830: douta=16'h6456;
2831: douta=16'h6c57;
2832: douta=16'h6416;
2833: douta=16'h63f5;
2834: douta=16'h5b93;
2835: douta=16'h5372;
2836: douta=16'h426e;
2837: douta=16'h322d;
2838: douta=16'h3aae;
2839: douta=16'h21a9;
2840: douta=16'h10e5;
2841: douta=16'h1084;
2842: douta=16'h0042;
2843: douta=16'h0883;
2844: douta=16'h08a3;
2845: douta=16'h08a4;
2846: douta=16'h08c4;
2847: douta=16'h08a4;
2848: douta=16'h0001;
2849: douta=16'h29e9;
2850: douta=16'h42cf;
2851: douta=16'h6415;
2852: douta=16'h6c54;
2853: douta=16'h9538;
2854: douta=16'h6415;
2855: douta=16'h1128;
2856: douta=16'h42d1;
2857: douta=16'h42ce;
2858: douta=16'h63f3;
2859: douta=16'had56;
2860: douta=16'h7c34;
2861: douta=16'h5b72;
2862: douta=16'h3a6f;
2863: douta=16'h3ad0;
2864: douta=16'h116a;
2865: douta=16'h4310;
2866: douta=16'h6c34;
2867: douta=16'h7455;
2868: douta=16'h5bf5;
2869: douta=16'h222e;
2870: douta=16'h5b92;
2871: douta=16'h7455;
2872: douta=16'h8cd6;
2873: douta=16'h5c58;
2874: douta=16'h7d1a;
2875: douta=16'h5bf6;
2876: douta=16'h6cb9;
2877: douta=16'h3b33;
2878: douta=16'h6458;
2879: douta=16'h959b;
2880: douta=16'h6478;
2881: douta=16'h6c36;
2882: douta=16'h5c16;
2883: douta=16'h4312;
2884: douta=16'h5371;
2885: douta=16'h3a8e;
2886: douta=16'h84d8;
2887: douta=16'h8d17;
2888: douta=16'h8495;
2889: douta=16'h6bf4;
2890: douta=16'h428d;
2891: douta=16'h6370;
2892: douta=16'h5351;
2893: douta=16'h8497;
2894: douta=16'hdeba;
2895: douta=16'hbe19;
2896: douta=16'hc67a;
2897: douta=16'h8454;
2898: douta=16'h9452;
2899: douta=16'h42d0;
2900: douta=16'h32ae;
2901: douta=16'h94f5;
2902: douta=16'hc5f8;
2903: douta=16'hc639;
2904: douta=16'hb577;
2905: douta=16'h8453;
2906: douta=16'h73d1;
2907: douta=16'h94d5;
2908: douta=16'hce37;
2909: douta=16'hef5b;
2910: douta=16'hd679;
2911: douta=16'ha556;
2912: douta=16'ha535;
2913: douta=16'h9473;
2914: douta=16'hce38;
2915: douta=16'hef1a;
2916: douta=16'hde78;
2917: douta=16'h6391;
2918: douta=16'had13;
2919: douta=16'h8cb3;
2920: douta=16'hb574;
2921: douta=16'hce15;
2922: douta=16'hd678;
2923: douta=16'h9d35;
2924: douta=16'h734e;
2925: douta=16'h9c70;
2926: douta=16'h52a9;
2927: douta=16'hc5f4;
2928: douta=16'hf75a;
2929: douta=16'hc5d4;
2930: douta=16'h5aed;
2931: douta=16'h5aeb;
2932: douta=16'hbdd5;
2933: douta=16'h73af;
2934: douta=16'hbdd5;
2935: douta=16'hdeb9;
2936: douta=16'h6c34;
2937: douta=16'hbdb6;
2938: douta=16'h8493;
2939: douta=16'h84d5;
2940: douta=16'h6390;
2941: douta=16'h9d56;
2942: douta=16'he71a;
2943: douta=16'ha4f5;
2944: douta=16'h3b11;
2945: douta=16'h5373;
2946: douta=16'h8517;
2947: douta=16'h9db9;
2948: douta=16'h6c56;
2949: douta=16'hce7b;
2950: douta=16'h7c75;
2951: douta=16'h4b73;
2952: douta=16'h9d37;
2953: douta=16'h222d;
2954: douta=16'h42d0;
2955: douta=16'h7455;
2956: douta=16'h7455;
2957: douta=16'ha61b;
2958: douta=16'h6c98;
2959: douta=16'h8d19;
2960: douta=16'h9d99;
2961: douta=16'h222f;
2962: douta=16'h7cd7;
2963: douta=16'h42f0;
2964: douta=16'h7476;
2965: douta=16'h94d6;
2966: douta=16'h9d77;
2967: douta=16'ha558;
2968: douta=16'h73f2;
2969: douta=16'hc5f7;
2970: douta=16'h3a2c;
2971: douta=16'h320d;
2972: douta=16'h326d;
2973: douta=16'h6bf2;
2974: douta=16'h9d56;
2975: douta=16'h6c13;
2976: douta=16'hd679;
2977: douta=16'h8494;
2978: douta=16'h6c14;
2979: douta=16'h5330;
2980: douta=16'h8cd5;
2981: douta=16'h9537;
2982: douta=16'h4b2f;
2983: douta=16'h4acf;
2984: douta=16'h31ca;
2985: douta=16'h5b71;
2986: douta=16'h9d15;
2987: douta=16'h8431;
2988: douta=16'h2925;
2989: douta=16'h18e4;
2990: douta=16'h426b;
2991: douta=16'h638f;
2992: douta=16'h2167;
2993: douta=16'h0042;
2994: douta=16'h10a4;
2995: douta=16'h10a5;
2996: douta=16'h10e5;
2997: douta=16'h10e5;
2998: douta=16'h10c4;
2999: douta=16'h0884;
3000: douta=16'h0843;
3001: douta=16'h2988;
3002: douta=16'h39eb;
3003: douta=16'h426c;
3004: douta=16'h5310;
3005: douta=16'h5332;
3006: douta=16'h63d4;
3007: douta=16'h6c15;
3008: douta=16'h63d4;
3009: douta=16'h74d9;
3010: douta=16'h74fa;
3011: douta=16'h7d1b;
3012: douta=16'h74b9;
3013: douta=16'h5c37;
3014: douta=16'h6c98;
3015: douta=16'h6c78;
3016: douta=16'h6cb9;
3017: douta=16'h6457;
3018: douta=16'h6c77;
3019: douta=16'h8d5b;
3020: douta=16'h7d1a;
3021: douta=16'h7d1a;
3022: douta=16'h5bf6;
3023: douta=16'h6437;
3024: douta=16'h6cb9;
3025: douta=16'h753b;
3026: douta=16'h7cfa;
3027: douta=16'h74f9;
3028: douta=16'h6c56;
3029: douta=16'h4b52;
3030: douta=16'h5bb4;
3031: douta=16'h4310;
3032: douta=16'h3a4c;
3033: douta=16'h29ca;
3034: douta=16'h2147;
3035: douta=16'h0042;
3036: douta=16'h0062;
3037: douta=16'h1084;
3038: douta=16'h08c4;
3039: douta=16'h08a4;
3040: douta=16'h10a4;
3041: douta=16'h0002;
3042: douta=16'h0001;
3043: douta=16'h3af0;
3044: douta=16'h6c54;
3045: douta=16'h9d99;
3046: douta=16'h63f5;
3047: douta=16'h8473;
3048: douta=16'h7c76;
3049: douta=16'h0149;
3050: douta=16'h328f;
3051: douta=16'h5b92;
3052: douta=16'h8cb5;
3053: douta=16'h4b11;
3054: douta=16'ha557;
3055: douta=16'h4b31;
3056: douta=16'h21ab;
3057: douta=16'h21aa;
3058: douta=16'h6c14;
3059: douta=16'h8cf6;
3060: douta=16'h7477;
3061: douta=16'h3af1;
3062: douta=16'h3ad1;
3063: douta=16'h4352;
3064: douta=16'h9d9a;
3065: douta=16'h6cb8;
3066: douta=16'h9e1d;
3067: douta=16'h74fa;
3068: douta=16'h4b96;
3069: douta=16'h4375;
3070: douta=16'h4374;
3071: douta=16'h74b8;
3072: douta=16'h74fa;
3073: douta=16'h6c78;
3074: douta=16'h7d1a;
3075: douta=16'h4b95;
3076: douta=16'h5bb4;
3077: douta=16'h5331;
3078: douta=16'h63b3;
3079: douta=16'h7456;
3080: douta=16'h6371;
3081: douta=16'h5b72;
3082: douta=16'h42ae;
3083: douta=16'h7c34;
3084: douta=16'hb5b8;
3085: douta=16'h9538;
3086: douta=16'hb576;
3087: douta=16'ha577;
3088: douta=16'h8454;
3089: douta=16'h5b0f;
3090: douta=16'h7bf2;
3091: douta=16'hb597;
3092: douta=16'h9d56;
3093: douta=16'hb5d8;
3094: douta=16'hbdd8;
3095: douta=16'h8c95;
3096: douta=16'hbd76;
3097: douta=16'ha576;
3098: douta=16'h7c53;
3099: douta=16'hbdb7;
3100: douta=16'hd6ba;
3101: douta=16'he657;
3102: douta=16'hb65a;
3103: douta=16'h7c53;
3104: douta=16'h8432;
3105: douta=16'hc616;
3106: douta=16'hd617;
3107: douta=16'hd698;
3108: douta=16'had34;
3109: douta=16'h3a8d;
3110: douta=16'hc616;
3111: douta=16'ha514;
3112: douta=16'had33;
3113: douta=16'hde57;
3114: douta=16'h6bcf;
3115: douta=16'h6bf0;
3116: douta=16'hb512;
3117: douta=16'hbdd4;
3118: douta=16'hde57;
3119: douta=16'h8c71;
3120: douta=16'hce57;
3121: douta=16'h9491;
3122: douta=16'h8c71;
3123: douta=16'h6b4b;
3124: douta=16'hce76;
3125: douta=16'h9c0f;
3126: douta=16'he6d7;
3127: douta=16'ha576;
3128: douta=16'h6bb1;
3129: douta=16'h6bd1;
3130: douta=16'hd637;
3131: douta=16'h6413;
3132: douta=16'h8c52;
3133: douta=16'h5372;
3134: douta=16'hdeba;
3135: douta=16'h52cd;
3136: douta=16'h3acf;
3137: douta=16'h9d16;
3138: douta=16'h5bb2;
3139: douta=16'hae3b;
3140: douta=16'h9cd7;
3141: douta=16'hd6dc;
3142: douta=16'had98;
3143: douta=16'h220e;
3144: douta=16'h7c34;
3145: douta=16'h5c15;
3146: douta=16'h32d2;
3147: douta=16'h8d38;
3148: douta=16'h9518;
3149: douta=16'h859b;
3150: douta=16'h4bf6;
3151: douta=16'h6c56;
3152: douta=16'h5bb4;
3153: douta=16'h84b8;
3154: douta=16'h5415;
3155: douta=16'h6c76;
3156: douta=16'h5bf5;
3157: douta=16'h94f6;
3158: douta=16'h5b92;
3159: douta=16'h6c76;
3160: douta=16'h632f;
3161: douta=16'h9d15;
3162: douta=16'h3a4d;
3163: douta=16'h5351;
3164: douta=16'h6bd2;
3165: douta=16'h6c13;
3166: douta=16'h7434;
3167: douta=16'h8cf6;
3168: douta=16'h9d57;
3169: douta=16'ha577;
3170: douta=16'h324e;
3171: douta=16'h63b2;
3172: douta=16'hc618;
3173: douta=16'h7454;
3174: douta=16'h9d17;
3175: douta=16'h7413;
3176: douta=16'h84d7;
3177: douta=16'h6c14;
3178: douta=16'h9536;
3179: douta=16'hbdf9;
3180: douta=16'h63b1;
3181: douta=16'h2125;
3182: douta=16'h18e5;
3183: douta=16'h18e5;
3184: douta=16'h10e5;
3185: douta=16'h18e5;
3186: douta=16'h10e4;
3187: douta=16'h10a3;
3188: douta=16'h31a8;
3189: douta=16'h5acd;
3190: douta=16'h7414;
3191: douta=16'h7414;
3192: douta=16'h84f9;
3193: douta=16'h74d9;
3194: douta=16'h6457;
3195: douta=16'h74f9;
3196: douta=16'h853a;
3197: douta=16'h7d1a;
3198: douta=16'h6cb9;
3199: douta=16'h6cb9;
3200: douta=16'h74d9;
3201: douta=16'h4bf7;
3202: douta=16'h6478;
3203: douta=16'h6c78;
3204: douta=16'h6437;
3205: douta=16'h7cfa;
3206: douta=16'h74b9;
3207: douta=16'h5c16;
3208: douta=16'h7499;
3209: douta=16'h7d1a;
3210: douta=16'h7cf9;
3211: douta=16'h7cd9;
3212: douta=16'h6c57;
3213: douta=16'h6c78;
3214: douta=16'h6cb9;
3215: douta=16'h74da;
3216: douta=16'h855b;
3217: douta=16'h7d3b;
3218: douta=16'h6cb9;
3219: douta=16'h6cb9;
3220: douta=16'h855c;
3221: douta=16'h857b;
3222: douta=16'h74da;
3223: douta=16'h6cb8;
3224: douta=16'h751a;
3225: douta=16'h74da;
3226: douta=16'h857c;
3227: douta=16'h6436;
3228: douta=16'h5bf5;
3229: douta=16'h42d0;
3230: douta=16'h42af;
3231: douta=16'h2989;
3232: douta=16'h0062;
3233: douta=16'h08a4;
3234: douta=16'h10a4;
3235: douta=16'h08a4;
3236: douta=16'h10c4;
3237: douta=16'h0863;
3238: douta=16'h32af;
3239: douta=16'h5b92;
3240: douta=16'h7cb5;
3241: douta=16'h8454;
3242: douta=16'h6bb2;
3243: douta=16'h7413;
3244: douta=16'h328e;
3245: douta=16'h3acf;
3246: douta=16'h3acf;
3247: douta=16'h7c94;
3248: douta=16'h6bf2;
3249: douta=16'h94b5;
3250: douta=16'h53b4;
3251: douta=16'h21ec;
3252: douta=16'h4b32;
3253: douta=16'h6c35;
3254: douta=16'h3ad1;
3255: douta=16'h53b4;
3256: douta=16'h957a;
3257: douta=16'h4375;
3258: douta=16'h4bb5;
3259: douta=16'h3b33;
3260: douta=16'h5bf5;
3261: douta=16'h5416;
3262: douta=16'h5bb3;
3263: douta=16'h8519;
3264: douta=16'h4374;
3265: douta=16'h32b0;
3266: douta=16'h6416;
3267: douta=16'h6437;
3268: douta=16'h63d4;
3269: douta=16'h42cf;
3270: douta=16'h6436;
3271: douta=16'h4b52;
3272: douta=16'h6371;
3273: douta=16'h94f6;
3274: douta=16'h8cf7;
3275: douta=16'h8c74;
3276: douta=16'ha579;
3277: douta=16'h84d8;
3278: douta=16'ha536;
3279: douta=16'h5b50;
3280: douta=16'had56;
3281: douta=16'hd658;
3282: douta=16'hce79;
3283: douta=16'hbdf8;
3284: douta=16'h6c34;
3285: douta=16'h73d1;
3286: douta=16'had36;
3287: douta=16'h7433;
3288: douta=16'h9d15;
3289: douta=16'hce58;
3290: douta=16'hef3a;
3291: douta=16'ha535;
3292: douta=16'h9d36;
3293: douta=16'hd678;
3294: douta=16'hd678;
3295: douta=16'he698;
3296: douta=16'hd698;
3297: douta=16'hef3a;
3298: douta=16'ha4b3;
3299: douta=16'hce37;
3300: douta=16'h8411;
3301: douta=16'h9c91;
3302: douta=16'hef5a;
3303: douta=16'hb595;
3304: douta=16'h632d;
3305: douta=16'h83ae;
3306: douta=16'ha511;
3307: douta=16'h9470;
3308: douta=16'he6b8;
3309: douta=16'hde77;
3310: douta=16'h6b2c;
3311: douta=16'h4aad;
3312: douta=16'hd676;
3313: douta=16'he6d7;
3314: douta=16'hc5d4;
3315: douta=16'hacf2;
3316: douta=16'h532d;
3317: douta=16'h9450;
3318: douta=16'h7c51;
3319: douta=16'h9d55;
3320: douta=16'h8431;
3321: douta=16'hb5d7;
3322: douta=16'hb5d7;
3323: douta=16'h5b50;
3324: douta=16'h7c74;
3325: douta=16'h73f1;
3326: douta=16'had96;
3327: douta=16'hc638;
3328: douta=16'h9d36;
3329: douta=16'hc658;
3330: douta=16'h8476;
3331: douta=16'h4353;
3332: douta=16'h6bd3;
3333: douta=16'h7433;
3334: douta=16'h8cf6;
3335: douta=16'h6477;
3336: douta=16'hbe39;
3337: douta=16'h5bb2;
3338: douta=16'h5c15;
3339: douta=16'h4311;
3340: douta=16'h4332;
3341: douta=16'h4b73;
3342: douta=16'h6c98;
3343: douta=16'h7c96;
3344: douta=16'h855a;
3345: douta=16'h7cd8;
3346: douta=16'h6436;
3347: douta=16'h53d4;
3348: douta=16'h32b1;
3349: douta=16'ha5b9;
3350: douta=16'h3aaf;
3351: douta=16'h4b31;
3352: douta=16'ha535;
3353: douta=16'hbe59;
3354: douta=16'h8517;
3355: douta=16'h84d7;
3356: douta=16'hbe3a;
3357: douta=16'h6bf4;
3358: douta=16'h5371;
3359: douta=16'h4aad;
3360: douta=16'h3a4c;
3361: douta=16'h5392;
3362: douta=16'h7c96;
3363: douta=16'h9515;
3364: douta=16'h9d56;
3365: douta=16'h3a4e;
3366: douta=16'h5bd3;
3367: douta=16'hb659;
3368: douta=16'h6c35;
3369: douta=16'h84f8;
3370: douta=16'h8d37;
3371: douta=16'h1127;
3372: douta=16'h18e5;
3373: douta=16'h2125;
3374: douta=16'h1905;
3375: douta=16'h1905;
3376: douta=16'h1083;
3377: douta=16'h39c8;
3378: douta=16'h422a;
3379: douta=16'h8434;
3380: douta=16'h7c55;
3381: douta=16'h7cd9;
3382: douta=16'h853a;
3383: douta=16'h855a;
3384: douta=16'h7cd9;
3385: douta=16'h9dbc;
3386: douta=16'ha61c;
3387: douta=16'h959b;
3388: douta=16'h74fa;
3389: douta=16'h74d9;
3390: douta=16'h74fa;
3391: douta=16'h6c57;
3392: douta=16'h6c98;
3393: douta=16'h855b;
3394: douta=16'h6479;
3395: douta=16'h6478;
3396: douta=16'h6478;
3397: douta=16'h6457;
3398: douta=16'h6458;
3399: douta=16'h7d1a;
3400: douta=16'h7499;
3401: douta=16'h6c98;
3402: douta=16'h74da;
3403: douta=16'h7d3b;
3404: douta=16'h74d9;
3405: douta=16'h7d1a;
3406: douta=16'h74d9;
3407: douta=16'h74d9;
3408: douta=16'h6c98;
3409: douta=16'h74d9;
3410: douta=16'h8d9b;
3411: douta=16'h855b;
3412: douta=16'h751a;
3413: douta=16'h751a;
3414: douta=16'h7d1b;
3415: douta=16'h6cb9;
3416: douta=16'h6498;
3417: douta=16'h6cb8;
3418: douta=16'h6457;
3419: douta=16'h7d3b;
3420: douta=16'h751b;
3421: douta=16'h755b;
3422: douta=16'h74fa;
3423: douta=16'h6c77;
3424: douta=16'h42cf;
3425: douta=16'h29eb;
3426: douta=16'h2189;
3427: douta=16'h08a4;
3428: douta=16'h10c5;
3429: douta=16'h10e5;
3430: douta=16'h08c4;
3431: douta=16'h0064;
3432: douta=16'h0907;
3433: douta=16'h6414;
3434: douta=16'h7c53;
3435: douta=16'h7c13;
3436: douta=16'h9d16;
3437: douta=16'h8cb6;
3438: douta=16'h7c55;
3439: douta=16'h1989;
3440: douta=16'h6bd3;
3441: douta=16'h42cf;
3442: douta=16'h3b12;
3443: douta=16'h5b72;
3444: douta=16'h3b33;
3445: douta=16'h11cc;
3446: douta=16'h3ad0;
3447: douta=16'h4312;
3448: douta=16'h7498;
3449: douta=16'h6c56;
3450: douta=16'h955a;
3451: douta=16'h53d5;
3452: douta=16'h53d5;
3453: douta=16'h3af2;
3454: douta=16'h2a4e;
3455: douta=16'h53d4;
3456: douta=16'h5c37;
3457: douta=16'h42d1;
3458: douta=16'h6c77;
3459: douta=16'h3b33;
3460: douta=16'h6c36;
3461: douta=16'h7cb8;
3462: douta=16'h5b93;
3463: douta=16'h953a;
3464: douta=16'h5310;
3465: douta=16'h6bd3;
3466: douta=16'h5b51;
3467: douta=16'h8454;
3468: douta=16'h94f6;
3469: douta=16'ha5ba;
3470: douta=16'h8cb5;
3471: douta=16'h6391;
3472: douta=16'h6b90;
3473: douta=16'h8432;
3474: douta=16'had55;
3475: douta=16'he6da;
3476: douta=16'hadd9;
3477: douta=16'hc5f9;
3478: douta=16'h8494;
3479: douta=16'ha557;
3480: douta=16'h6392;
3481: douta=16'h94f5;
3482: douta=16'h94d3;
3483: douta=16'hd679;
3484: douta=16'hb5d8;
3485: douta=16'hd698;
3486: douta=16'h9d56;
3487: douta=16'h8472;
3488: douta=16'hb595;
3489: douta=16'hd698;
3490: douta=16'he6f9;
3491: douta=16'hde99;
3492: douta=16'h73f1;
3493: douta=16'h326c;
3494: douta=16'hbd94;
3495: douta=16'hbdb4;
3496: douta=16'hcdd4;
3497: douta=16'hde77;
3498: douta=16'h5b0d;
3499: douta=16'h52cd;
3500: douta=16'hc5d4;
3501: douta=16'hd657;
3502: douta=16'hd616;
3503: douta=16'h632c;
3504: douta=16'hd697;
3505: douta=16'h8c4f;
3506: douta=16'ha512;
3507: douta=16'ha4f1;
3508: douta=16'h8431;
3509: douta=16'hc5d4;
3510: douta=16'h7c30;
3511: douta=16'h530f;
3512: douta=16'h7b8e;
3513: douta=16'h9d34;
3514: douta=16'he71a;
3515: douta=16'h73f2;
3516: douta=16'h9d16;
3517: douta=16'h5b51;
3518: douta=16'h9d76;
3519: douta=16'h42ee;
3520: douta=16'h7433;
3521: douta=16'h4b30;
3522: douta=16'h8cd6;
3523: douta=16'h5bf5;
3524: douta=16'h94f6;
3525: douta=16'ha598;
3526: douta=16'h3aaf;
3527: douta=16'h5373;
3528: douta=16'h9517;
3529: douta=16'h9579;
3530: douta=16'h6478;
3531: douta=16'h8496;
3532: douta=16'h7c76;
3533: douta=16'h3312;
3534: douta=16'h4b94;
3535: douta=16'h63d5;
3536: douta=16'h3af1;
3537: douta=16'h95bb;
3538: douta=16'h7497;
3539: douta=16'h7498;
3540: douta=16'h4b94;
3541: douta=16'h6c55;
3542: douta=16'h5b2f;
3543: douta=16'h220d;
3544: douta=16'h5351;
3545: douta=16'h5372;
3546: douta=16'h63b3;
3547: douta=16'h6c14;
3548: douta=16'h7c96;
3549: douta=16'h5351;
3550: douta=16'h7455;
3551: douta=16'h9d36;
3552: douta=16'h6bd3;
3553: douta=16'h428f;
3554: douta=16'h428e;
3555: douta=16'h424b;
3556: douta=16'h7cb5;
3557: douta=16'h84b6;
3558: douta=16'h84d7;
3559: douta=16'h5bb3;
3560: douta=16'h21ec;
3561: douta=16'h7c54;
3562: douta=16'h322b;
3563: douta=16'h18c4;
3564: douta=16'h2126;
3565: douta=16'h2125;
3566: douta=16'h10e5;
3567: douta=16'h1083;
3568: douta=16'h522a;
3569: douta=16'h5b0e;
3570: douta=16'h7c74;
3571: douta=16'h7c98;
3572: douta=16'h851a;
3573: douta=16'h853a;
3574: douta=16'h8519;
3575: douta=16'h8d5b;
3576: douta=16'h8519;
3577: douta=16'h853b;
3578: douta=16'h959b;
3579: douta=16'ha5fc;
3580: douta=16'h853a;
3581: douta=16'h8d5b;
3582: douta=16'h74d9;
3583: douta=16'h6478;
3584: douta=16'h5c16;
3585: douta=16'h7cfa;
3586: douta=16'h74da;
3587: douta=16'h6cba;
3588: douta=16'h74da;
3589: douta=16'h74f9;
3590: douta=16'h7cf9;
3591: douta=16'h6cb9;
3592: douta=16'h74d9;
3593: douta=16'h6c99;
3594: douta=16'h6cb9;
3595: douta=16'h855b;
3596: douta=16'h7d5a;
3597: douta=16'h6cb9;
3598: douta=16'h857b;
3599: douta=16'h95bc;
3600: douta=16'h6437;
3601: douta=16'h74f9;
3602: douta=16'h7d3a;
3603: douta=16'h859b;
3604: douta=16'h74fa;
3605: douta=16'h74fa;
3606: douta=16'h7d1a;
3607: douta=16'h855b;
3608: douta=16'h74d9;
3609: douta=16'h6cb9;
3610: douta=16'h7d1a;
3611: douta=16'h5c37;
3612: douta=16'h7d5b;
3613: douta=16'h7d3b;
3614: douta=16'h7d5c;
3615: douta=16'h753b;
3616: douta=16'h6c37;
3617: douta=16'h4310;
3618: douta=16'h3a8e;
3619: douta=16'h10e4;
3620: douta=16'h0063;
3621: douta=16'h10e5;
3622: douta=16'h08c5;
3623: douta=16'h10c5;
3624: douta=16'h0884;
3625: douta=16'h42ef;
3626: douta=16'h7434;
3627: douta=16'h8473;
3628: douta=16'h9d35;
3629: douta=16'had77;
3630: douta=16'h7c53;
3631: douta=16'h7412;
3632: douta=16'h2a4e;
3633: douta=16'h2a4e;
3634: douta=16'h4b11;
3635: douta=16'h8cb6;
3636: douta=16'h5bb4;
3637: douta=16'h32b0;
3638: douta=16'h4332;
3639: douta=16'h2a6f;
3640: douta=16'h1a2f;
3641: douta=16'h851a;
3642: douta=16'h7497;
3643: douta=16'h6c57;
3644: douta=16'h6436;
3645: douta=16'h7498;
3646: douta=16'h19cd;
3647: douta=16'h4b73;
3648: douta=16'h3b34;
3649: douta=16'h3af1;
3650: douta=16'h6457;
3651: douta=16'h4b94;
3652: douta=16'h6c36;
3653: douta=16'h74b8;
3654: douta=16'h6c15;
3655: douta=16'h953a;
3656: douta=16'h6bd3;
3657: douta=16'h5330;
3658: douta=16'h7c34;
3659: douta=16'h8475;
3660: douta=16'hce39;
3661: douta=16'hadd9;
3662: douta=16'h7433;
3663: douta=16'h73d1;
3664: douta=16'h73f2;
3665: douta=16'h9cf5;
3666: douta=16'heefa;
3667: douta=16'hbd76;
3668: douta=16'hd69a;
3669: douta=16'h9cd5;
3670: douta=16'h6bf3;
3671: douta=16'h8cb4;
3672: douta=16'h94d5;
3673: douta=16'hd679;
3674: douta=16'hdeb8;
3675: douta=16'h4aae;
3676: douta=16'h9d15;
3677: douta=16'h8c52;
3678: douta=16'h94d4;
3679: douta=16'hb554;
3680: douta=16'hce36;
3681: douta=16'hfffc;
3682: douta=16'hbdb5;
3683: douta=16'hde78;
3684: douta=16'ha514;
3685: douta=16'h9450;
3686: douta=16'hde97;
3687: douta=16'hb552;
3688: douta=16'h9410;
3689: douta=16'hcdf5;
3690: douta=16'h5b6f;
3691: douta=16'h63af;
3692: douta=16'hef18;
3693: douta=16'he6d8;
3694: douta=16'hc5d4;
3695: douta=16'h8c0e;
3696: douta=16'hbdd4;
3697: douta=16'had31;
3698: douta=16'hbe15;
3699: douta=16'hbd93;
3700: douta=16'h634d;
3701: douta=16'hc615;
3702: douta=16'h328c;
3703: douta=16'h4a8d;
3704: douta=16'hacd3;
3705: douta=16'h94b4;
3706: douta=16'hbe59;
3707: douta=16'h52ef;
3708: douta=16'h7c11;
3709: douta=16'h6b90;
3710: douta=16'h5b4e;
3711: douta=16'h4a8c;
3712: douta=16'h9d14;
3713: douta=16'h9515;
3714: douta=16'h4b2f;
3715: douta=16'h7496;
3716: douta=16'h63b1;
3717: douta=16'h8cb5;
3718: douta=16'h328e;
3719: douta=16'h4b73;
3720: douta=16'h74d8;
3721: douta=16'h84f7;
3722: douta=16'h53d4;
3723: douta=16'h6c15;
3724: douta=16'h6c56;
3725: douta=16'h3b11;
3726: douta=16'h4b52;
3727: douta=16'h5c16;
3728: douta=16'h3af1;
3729: douta=16'h8d39;
3730: douta=16'h8d38;
3731: douta=16'h32b1;
3732: douta=16'h326f;
3733: douta=16'h52f0;
3734: douta=16'h4b52;
3735: douta=16'h7497;
3736: douta=16'h84d6;
3737: douta=16'h7496;
3738: douta=16'h7476;
3739: douta=16'had96;
3740: douta=16'h7c96;
3741: douta=16'h8495;
3742: douta=16'h52ef;
3743: douta=16'h73d1;
3744: douta=16'h63b2;
3745: douta=16'h94f5;
3746: douta=16'h9d36;
3747: douta=16'h8cf5;
3748: douta=16'h7c96;
3749: douta=16'h8cb7;
3750: douta=16'h5b93;
3751: douta=16'h31ea;
3752: douta=16'h1926;
3753: douta=16'h2146;
3754: douta=16'h2146;
3755: douta=16'h10c4;
3756: douta=16'h1063;
3757: douta=16'h7b8f;
3758: douta=16'h6b70;
3759: douta=16'h84b7;
3760: douta=16'h853a;
3761: douta=16'h74b9;
3762: douta=16'h8d1a;
3763: douta=16'h853a;
3764: douta=16'h8519;
3765: douta=16'h8d3a;
3766: douta=16'h8519;
3767: douta=16'h8519;
3768: douta=16'h853b;
3769: douta=16'h8d5b;
3770: douta=16'h851a;
3771: douta=16'h851a;
3772: douta=16'h7c77;
3773: douta=16'h7c97;
3774: douta=16'h851a;
3775: douta=16'h74b9;
3776: douta=16'h7d1a;
3777: douta=16'h8d7b;
3778: douta=16'h74ba;
3779: douta=16'h74fa;
3780: douta=16'h6cb9;
3781: douta=16'h7d3a;
3782: douta=16'h6478;
3783: douta=16'h751a;
3784: douta=16'h74da;
3785: douta=16'h74fa;
3786: douta=16'h7d1b;
3787: douta=16'h7d3a;
3788: douta=16'h7d3a;
3789: douta=16'h7d3a;
3790: douta=16'h751a;
3791: douta=16'h8d9c;
3792: douta=16'h7d1a;
3793: douta=16'h74b9;
3794: douta=16'h7d1a;
3795: douta=16'h74b9;
3796: douta=16'h6cb8;
3797: douta=16'h6478;
3798: douta=16'h7d1b;
3799: douta=16'h85bc;
3800: douta=16'h7d1a;
3801: douta=16'h6cb9;
3802: douta=16'h8dbc;
3803: douta=16'h6cd9;
3804: douta=16'h6cd9;
3805: douta=16'h6cd9;
3806: douta=16'h6cda;
3807: douta=16'h753b;
3808: douta=16'h6cba;
3809: douta=16'h7d7c;
3810: douta=16'h74fa;
3811: douta=16'h74d9;
3812: douta=16'h6c16;
3813: douta=16'h42cf;
3814: douta=16'h2168;
3815: douta=16'h0884;
3816: douta=16'h10c5;
3817: douta=16'h10e6;
3818: douta=16'h10c4;
3819: douta=16'h1169;
3820: douta=16'ha557;
3821: douta=16'h6bd3;
3822: douta=16'h6bb1;
3823: douta=16'h4b0f;
3824: douta=16'hb5d8;
3825: douta=16'h63b2;
3826: douta=16'h222f;
3827: douta=16'h3af1;
3828: douta=16'h2a6e;
3829: douta=16'h5392;
3830: douta=16'h7498;
3831: douta=16'h7cd9;
3832: douta=16'h9559;
3833: douta=16'h8cf8;
3834: douta=16'h6478;
3835: douta=16'h4332;
3836: douta=16'h4b95;
3837: douta=16'h32b0;
3838: douta=16'h6478;
3839: douta=16'ha5bc;
3840: douta=16'h224f;
3841: douta=16'h32b0;
3842: douta=16'h6415;
3843: douta=16'h6415;
3844: douta=16'h5bf5;
3845: douta=16'h6c57;
3846: douta=16'h4b11;
3847: douta=16'h4b73;
3848: douta=16'h6bd4;
3849: douta=16'h9cb6;
3850: douta=16'h8cb5;
3851: douta=16'h6bf4;
3852: douta=16'hce39;
3853: douta=16'h8474;
3854: douta=16'h5b92;
3855: douta=16'ha536;
3856: douta=16'hd659;
3857: douta=16'had97;
3858: douta=16'hbd97;
3859: douta=16'had76;
3860: douta=16'hb5b7;
3861: douta=16'h8cb5;
3862: douta=16'h94d5;
3863: douta=16'hffdb;
3864: douta=16'hb5b7;
3865: douta=16'h8473;
3866: douta=16'ha534;
3867: douta=16'h8c73;
3868: douta=16'hb5d6;
3869: douta=16'hff7b;
3870: douta=16'hffbc;
3871: douta=16'hc5b4;
3872: douta=16'h4acd;
3873: douta=16'h83ef;
3874: douta=16'h9c92;
3875: douta=16'hde98;
3876: douta=16'hce16;
3877: douta=16'h8bce;
3878: douta=16'hce57;
3879: douta=16'h634e;
3880: douta=16'h428a;
3881: douta=16'hbd74;
3882: douta=16'h946f;
3883: douta=16'ha4b1;
3884: douta=16'ha4d0;
3885: douta=16'hbd72;
3886: douta=16'h6b8c;
3887: douta=16'h5b0c;
3888: douta=16'hb593;
3889: douta=16'hfffb;
3890: douta=16'h840f;
3891: douta=16'hd615;
3892: douta=16'h630c;
3893: douta=16'h94b2;
3894: douta=16'h634d;
3895: douta=16'h5b0e;
3896: douta=16'hde77;
3897: douta=16'h5b50;
3898: douta=16'h5b90;
3899: douta=16'h5aaa;
3900: douta=16'ha4f3;
3901: douta=16'hbd94;
3902: douta=16'h3a2a;
3903: douta=16'h7c11;
3904: douta=16'h63b0;
3905: douta=16'h324d;
3906: douta=16'h4b71;
3907: douta=16'h0044;
3908: douta=16'h5bb3;
3909: douta=16'h3b11;
3910: douta=16'h5393;
3911: douta=16'h5372;
3912: douta=16'h6414;
3913: douta=16'h42f0;
3914: douta=16'h4311;
3915: douta=16'h5351;
3916: douta=16'h7519;
3917: douta=16'h4bd6;
3918: douta=16'h957a;
3919: douta=16'h859d;
3920: douta=16'h5395;
3921: douta=16'h4aaf;
3922: douta=16'h3ad1;
3923: douta=16'h53d5;
3924: douta=16'h53b4;
3925: douta=16'h7cb6;
3926: douta=16'h53f5;
3927: douta=16'h5b73;
3928: douta=16'h6456;
3929: douta=16'h42b0;
3930: douta=16'h2a4e;
3931: douta=16'h5b91;
3932: douta=16'h4b11;
3933: douta=16'h6bf2;
3934: douta=16'ha598;
3935: douta=16'ha578;
3936: douta=16'h9d77;
3937: douta=16'h6392;
3938: douta=16'h324e;
3939: douta=16'h5b50;
3940: douta=16'h5b71;
3941: douta=16'h5b71;
3942: douta=16'h3a4b;
3943: douta=16'h2966;
3944: douta=16'h2966;
3945: douta=16'h2146;
3946: douta=16'h49e8;
3947: douta=16'h7b6e;
3948: douta=16'h8cb5;
3949: douta=16'h7498;
3950: douta=16'h8519;
3951: douta=16'h953a;
3952: douta=16'h7d19;
3953: douta=16'h851a;
3954: douta=16'h8d5b;
3955: douta=16'h851a;
3956: douta=16'h851a;
3957: douta=16'h8d7b;
3958: douta=16'h8d5b;
3959: douta=16'h851a;
3960: douta=16'h853a;
3961: douta=16'h8519;
3962: douta=16'h8d5b;
3963: douta=16'h853a;
3964: douta=16'h855a;
3965: douta=16'h8d7b;
3966: douta=16'h8519;
3967: douta=16'h959b;
3968: douta=16'h8d7b;
3969: douta=16'h853a;
3970: douta=16'h853a;
3971: douta=16'h6cb9;
3972: douta=16'h6458;
3973: douta=16'h6438;
3974: douta=16'h6c99;
3975: douta=16'h6478;
3976: douta=16'h6c99;
3977: douta=16'h7d3b;
3978: douta=16'h6478;
3979: douta=16'h7d1b;
3980: douta=16'h7d3a;
3981: douta=16'h8dbc;
3982: douta=16'h95dd;
3983: douta=16'h7d3a;
3984: douta=16'h7d1a;
3985: douta=16'h855b;
3986: douta=16'h855a;
3987: douta=16'h7d1a;
3988: douta=16'h6cd9;
3989: douta=16'h6c99;
3990: douta=16'h8d9b;
3991: douta=16'h6478;
3992: douta=16'h7d1a;
3993: douta=16'h74da;
3994: douta=16'h7d3a;
3995: douta=16'h7d1a;
3996: douta=16'h7d1a;
3997: douta=16'h6478;
3998: douta=16'h751a;
3999: douta=16'h753b;
4000: douta=16'h6478;
4001: douta=16'h74d9;
4002: douta=16'h74f9;
4003: douta=16'h74fb;
4004: douta=16'h751a;
4005: douta=16'h6cda;
4006: douta=16'h5353;
4007: douta=16'h29aa;
4008: douta=16'h2168;
4009: douta=16'h08c5;
4010: douta=16'h1107;
4011: douta=16'h1127;
4012: douta=16'h00c6;
4013: douta=16'h42ee;
4014: douta=16'ha516;
4015: douta=16'h73f4;
4016: douta=16'h19ab;
4017: douta=16'h42d0;
4018: douta=16'hb63b;
4019: douta=16'h9d79;
4020: douta=16'h73f4;
4021: douta=16'h6416;
4022: douta=16'h5c38;
4023: douta=16'h4374;
4024: douta=16'h2ad2;
4025: douta=16'h6c97;
4026: douta=16'h7c76;
4027: douta=16'h6cb9;
4028: douta=16'h6c57;
4029: douta=16'h32f2;
4030: douta=16'h2a8f;
4031: douta=16'h3b12;
4032: douta=16'h3b33;
4033: douta=16'h2a90;
4034: douta=16'h6436;
4035: douta=16'h5bd4;
4036: douta=16'h5b94;
4037: douta=16'h7d19;
4038: douta=16'h5b92;
4039: douta=16'h8d19;
4040: douta=16'h5b93;
4041: douta=16'h5330;
4042: douta=16'h6c14;
4043: douta=16'h6bd3;
4044: douta=16'hbdd7;
4045: douta=16'ha577;
4046: douta=16'h84b6;
4047: douta=16'h6bb1;
4048: douta=16'h7c32;
4049: douta=16'h7412;
4050: douta=16'he6b9;
4051: douta=16'hb596;
4052: douta=16'hce59;
4053: douta=16'h6bd2;
4054: douta=16'h6bf3;
4055: douta=16'hb596;
4056: douta=16'hb556;
4057: douta=16'hb576;
4058: douta=16'hb5b6;
4059: douta=16'h52ef;
4060: douta=16'hb5f8;
4061: douta=16'hc5d6;
4062: douta=16'hffbb;
4063: douta=16'hef19;
4064: douta=16'hb575;
4065: douta=16'ha4b3;
4066: douta=16'h62ee;
4067: douta=16'hcdd6;
4068: douta=16'ha4f3;
4069: douta=16'he696;
4070: douta=16'hd676;
4071: douta=16'h7bed;
4072: douta=16'h528b;
4073: douta=16'h8c0f;
4074: douta=16'h840f;
4075: douta=16'had31;
4076: douta=16'heef8;
4077: douta=16'he6f8;
4078: douta=16'hc615;
4079: douta=16'h41c8;
4080: douta=16'hb593;
4081: douta=16'he6d7;
4082: douta=16'had10;
4083: douta=16'hef18;
4084: douta=16'h734c;
4085: douta=16'h8cd3;
4086: douta=16'h2a0a;
4087: douta=16'h4aad;
4088: douta=16'hbd95;
4089: douta=16'h73d1;
4090: douta=16'h6bf1;
4091: douta=16'h7bcf;
4092: douta=16'h8410;
4093: douta=16'h7bcf;
4094: douta=16'h4a8b;
4095: douta=16'h29a7;
4096: douta=16'h3a8d;
4097: douta=16'h31ea;
4098: douta=16'h3acf;
4099: douta=16'h29aa;
4100: douta=16'h00c6;
4101: douta=16'h1968;
4102: douta=16'h2a2d;
4103: douta=16'h5373;
4104: douta=16'h6415;
4105: douta=16'h5352;
4106: douta=16'h222d;
4107: douta=16'h5b71;
4108: douta=16'h5c15;
4109: douta=16'h4b73;
4110: douta=16'h63f4;
4111: douta=16'h4bf6;
4112: douta=16'h3b13;
4113: douta=16'h8d59;
4114: douta=16'h4b74;
4115: douta=16'h3af2;
4116: douta=16'h32d1;
4117: douta=16'h5bb4;
4118: douta=16'h2a4e;
4119: douta=16'h8d7a;
4120: douta=16'h7cd8;
4121: douta=16'h63d3;
4122: douta=16'h5372;
4123: douta=16'h7c55;
4124: douta=16'h7413;
4125: douta=16'h6b91;
4126: douta=16'h7453;
4127: douta=16'h5b91;
4128: douta=16'h9d77;
4129: douta=16'h8cf5;
4130: douta=16'h4312;
4131: douta=16'h4310;
4132: douta=16'h4b10;
4133: douta=16'h5350;
4134: douta=16'h2105;
4135: douta=16'h2967;
4136: douta=16'h2145;
4137: douta=16'h10a4;
4138: douta=16'h83af;
4139: douta=16'h73d1;
4140: douta=16'h7c96;
4141: douta=16'h7498;
4142: douta=16'h7457;
4143: douta=16'h8d3a;
4144: douta=16'h851a;
4145: douta=16'h8519;
4146: douta=16'h7cf9;
4147: douta=16'h959c;
4148: douta=16'h7cf9;
4149: douta=16'h853a;
4150: douta=16'h8d7b;
4151: douta=16'h959b;
4152: douta=16'h8d5b;
4153: douta=16'h7cf9;
4154: douta=16'h8d5a;
4155: douta=16'h851a;
4156: douta=16'h95bc;
4157: douta=16'h8d7b;
4158: douta=16'h851a;
4159: douta=16'h8d7b;
4160: douta=16'h8d5a;
4161: douta=16'h95bc;
4162: douta=16'h7cf9;
4163: douta=16'h7d3b;
4164: douta=16'h7cd9;
4165: douta=16'h6498;
4166: douta=16'h859c;
4167: douta=16'h6cba;
4168: douta=16'h4b75;
4169: douta=16'h7d7c;
4170: douta=16'h9e5f;
4171: douta=16'h6499;
4172: douta=16'h74d9;
4173: douta=16'h74fa;
4174: douta=16'h95bc;
4175: douta=16'h961d;
4176: douta=16'h7d3b;
4177: douta=16'h857b;
4178: douta=16'h857b;
4179: douta=16'h8d9b;
4180: douta=16'h8d9b;
4181: douta=16'h855b;
4182: douta=16'h74f9;
4183: douta=16'h74d9;
4184: douta=16'h7cfa;
4185: douta=16'h7d1a;
4186: douta=16'h6c98;
4187: douta=16'h6498;
4188: douta=16'h7d1a;
4189: douta=16'h74d9;
4190: douta=16'h74d9;
4191: douta=16'h6498;
4192: douta=16'h6c98;
4193: douta=16'h6c98;
4194: douta=16'h6cb9;
4195: douta=16'h753b;
4196: douta=16'h751a;
4197: douta=16'h6cfa;
4198: douta=16'h74fa;
4199: douta=16'h5332;
4200: douta=16'h324d;
4201: douta=16'h2168;
4202: douta=16'h08c5;
4203: douta=16'h1106;
4204: douta=16'h10e7;
4205: douta=16'h08e6;
4206: douta=16'h4310;
4207: douta=16'h94b6;
4208: douta=16'h5351;
4209: douta=16'h5372;
4210: douta=16'h42f1;
4211: douta=16'h4b11;
4212: douta=16'h9d16;
4213: douta=16'h955a;
4214: douta=16'h6c98;
4215: douta=16'h74b8;
4216: douta=16'h53d5;
4217: douta=16'h2291;
4218: douta=16'h7cb7;
4219: douta=16'h84d8;
4220: douta=16'ha59a;
4221: douta=16'h5c16;
4222: douta=16'h6477;
4223: douta=16'h53d4;
4224: douta=16'h2a6f;
4225: douta=16'h19ad;
4226: douta=16'h42d1;
4227: douta=16'h32b0;
4228: douta=16'h5c15;
4229: douta=16'h63d4;
4230: douta=16'h63f4;
4231: douta=16'h7c96;
4232: douta=16'h5bb3;
4233: douta=16'h6b91;
4234: douta=16'h9517;
4235: douta=16'h7c74;
4236: douta=16'hce38;
4237: douta=16'h8474;
4238: douta=16'h2a70;
4239: douta=16'h8454;
4240: douta=16'had75;
4241: douta=16'had56;
4242: douta=16'hce38;
4243: douta=16'hb597;
4244: douta=16'h8c93;
4245: douta=16'h63d3;
4246: douta=16'hbdb6;
4247: douta=16'had95;
4248: douta=16'h94b4;
4249: douta=16'h6bb2;
4250: douta=16'h94b2;
4251: douta=16'h8411;
4252: douta=16'hded8;
4253: douta=16'hd637;
4254: douta=16'hffdb;
4255: douta=16'h9cd3;
4256: douta=16'hce36;
4257: douta=16'hb575;
4258: douta=16'h7bd0;
4259: douta=16'hce16;
4260: douta=16'hb533;
4261: douta=16'h9430;
4262: douta=16'had53;
4263: douta=16'h632d;
4264: douta=16'h3a2a;
4265: douta=16'h8c2e;
4266: douta=16'h944e;
4267: douta=16'h734b;
4268: douta=16'hffba;
4269: douta=16'hd698;
4270: douta=16'hb5f4;
4271: douta=16'h62ec;
4272: douta=16'h5b4c;
4273: douta=16'h7c2f;
4274: douta=16'h4a8a;
4275: douta=16'h740f;
4276: douta=16'h4a28;
4277: douta=16'h6bf0;
4278: douta=16'h426b;
4279: douta=16'h7bcf;
4280: douta=16'hce76;
4281: douta=16'h8c30;
4282: douta=16'h634e;
4283: douta=16'h840f;
4284: douta=16'h73cf;
4285: douta=16'h8c4f;
4286: douta=16'h2945;
4287: douta=16'h63d1;
4288: douta=16'h4aef;
4289: douta=16'h63d2;
4290: douta=16'h0881;
4291: douta=16'h0840;
4292: douta=16'h2147;
4293: douta=16'h320b;
4294: douta=16'h3a8f;
4295: douta=16'h2a4d;
4296: douta=16'h3ab0;
4297: douta=16'h328f;
4298: douta=16'h5371;
4299: douta=16'h2a4e;
4300: douta=16'h32b0;
4301: douta=16'h63f4;
4302: douta=16'h8d38;
4303: douta=16'h3b34;
4304: douta=16'h5bd4;
4305: douta=16'h7497;
4306: douta=16'h3b11;
4307: douta=16'h5352;
4308: douta=16'h84d6;
4309: douta=16'h7c96;
4310: douta=16'h6436;
4311: douta=16'h9d16;
4312: douta=16'h5b93;
4313: douta=16'h5bd4;
4314: douta=16'h4b31;
4315: douta=16'h324e;
4316: douta=16'h42ef;
4317: douta=16'h21ec;
4318: douta=16'h8cd5;
4319: douta=16'h6bf4;
4320: douta=16'h8d59;
4321: douta=16'h8433;
4322: douta=16'h7433;
4323: douta=16'h6c13;
4324: douta=16'h2945;
4325: douta=16'h31a7;
4326: douta=16'h10e5;
4327: douta=16'h8b8d;
4328: douta=16'h9452;
4329: douta=16'h7c76;
4330: douta=16'h84d8;
4331: douta=16'h7c98;
4332: douta=16'h7497;
4333: douta=16'h7c98;
4334: douta=16'h7477;
4335: douta=16'h8d5a;
4336: douta=16'h63f5;
4337: douta=16'h63f6;
4338: douta=16'h7cd9;
4339: douta=16'h9dbc;
4340: douta=16'h959c;
4341: douta=16'h853a;
4342: douta=16'h8d5a;
4343: douta=16'h8d5a;
4344: douta=16'h8519;
4345: douta=16'h7cf9;
4346: douta=16'h8d7b;
4347: douta=16'h853a;
4348: douta=16'h8d5b;
4349: douta=16'h8d9b;
4350: douta=16'h851a;
4351: douta=16'h95bc;
4352: douta=16'h95bc;
4353: douta=16'h957b;
4354: douta=16'h8d5b;
4355: douta=16'h8d5b;
4356: douta=16'h8d5b;
4357: douta=16'h8d7b;
4358: douta=16'h8d9b;
4359: douta=16'h6cba;
4360: douta=16'h6478;
4361: douta=16'h8dbd;
4362: douta=16'h859c;
4363: douta=16'h6cba;
4364: douta=16'h74fa;
4365: douta=16'h7d5b;
4366: douta=16'h7d1a;
4367: douta=16'h74f9;
4368: douta=16'h6cb9;
4369: douta=16'h8d9c;
4370: douta=16'h6cb9;
4371: douta=16'h6c99;
4372: douta=16'h7d5b;
4373: douta=16'h74d9;
4374: douta=16'h855b;
4375: douta=16'h8d9b;
4376: douta=16'h74d9;
4377: douta=16'h855b;
4378: douta=16'h7d3a;
4379: douta=16'h7d1a;
4380: douta=16'h74fa;
4381: douta=16'h857b;
4382: douta=16'h857b;
4383: douta=16'h6cb9;
4384: douta=16'h753a;
4385: douta=16'h857b;
4386: douta=16'h7d3b;
4387: douta=16'h6c78;
4388: douta=16'h6cd9;
4389: douta=16'h6cb9;
4390: douta=16'h6cb9;
4391: douta=16'h74fa;
4392: douta=16'h753b;
4393: douta=16'h6cba;
4394: douta=16'h3a4c;
4395: douta=16'h2168;
4396: douta=16'h1106;
4397: douta=16'h1127;
4398: douta=16'h1127;
4399: douta=16'h7456;
4400: douta=16'h4332;
4401: douta=16'h5393;
4402: douta=16'h9d16;
4403: douta=16'hb5da;
4404: douta=16'h9539;
4405: douta=16'h4b53;
4406: douta=16'h2a90;
4407: douta=16'h222f;
4408: douta=16'h2ab0;
4409: douta=16'h7497;
4410: douta=16'h959b;
4411: douta=16'h4b75;
4412: douta=16'h5bd4;
4413: douta=16'h3b12;
4414: douta=16'h53d4;
4415: douta=16'h4b94;
4416: douta=16'h32f2;
4417: douta=16'h53d5;
4418: douta=16'h7457;
4419: douta=16'h6477;
4420: douta=16'h4373;
4421: douta=16'h5373;
4422: douta=16'h198b;
4423: douta=16'h6c14;
4424: douta=16'h7455;
4425: douta=16'h94d6;
4426: douta=16'h8454;
4427: douta=16'h73f3;
4428: douta=16'h8473;
4429: douta=16'h7c12;
4430: douta=16'h9d56;
4431: douta=16'hbdd8;
4432: douta=16'h8c94;
4433: douta=16'ha557;
4434: douta=16'h9cb5;
4435: douta=16'h9d15;
4436: douta=16'hc5f7;
4437: douta=16'ha556;
4438: douta=16'h9cd4;
4439: douta=16'hb575;
4440: douta=16'h8cb3;
4441: douta=16'had55;
4442: douta=16'hbdb5;
4443: douta=16'hde98;
4444: douta=16'h8474;
4445: douta=16'hde98;
4446: douta=16'h8c72;
4447: douta=16'ha514;
4448: douta=16'h73f0;
4449: douta=16'hce15;
4450: douta=16'hcdf5;
4451: douta=16'hef19;
4452: douta=16'hacd1;
4453: douta=16'h5acb;
4454: douta=16'hd655;
4455: douta=16'hacf1;
4456: douta=16'hac8f;
4457: douta=16'hff38;
4458: douta=16'h5289;
4459: douta=16'h8410;
4460: douta=16'hb510;
4461: douta=16'had92;
4462: douta=16'h7bcd;
4463: douta=16'h62cb;
4464: douta=16'h10e4;
4465: douta=16'h1926;
4466: douta=16'h18e5;
4467: douta=16'h1905;
4468: douta=16'h736d;
4469: douta=16'h73ae;
4470: douta=16'h9c91;
4471: douta=16'hc5b5;
4472: douta=16'had32;
4473: douta=16'h31ea;
4474: douta=16'h4a8c;
4475: douta=16'h9cb0;
4476: douta=16'h8470;
4477: douta=16'ha574;
4478: douta=16'h5b4e;
4479: douta=16'h3a6e;
4480: douta=16'h4aae;
4481: douta=16'h4a4b;
4482: douta=16'h0840;
4483: douta=16'h1083;
4484: douta=16'h1082;
4485: douta=16'h0860;
4486: douta=16'h2967;
4487: douta=16'h3aaf;
4488: douta=16'h0108;
4489: douta=16'h2a2c;
4490: douta=16'h5393;
4491: douta=16'h322d;
4492: douta=16'h3b73;
4493: douta=16'h6c56;
4494: douta=16'h5393;
4495: douta=16'h42f1;
4496: douta=16'h4b53;
4497: douta=16'h6436;
4498: douta=16'h5c37;
4499: douta=16'h6bf2;
4500: douta=16'h9dba;
4501: douta=16'h6c35;
4502: douta=16'h5352;
4503: douta=16'h6bf5;
4504: douta=16'h4b94;
4505: douta=16'h32b1;
4506: douta=16'h7c56;
4507: douta=16'h6c15;
4508: douta=16'h63d3;
4509: douta=16'h6414;
4510: douta=16'h63d3;
4511: douta=16'ha599;
4512: douta=16'h42ef;
4513: douta=16'h42ae;
4514: douta=16'h4aad;
4515: douta=16'h3147;
4516: douta=16'h2988;
4517: douta=16'h41a6;
4518: douta=16'h9bee;
4519: douta=16'h7477;
4520: douta=16'h84f8;
4521: douta=16'h7cb7;
4522: douta=16'h84f8;
4523: douta=16'h7c97;
4524: douta=16'h7c97;
4525: douta=16'h7cb8;
4526: douta=16'h84f9;
4527: douta=16'h84d8;
4528: douta=16'h6c36;
4529: douta=16'h84f9;
4530: douta=16'h7cd8;
4531: douta=16'h4b12;
4532: douta=16'h8d7b;
4533: douta=16'h957b;
4534: douta=16'h9dbc;
4535: douta=16'h8d5a;
4536: douta=16'h851a;
4537: douta=16'h6c36;
4538: douta=16'h84d9;
4539: douta=16'h84d9;
4540: douta=16'h8d3a;
4541: douta=16'h8d5b;
4542: douta=16'h851a;
4543: douta=16'h851a;
4544: douta=16'h74b8;
4545: douta=16'h8d5a;
4546: douta=16'h959b;
4547: douta=16'h957b;
4548: douta=16'h957b;
4549: douta=16'h959c;
4550: douta=16'h95bc;
4551: douta=16'h95bc;
4552: douta=16'h6c98;
4553: douta=16'h74da;
4554: douta=16'h6c99;
4555: douta=16'h6cb9;
4556: douta=16'h859c;
4557: douta=16'h4b75;
4558: douta=16'h857c;
4559: douta=16'h8dbc;
4560: douta=16'h7d3b;
4561: douta=16'h74d9;
4562: douta=16'h855b;
4563: douta=16'h9e3e;
4564: douta=16'h6cb9;
4565: douta=16'h859c;
4566: douta=16'h855b;
4567: douta=16'h7d5b;
4568: douta=16'h7d3b;
4569: douta=16'h7d5b;
4570: douta=16'h6478;
4571: douta=16'h8d9b;
4572: douta=16'h7d3a;
4573: douta=16'h855b;
4574: douta=16'h7d3a;
4575: douta=16'h7d3b;
4576: douta=16'h7d5b;
4577: douta=16'h753a;
4578: douta=16'h8dbc;
4579: douta=16'h7d7b;
4580: douta=16'h7d7c;
4581: douta=16'h6cba;
4582: douta=16'h7d3a;
4583: douta=16'h74fa;
4584: douta=16'h74da;
4585: douta=16'h755b;
4586: douta=16'h753b;
4587: douta=16'h74b8;
4588: douta=16'h21a8;
4589: douta=16'h21a8;
4590: douta=16'h1107;
4591: douta=16'h1107;
4592: douta=16'h32af;
4593: douta=16'h8518;
4594: douta=16'h7455;
4595: douta=16'h63f5;
4596: douta=16'h1a0e;
4597: douta=16'h5373;
4598: douta=16'haddb;
4599: douta=16'hadfc;
4600: douta=16'h957a;
4601: douta=16'h2a90;
4602: douta=16'h2a70;
4603: douta=16'h5bb3;
4604: douta=16'h8518;
4605: douta=16'hbe3b;
4606: douta=16'h6416;
4607: douta=16'h8d5a;
4608: douta=16'h2a4f;
4609: douta=16'h1a0e;
4610: douta=16'h5374;
4611: douta=16'h74b9;
4612: douta=16'h6437;
4613: douta=16'h4b53;
4614: douta=16'h3a8e;
4615: douta=16'h2a2e;
4616: douta=16'h42f2;
4617: douta=16'h8475;
4618: douta=16'had97;
4619: douta=16'h8cb5;
4620: douta=16'h9453;
4621: douta=16'h8c75;
4622: douta=16'h63f4;
4623: douta=16'h9d15;
4624: douta=16'had36;
4625: douta=16'hbdf8;
4626: douta=16'hbdb7;
4627: douta=16'h6bf3;
4628: douta=16'h8412;
4629: douta=16'h5bb1;
4630: douta=16'hc5f7;
4631: douta=16'hde98;
4632: douta=16'hbdb6;
4633: douta=16'h7c33;
4634: douta=16'h94d4;
4635: douta=16'h8432;
4636: douta=16'hde98;
4637: douta=16'he6d9;
4638: douta=16'hbdb5;
4639: douta=16'hb595;
4640: douta=16'h94d3;
4641: douta=16'had13;
4642: douta=16'hd655;
4643: douta=16'hd677;
4644: douta=16'hde55;
4645: douta=16'h9430;
4646: douta=16'hbdd3;
4647: douta=16'h52ac;
4648: douta=16'h9c8e;
4649: douta=16'hb551;
4650: douta=16'h8bcc;
4651: douta=16'h6b4c;
4652: douta=16'hf779;
4653: douta=16'h9d12;
4654: douta=16'h41c7;
4655: douta=16'h2967;
4656: douta=16'h2967;
4657: douta=16'h2126;
4658: douta=16'h1926;
4659: douta=16'h1925;
4660: douta=16'h0042;
4661: douta=16'h3a4b;
4662: douta=16'h738e;
4663: douta=16'h9450;
4664: douta=16'had53;
4665: douta=16'h9430;
4666: douta=16'h42ac;
4667: douta=16'h83ee;
4668: douta=16'h5b2c;
4669: douta=16'h9cf2;
4670: douta=16'h63f3;
4671: douta=16'h29eb;
4672: douta=16'h5bb1;
4673: douta=16'h5350;
4674: douta=16'h4a8b;
4675: douta=16'h1883;
4676: douta=16'h18a2;
4677: douta=16'h18a3;
4678: douta=16'h0800;
4679: douta=16'h320b;
4680: douta=16'h21ea;
4681: douta=16'h21aa;
4682: douta=16'h3af0;
4683: douta=16'h4bb3;
4684: douta=16'h19ac;
4685: douta=16'h6435;
4686: douta=16'h4b93;
4687: douta=16'h7476;
4688: douta=16'h8559;
4689: douta=16'h5373;
4690: douta=16'h2a6f;
4691: douta=16'h84d6;
4692: douta=16'h7d19;
4693: douta=16'h6477;
4694: douta=16'h74b7;
4695: douta=16'h9d9a;
4696: douta=16'h5394;
4697: douta=16'h3b12;
4698: douta=16'h8475;
4699: douta=16'h5311;
4700: douta=16'h3aaf;
4701: douta=16'h6c35;
4702: douta=16'h6bf4;
4703: douta=16'ha5b9;
4704: douta=16'h4b31;
4705: douta=16'h428d;
4706: douta=16'h3168;
4707: douta=16'h39a8;
4708: douta=16'h20e5;
4709: douta=16'ha40e;
4710: douta=16'h6bb3;
4711: douta=16'h8518;
4712: douta=16'h7c97;
4713: douta=16'h7456;
4714: douta=16'h7c97;
4715: douta=16'h8d18;
4716: douta=16'h84f8;
4717: douta=16'h8519;
4718: douta=16'h7cb7;
4719: douta=16'h84f8;
4720: douta=16'h7c97;
4721: douta=16'h8519;
4722: douta=16'h74b8;
4723: douta=16'h7477;
4724: douta=16'h4b74;
4725: douta=16'h84f9;
4726: douta=16'h851a;
4727: douta=16'h957b;
4728: douta=16'h8519;
4729: douta=16'h7497;
4730: douta=16'h8d5a;
4731: douta=16'h7cb8;
4732: douta=16'h95bc;
4733: douta=16'h9dbc;
4734: douta=16'h957b;
4735: douta=16'h8d5b;
4736: douta=16'h8d3a;
4737: douta=16'h8d5a;
4738: douta=16'h8d5b;
4739: douta=16'h95bc;
4740: douta=16'h95bc;
4741: douta=16'h853a;
4742: douta=16'h8d7b;
4743: douta=16'h9dbc;
4744: douta=16'h95bc;
4745: douta=16'h6cb9;
4746: douta=16'h6c58;
4747: douta=16'h4353;
4748: douta=16'h6498;
4749: douta=16'h753b;
4750: douta=16'h53f7;
4751: douta=16'h74da;
4752: douta=16'h857c;
4753: douta=16'h7d3b;
4754: douta=16'h74da;
4755: douta=16'h74fa;
4756: douta=16'h7d3b;
4757: douta=16'h74da;
4758: douta=16'h74d9;
4759: douta=16'h859c;
4760: douta=16'h857b;
4761: douta=16'h7d5b;
4762: douta=16'h74fa;
4763: douta=16'h74d9;
4764: douta=16'h8d9b;
4765: douta=16'h6cd9;
4766: douta=16'h7d3b;
4767: douta=16'h74da;
4768: douta=16'h753a;
4769: douta=16'h7d3b;
4770: douta=16'h857b;
4771: douta=16'h8dbc;
4772: douta=16'h95dc;
4773: douta=16'h855b;
4774: douta=16'h6c99;
4775: douta=16'h857c;
4776: douta=16'h753b;
4777: douta=16'h6cda;
4778: douta=16'h753b;
4779: douta=16'h74b9;
4780: douta=16'h29e9;
4781: douta=16'h2147;
4782: douta=16'h1968;
4783: douta=16'h1148;
4784: douta=16'h08c6;
4785: douta=16'h21eb;
4786: douta=16'h84d7;
4787: douta=16'h8539;
4788: douta=16'h63f5;
4789: douta=16'h222f;
4790: douta=16'h53d4;
4791: douta=16'h5bf5;
4792: douta=16'h955a;
4793: douta=16'h84d7;
4794: douta=16'h5c16;
4795: douta=16'h2ab1;
4796: douta=16'h3b32;
4797: douta=16'ha5da;
4798: douta=16'h8d39;
4799: douta=16'h7cf9;
4800: douta=16'h32d1;
4801: douta=16'h32f2;
4802: douta=16'h4b73;
4803: douta=16'h8d9b;
4804: douta=16'h74b8;
4805: douta=16'h6436;
4806: douta=16'h5352;
4807: douta=16'h7456;
4808: douta=16'h6c36;
4809: douta=16'h6bf4;
4810: douta=16'h9d16;
4811: douta=16'h9cf6;
4812: douta=16'h8c74;
4813: douta=16'h8cb5;
4814: douta=16'h6bd2;
4815: douta=16'h6bd2;
4816: douta=16'hc5f8;
4817: douta=16'hd699;
4818: douta=16'h9453;
4819: douta=16'h6372;
4820: douta=16'h83f1;
4821: douta=16'h7c52;
4822: douta=16'hd677;
4823: douta=16'heed9;
4824: douta=16'ha514;
4825: douta=16'h7413;
4826: douta=16'h8c52;
4827: douta=16'h7c11;
4828: douta=16'he6b8;
4829: douta=16'he6d8;
4830: douta=16'h9cf3;
4831: douta=16'hb573;
4832: douta=16'h73b0;
4833: douta=16'ha553;
4834: douta=16'he6b6;
4835: douta=16'he719;
4836: douta=16'hd616;
4837: douta=16'h942f;
4838: douta=16'h8c4f;
4839: douta=16'h62eb;
4840: douta=16'h8c2e;
4841: douta=16'hdeb7;
4842: douta=16'h8bec;
4843: douta=16'h732b;
4844: douta=16'h6b2a;
4845: douta=16'h62aa;
4846: douta=16'h5249;
4847: douta=16'h2987;
4848: douta=16'h3a09;
4849: douta=16'h1906;
4850: douta=16'h1926;
4851: douta=16'h1905;
4852: douta=16'h10e4;
4853: douta=16'h0042;
4854: douta=16'h736d;
4855: douta=16'he717;
4856: douta=16'h73f0;
4857: douta=16'hb512;
4858: douta=16'h52aa;
4859: douta=16'h5b2c;
4860: douta=16'h18e4;
4861: douta=16'h324d;
4862: douta=16'h5bd3;
4863: douta=16'h328d;
4864: douta=16'h5351;
4865: douta=16'h5b6f;
4866: douta=16'h4b30;
4867: douta=16'ha5b7;
4868: douta=16'h39e9;
4869: douta=16'h2945;
4870: douta=16'h20e3;
4871: douta=16'h18e3;
4872: douta=16'h1082;
4873: douta=16'h3a2a;
4874: douta=16'h4aef;
4875: douta=16'h19ec;
4876: douta=16'h19ab;
4877: douta=16'h4bb5;
4878: douta=16'h5394;
4879: douta=16'h7c97;
4880: douta=16'h4b72;
4881: douta=16'h3aaf;
4882: douta=16'h3aaf;
4883: douta=16'h6477;
4884: douta=16'h53d5;
4885: douta=16'h53b4;
4886: douta=16'h9d38;
4887: douta=16'h4333;
4888: douta=16'h3270;
4889: douta=16'h63f4;
4890: douta=16'h53d4;
4891: douta=16'h6c76;
4892: douta=16'h6c36;
4893: douta=16'h63f4;
4894: douta=16'h9579;
4895: douta=16'h63f5;
4896: douta=16'h4a8c;
4897: douta=16'h4209;
4898: douta=16'h2127;
4899: douta=16'h934b;
4900: douta=16'h73f3;
4901: douta=16'h7496;
4902: douta=16'h955a;
4903: douta=16'h9d9a;
4904: douta=16'h84d7;
4905: douta=16'h7476;
4906: douta=16'h84d7;
4907: douta=16'h6c15;
4908: douta=16'h6c15;
4909: douta=16'h7c97;
4910: douta=16'h84d8;
4911: douta=16'h8d59;
4912: douta=16'h7cf8;
4913: douta=16'h7cb8;
4914: douta=16'h84f9;
4915: douta=16'h8d3a;
4916: douta=16'h7cb8;
4917: douta=16'h957a;
4918: douta=16'h8d5a;
4919: douta=16'h8d39;
4920: douta=16'h7d19;
4921: douta=16'h8d9b;
4922: douta=16'h853a;
4923: douta=16'h84f9;
4924: douta=16'h7cf9;
4925: douta=16'h8d5b;
4926: douta=16'h959c;
4927: douta=16'h7cf9;
4928: douta=16'h7cf9;
4929: douta=16'h8d5b;
4930: douta=16'h8d5b;
4931: douta=16'h8519;
4932: douta=16'h853a;
4933: douta=16'h8d5b;
4934: douta=16'h853a;
4935: douta=16'h8d5a;
4936: douta=16'h8539;
4937: douta=16'h8d7b;
4938: douta=16'h8d7b;
4939: douta=16'h8d7b;
4940: douta=16'h959c;
4941: douta=16'h74b9;
4942: douta=16'h53d6;
4943: douta=16'h5c58;
4944: douta=16'h6478;
4945: douta=16'h7d5b;
4946: douta=16'h6478;
4947: douta=16'h753b;
4948: douta=16'h7d3b;
4949: douta=16'h74da;
4950: douta=16'h857b;
4951: douta=16'h8dbc;
4952: douta=16'h6c99;
4953: douta=16'h6cfa;
4954: douta=16'h8dbc;
4955: douta=16'h751a;
4956: douta=16'h7d1a;
4957: douta=16'h74fa;
4958: douta=16'h7d3b;
4959: douta=16'h859c;
4960: douta=16'h7d7b;
4961: douta=16'h7d5b;
4962: douta=16'h751a;
4963: douta=16'h7d3b;
4964: douta=16'h8dbc;
4965: douta=16'h7d1a;
4966: douta=16'h8dbc;
4967: douta=16'h857b;
4968: douta=16'h6c78;
4969: douta=16'h74d9;
4970: douta=16'h859c;
4971: douta=16'h74da;
4972: douta=16'h753a;
4973: douta=16'h6cd9;
4974: douta=16'h7c98;
4975: douta=16'h29ca;
4976: douta=16'h1927;
4977: douta=16'h1948;
4978: douta=16'h5c37;
4979: douta=16'h5bf5;
4980: douta=16'h5394;
4981: douta=16'h1a4f;
4982: douta=16'ha579;
4983: douta=16'hc69d;
4984: douta=16'h6457;
4985: douta=16'h4bb5;
4986: douta=16'h5393;
4987: douta=16'h84f7;
4988: douta=16'h9559;
4989: douta=16'hadb9;
4990: douta=16'h6416;
4991: douta=16'h7cda;
4992: douta=16'h32f2;
4993: douta=16'h74d9;
4994: douta=16'h4312;
4995: douta=16'h74b9;
4996: douta=16'h3af1;
4997: douta=16'h2a70;
4998: douta=16'h5b93;
4999: douta=16'h7414;
5000: douta=16'h6bd4;
5001: douta=16'h8475;
5002: douta=16'h8cd5;
5003: douta=16'h6bd2;
5004: douta=16'h6b71;
5005: douta=16'hc5f8;
5006: douta=16'h8c94;
5007: douta=16'had56;
5008: douta=16'hc5f7;
5009: douta=16'h8453;
5010: douta=16'h8453;
5011: douta=16'hb555;
5012: douta=16'hd657;
5013: douta=16'h94b5;
5014: douta=16'h8cb5;
5015: douta=16'ha4d2;
5016: douta=16'had75;
5017: douta=16'hbdb4;
5018: douta=16'hf738;
5019: douta=16'ha4f2;
5020: douta=16'hf719;
5021: douta=16'hc5b5;
5022: douta=16'hce37;
5023: douta=16'hce14;
5024: douta=16'hde76;
5025: douta=16'hce76;
5026: douta=16'he6f9;
5027: douta=16'hce16;
5028: douta=16'h9c91;
5029: douta=16'hb531;
5030: douta=16'hb551;
5031: douta=16'had10;
5032: douta=16'hd5f4;
5033: douta=16'hde96;
5034: douta=16'h5269;
5035: douta=16'h732b;
5036: douta=16'h62ca;
5037: douta=16'h62a9;
5038: douta=16'h41e7;
5039: douta=16'h2167;
5040: douta=16'h2987;
5041: douta=16'h2968;
5042: douta=16'h2988;
5043: douta=16'h29a9;
5044: douta=16'h10c4;
5045: douta=16'h0084;
5046: douta=16'h39c7;
5047: douta=16'h9cf1;
5048: douta=16'h530c;
5049: douta=16'h6b4c;
5050: douta=16'hb552;
5051: douta=16'h7bce;
5052: douta=16'h634d;
5053: douta=16'h8d58;
5054: douta=16'h4b31;
5055: douta=16'h1148;
5056: douta=16'h3209;
5057: douta=16'h9472;
5058: douta=16'h84f7;
5059: douta=16'h53b3;
5060: douta=16'h4b0f;
5061: douta=16'h5bb2;
5062: douta=16'h31c7;
5063: douta=16'h1061;
5064: douta=16'h20e3;
5065: douta=16'h18e3;
5066: douta=16'h1061;
5067: douta=16'h1967;
5068: douta=16'h3b11;
5069: douta=16'h00e7;
5070: douta=16'h220c;
5071: douta=16'h3b11;
5072: douta=16'h3b31;
5073: douta=16'h53b4;
5074: douta=16'h6c33;
5075: douta=16'h29ec;
5076: douta=16'h5351;
5077: douta=16'h322c;
5078: douta=16'h4b31;
5079: douta=16'h5c15;
5080: douta=16'h53d5;
5081: douta=16'h74b8;
5082: douta=16'h6cb8;
5083: douta=16'h53d5;
5084: douta=16'h6bd2;
5085: douta=16'h7c96;
5086: douta=16'h4b10;
5087: douta=16'h52f0;
5088: douta=16'h4208;
5089: douta=16'h5a29;
5090: douta=16'h836c;
5091: douta=16'h528d;
5092: douta=16'h7476;
5093: douta=16'h9d9a;
5094: douta=16'h7c97;
5095: douta=16'h7cb7;
5096: douta=16'h9519;
5097: douta=16'h7cb7;
5098: douta=16'h8d18;
5099: douta=16'h7456;
5100: douta=16'h7456;
5101: douta=16'h7cb8;
5102: douta=16'h84d8;
5103: douta=16'h7c98;
5104: douta=16'h7cd8;
5105: douta=16'h84f9;
5106: douta=16'h7497;
5107: douta=16'h6c56;
5108: douta=16'h8d3a;
5109: douta=16'h7cd8;
5110: douta=16'h7cd8;
5111: douta=16'h8519;
5112: douta=16'h855a;
5113: douta=16'h7c98;
5114: douta=16'h7cb9;
5115: douta=16'h8d5a;
5116: douta=16'h851a;
5117: douta=16'h8d7b;
5118: douta=16'h8d7b;
5119: douta=16'h853a;
5120: douta=16'h853a;
5121: douta=16'h8d5a;
5122: douta=16'h8d7b;
5123: douta=16'h959c;
5124: douta=16'h9ddc;
5125: douta=16'h8d5a;
5126: douta=16'h8d7a;
5127: douta=16'h95bb;
5128: douta=16'h8d5a;
5129: douta=16'h8519;
5130: douta=16'h8d3a;
5131: douta=16'h959c;
5132: douta=16'h851a;
5133: douta=16'h959c;
5134: douta=16'h95bc;
5135: douta=16'h853a;
5136: douta=16'h6458;
5137: douta=16'h6c98;
5138: douta=16'h74fa;
5139: douta=16'h6478;
5140: douta=16'h7d5c;
5141: douta=16'h7d7b;
5142: douta=16'h857c;
5143: douta=16'h7d5b;
5144: douta=16'h8dbd;
5145: douta=16'h8d9c;
5146: douta=16'h6cba;
5147: douta=16'h95bc;
5148: douta=16'h857c;
5149: douta=16'h857c;
5150: douta=16'h7d3a;
5151: douta=16'h7d3b;
5152: douta=16'h855b;
5153: douta=16'h74fa;
5154: douta=16'h753b;
5155: douta=16'h751a;
5156: douta=16'h6499;
5157: douta=16'h751a;
5158: douta=16'h8dbc;
5159: douta=16'h74d9;
5160: douta=16'h74fa;
5161: douta=16'h74d9;
5162: douta=16'h5c16;
5163: douta=16'h753a;
5164: douta=16'h74b9;
5165: douta=16'h6cb9;
5166: douta=16'h6cfa;
5167: douta=16'h5b53;
5168: douta=16'h29a8;
5169: douta=16'h2188;
5170: douta=16'h1148;
5171: douta=16'h53d4;
5172: douta=16'h9538;
5173: douta=16'h84f8;
5174: douta=16'h5c16;
5175: douta=16'h32b0;
5176: douta=16'h3ad1;
5177: douta=16'h5392;
5178: douta=16'h8d17;
5179: douta=16'h53b4;
5180: douta=16'h7456;
5181: douta=16'h3b12;
5182: douta=16'h74d8;
5183: douta=16'h84d7;
5184: douta=16'h2ad0;
5185: douta=16'h4333;
5186: douta=16'h53f5;
5187: douta=16'h7d3b;
5188: douta=16'h6477;
5189: douta=16'h74da;
5190: douta=16'h5352;
5191: douta=16'h5353;
5192: douta=16'h4b31;
5193: douta=16'h5331;
5194: douta=16'had77;
5195: douta=16'h9d17;
5196: douta=16'h8c74;
5197: douta=16'h7433;
5198: douta=16'h6bd2;
5199: douta=16'h8cb5;
5200: douta=16'hbd96;
5201: douta=16'he6fa;
5202: douta=16'h8c74;
5203: douta=16'hb575;
5204: douta=16'hc5d6;
5205: douta=16'h73f2;
5206: douta=16'hce16;
5207: douta=16'hde97;
5208: douta=16'hde98;
5209: douta=16'h8c31;
5210: douta=16'hc5b5;
5211: douta=16'h8c51;
5212: douta=16'hdeb8;
5213: douta=16'he6b8;
5214: douta=16'hd637;
5215: douta=16'hc5f4;
5216: douta=16'he6f8;
5217: douta=16'ha4d0;
5218: douta=16'hce14;
5219: douta=16'hce35;
5220: douta=16'heeb7;
5221: douta=16'hbd12;
5222: douta=16'h94af;
5223: douta=16'h946f;
5224: douta=16'hcd93;
5225: douta=16'hf759;
5226: douta=16'h732b;
5227: douta=16'h732a;
5228: douta=16'h62ca;
5229: douta=16'h5a68;
5230: douta=16'h4208;
5231: douta=16'h1926;
5232: douta=16'h18e5;
5233: douta=16'h10e4;
5234: douta=16'h1905;
5235: douta=16'h2968;
5236: douta=16'h10e5;
5237: douta=16'h1105;
5238: douta=16'h0883;
5239: douta=16'hbdf5;
5240: douta=16'h322a;
5241: douta=16'h83ad;
5242: douta=16'h5aaa;
5243: douta=16'h6baf;
5244: douta=16'h7c53;
5245: douta=16'h74b5;
5246: douta=16'h5b4e;
5247: douta=16'h21a9;
5248: douta=16'h10a5;
5249: douta=16'h8c30;
5250: douta=16'h7cb6;
5251: douta=16'h4310;
5252: douta=16'h52ee;
5253: douta=16'h5330;
5254: douta=16'h94f5;
5255: douta=16'h1926;
5256: douta=16'h18a2;
5257: douta=16'h1082;
5258: douta=16'h10a2;
5259: douta=16'h0000;
5260: douta=16'h4b11;
5261: douta=16'h2a0d;
5262: douta=16'h1149;
5263: douta=16'h4bb5;
5264: douta=16'h53d5;
5265: douta=16'h2a4e;
5266: douta=16'h63d4;
5267: douta=16'h5392;
5268: douta=16'h5bd4;
5269: douta=16'h5b91;
5270: douta=16'h4b72;
5271: douta=16'h4332;
5272: douta=16'h53d5;
5273: douta=16'h6436;
5274: douta=16'h5c57;
5275: douta=16'h5c16;
5276: douta=16'h9579;
5277: douta=16'h8dbc;
5278: douta=16'h63b2;
5279: douta=16'h4a09;
5280: douta=16'h4229;
5281: douta=16'hc4cf;
5282: douta=16'h5a6c;
5283: douta=16'h8454;
5284: douta=16'h6bd4;
5285: douta=16'hadfb;
5286: douta=16'h9559;
5287: douta=16'h63f4;
5288: douta=16'h7c96;
5289: douta=16'h957a;
5290: douta=16'h6c15;
5291: douta=16'h9559;
5292: douta=16'h8d18;
5293: douta=16'h8d39;
5294: douta=16'h8d19;
5295: douta=16'h84d8;
5296: douta=16'h6c57;
5297: douta=16'h84f9;
5298: douta=16'h957a;
5299: douta=16'h84f9;
5300: douta=16'h5bd5;
5301: douta=16'h957a;
5302: douta=16'h84f8;
5303: douta=16'h8d5a;
5304: douta=16'h853a;
5305: douta=16'h8d5a;
5306: douta=16'h7498;
5307: douta=16'h7498;
5308: douta=16'h853a;
5309: douta=16'h7cf9;
5310: douta=16'h959c;
5311: douta=16'h8d7b;
5312: douta=16'h853a;
5313: douta=16'h8d7b;
5314: douta=16'h855a;
5315: douta=16'h8d5b;
5316: douta=16'h8d7b;
5317: douta=16'h959b;
5318: douta=16'h853a;
5319: douta=16'h957b;
5320: douta=16'ha5dc;
5321: douta=16'h851a;
5322: douta=16'h851a;
5323: douta=16'h853a;
5324: douta=16'h8d7b;
5325: douta=16'h8d5a;
5326: douta=16'h95bc;
5327: douta=16'h95bc;
5328: douta=16'h8d9b;
5329: douta=16'h5bf6;
5330: douta=16'h751a;
5331: douta=16'h7d5b;
5332: douta=16'h6cfa;
5333: douta=16'h7d3b;
5334: douta=16'h6cba;
5335: douta=16'h7d5c;
5336: douta=16'h859c;
5337: douta=16'h7d7b;
5338: douta=16'h8d9c;
5339: douta=16'h74fb;
5340: douta=16'h857b;
5341: douta=16'h8d9c;
5342: douta=16'h7d3b;
5343: douta=16'h7d3b;
5344: douta=16'h857b;
5345: douta=16'h7d3b;
5346: douta=16'h6cb9;
5347: douta=16'h85bc;
5348: douta=16'h857b;
5349: douta=16'h6cda;
5350: douta=16'h8dbc;
5351: douta=16'h7d3a;
5352: douta=16'h7499;
5353: douta=16'h855b;
5354: douta=16'h6437;
5355: douta=16'h6478;
5356: douta=16'h8dbc;
5357: douta=16'h7d3b;
5358: douta=16'h7d1a;
5359: douta=16'h74fa;
5360: douta=16'h31ea;
5361: douta=16'h31a8;
5362: douta=16'h1967;
5363: douta=16'h1968;
5364: douta=16'h5c16;
5365: douta=16'ha5ba;
5366: douta=16'h7497;
5367: douta=16'h7cb8;
5368: douta=16'h5351;
5369: douta=16'h1a0e;
5370: douta=16'h7cb7;
5371: douta=16'h84b7;
5372: douta=16'hb63b;
5373: douta=16'h6c55;
5374: douta=16'h1a50;
5375: douta=16'h8d39;
5376: douta=16'h32f2;
5377: douta=16'h32f1;
5378: douta=16'h5c37;
5379: douta=16'h53b4;
5380: douta=16'h6436;
5381: douta=16'h6c98;
5382: douta=16'h6c15;
5383: douta=16'h4b11;
5384: douta=16'h4311;
5385: douta=16'h5b72;
5386: douta=16'h94d6;
5387: douta=16'h9d17;
5388: douta=16'h73d3;
5389: douta=16'h8c95;
5390: douta=16'had98;
5391: douta=16'h6bd4;
5392: douta=16'hd637;
5393: douta=16'hbdb6;
5394: douta=16'h8c73;
5395: douta=16'h73f2;
5396: douta=16'h7391;
5397: douta=16'h7c10;
5398: douta=16'hd657;
5399: douta=16'hde77;
5400: douta=16'h9cb2;
5401: douta=16'hb554;
5402: douta=16'hd636;
5403: douta=16'h83ef;
5404: douta=16'hc5f5;
5405: douta=16'hef39;
5406: douta=16'hf75a;
5407: douta=16'he676;
5408: douta=16'hc5d3;
5409: douta=16'ha48f;
5410: douta=16'hef19;
5411: douta=16'he6d8;
5412: douta=16'hb532;
5413: douta=16'h6289;
5414: douta=16'hd675;
5415: douta=16'h5aca;
5416: douta=16'h83ab;
5417: douta=16'h730a;
5418: douta=16'h83ab;
5419: douta=16'h6b2b;
5420: douta=16'h62c9;
5421: douta=16'h5a69;
5422: douta=16'h2986;
5423: douta=16'h10c4;
5424: douta=16'h2125;
5425: douta=16'h10e5;
5426: douta=16'h10e4;
5427: douta=16'h10e5;
5428: douta=16'h1126;
5429: douta=16'h10e5;
5430: douta=16'h0884;
5431: douta=16'h42ab;
5432: douta=16'h4a29;
5433: douta=16'h7bad;
5434: douta=16'h6b4e;
5435: douta=16'h5371;
5436: douta=16'h5b50;
5437: douta=16'h4a6b;
5438: douta=16'h6bf2;
5439: douta=16'h3a29;
5440: douta=16'h4a6a;
5441: douta=16'had33;
5442: douta=16'h1906;
5443: douta=16'h4b51;
5444: douta=16'h6371;
5445: douta=16'h3aae;
5446: douta=16'h5bd3;
5447: douta=16'h3a6d;
5448: douta=16'h21ca;
5449: douta=16'h3a09;
5450: douta=16'h1041;
5451: douta=16'h18a2;
5452: douta=16'h0861;
5453: douta=16'h0000;
5454: douta=16'h0000;
5455: douta=16'h2a4e;
5456: douta=16'h32d1;
5457: douta=16'h1149;
5458: douta=16'h53f5;
5459: douta=16'h53b3;
5460: douta=16'h53d5;
5461: douta=16'h5351;
5462: douta=16'h32d0;
5463: douta=16'h19ed;
5464: douta=16'h63f4;
5465: douta=16'h7d1a;
5466: douta=16'h74b8;
5467: douta=16'h5c16;
5468: douta=16'h7d19;
5469: douta=16'h6cb9;
5470: douta=16'h422a;
5471: douta=16'h39c7;
5472: douta=16'ha42d;
5473: douta=16'h84d7;
5474: douta=16'h8d59;
5475: douta=16'h8497;
5476: douta=16'h8cd8;
5477: douta=16'h84f8;
5478: douta=16'h5bf5;
5479: douta=16'h6c36;
5480: douta=16'h84f9;
5481: douta=16'h84f9;
5482: douta=16'h7c97;
5483: douta=16'h7c97;
5484: douta=16'h6c35;
5485: douta=16'h8d39;
5486: douta=16'h8d39;
5487: douta=16'h6c36;
5488: douta=16'h7c97;
5489: douta=16'h955a;
5490: douta=16'h8d7a;
5491: douta=16'h7c77;
5492: douta=16'h6c56;
5493: douta=16'h7c98;
5494: douta=16'h8519;
5495: douta=16'h8519;
5496: douta=16'h6c56;
5497: douta=16'h6c36;
5498: douta=16'h5bf5;
5499: douta=16'h6c57;
5500: douta=16'h8d5a;
5501: douta=16'h8d7a;
5502: douta=16'h853a;
5503: douta=16'h9dbc;
5504: douta=16'h8d5b;
5505: douta=16'h7cd9;
5506: douta=16'h959b;
5507: douta=16'h959c;
5508: douta=16'h95bc;
5509: douta=16'h8d7b;
5510: douta=16'h853a;
5511: douta=16'h8d5a;
5512: douta=16'h851a;
5513: douta=16'h8d5b;
5514: douta=16'h957b;
5515: douta=16'h959b;
5516: douta=16'h959b;
5517: douta=16'h95bc;
5518: douta=16'h7d19;
5519: douta=16'h8d5b;
5520: douta=16'h8d5a;
5521: douta=16'h8d9b;
5522: douta=16'h95bc;
5523: douta=16'h9ddc;
5524: douta=16'h7d3b;
5525: douta=16'h961d;
5526: douta=16'h6cba;
5527: douta=16'h751b;
5528: douta=16'h6cba;
5529: douta=16'h7d3b;
5530: douta=16'h753b;
5531: douta=16'h7d5b;
5532: douta=16'h855c;
5533: douta=16'h857c;
5534: douta=16'h74fa;
5535: douta=16'h74fa;
5536: douta=16'h857b;
5537: douta=16'h74fa;
5538: douta=16'h751b;
5539: douta=16'h857b;
5540: douta=16'h7d3b;
5541: douta=16'h6cba;
5542: douta=16'h857c;
5543: douta=16'h7d3b;
5544: douta=16'h6c98;
5545: douta=16'h74f9;
5546: douta=16'h855b;
5547: douta=16'h8dbc;
5548: douta=16'h6499;
5549: douta=16'h6499;
5550: douta=16'h6478;
5551: douta=16'h751b;
5552: douta=16'h7d7c;
5553: douta=16'h74fa;
5554: douta=16'h29ca;
5555: douta=16'h1968;
5556: douta=16'h1106;
5557: douta=16'h53d4;
5558: douta=16'h32d1;
5559: douta=16'h32d0;
5560: douta=16'h2ab1;
5561: douta=16'hadda;
5562: douta=16'h5bd4;
5563: douta=16'h8519;
5564: douta=16'h6435;
5565: douta=16'h63d4;
5566: douta=16'h4353;
5567: douta=16'h322c;
5568: douta=16'h2ab0;
5569: douta=16'h4374;
5570: douta=16'h5c57;
5571: douta=16'h326f;
5572: douta=16'h4b52;
5573: douta=16'h5bd5;
5574: douta=16'h7c76;
5575: douta=16'h8497;
5576: douta=16'h9d59;
5577: douta=16'h84d7;
5578: douta=16'h4ad0;
5579: douta=16'h5b70;
5580: douta=16'h5b30;
5581: douta=16'ha536;
5582: douta=16'hce39;
5583: douta=16'hb5b8;
5584: douta=16'h8c93;
5585: douta=16'had35;
5586: douta=16'h3a4d;
5587: douta=16'hc5f6;
5588: douta=16'hde77;
5589: douta=16'had75;
5590: douta=16'had56;
5591: douta=16'h6b4d;
5592: douta=16'h9cb2;
5593: douta=16'hc5f6;
5594: douta=16'hde76;
5595: douta=16'ha4d1;
5596: douta=16'h8bf0;
5597: douta=16'h52ed;
5598: douta=16'h8c0f;
5599: douta=16'h9c6f;
5600: douta=16'hbdd3;
5601: douta=16'hde97;
5602: douta=16'ha4d1;
5603: douta=16'hd636;
5604: douta=16'h736c;
5605: douta=16'hc593;
5606: douta=16'hc614;
5607: douta=16'hb572;
5608: douta=16'h836b;
5609: douta=16'h83ac;
5610: douta=16'h836b;
5611: douta=16'h836b;
5612: douta=16'h62a9;
5613: douta=16'h5a68;
5614: douta=16'h31c8;
5615: douta=16'h2167;
5616: douta=16'h10c5;
5617: douta=16'h10a4;
5618: douta=16'h10e5;
5619: douta=16'h10a4;
5620: douta=16'h10e4;
5621: douta=16'h18e5;
5622: douta=16'h10e4;
5623: douta=16'h31e9;
5624: douta=16'h39a8;
5625: douta=16'h9cf1;
5626: douta=16'h63d1;
5627: douta=16'h63d2;
5628: douta=16'h6c33;
5629: douta=16'h1927;
5630: douta=16'h1927;
5631: douta=16'h638e;
5632: douta=16'h4a4a;
5633: douta=16'h8430;
5634: douta=16'h5acc;
5635: douta=16'h10e6;
5636: douta=16'h8474;
5637: douta=16'h3a8e;
5638: douta=16'h4b0f;
5639: douta=16'h5370;
5640: douta=16'h4b31;
5641: douta=16'h3a8f;
5642: douta=16'h5393;
5643: douta=16'h3aaf;
5644: douta=16'h1081;
5645: douta=16'h10e3;
5646: douta=16'h18e4;
5647: douta=16'h1926;
5648: douta=16'h428d;
5649: douta=16'h5330;
5650: douta=16'h1169;
5651: douta=16'h4374;
5652: douta=16'h3b32;
5653: douta=16'h4b11;
5654: douta=16'h3b11;
5655: douta=16'h4312;
5656: douta=16'h7cd8;
5657: douta=16'h53b4;
5658: douta=16'h74b8;
5659: douta=16'h3a4e;
5660: douta=16'h6498;
5661: douta=16'h5372;
5662: douta=16'hc48e;
5663: douta=16'hacaf;
5664: douta=16'h94b6;
5665: douta=16'h957b;
5666: douta=16'h6478;
5667: douta=16'h4bd6;
5668: douta=16'h9dbb;
5669: douta=16'h957a;
5670: douta=16'h7498;
5671: douta=16'h5bf5;
5672: douta=16'h5bb5;
5673: douta=16'h6c56;
5674: douta=16'h7cb8;
5675: douta=16'h7c76;
5676: douta=16'h7476;
5677: douta=16'h6415;
5678: douta=16'h6c36;
5679: douta=16'h5bd4;
5680: douta=16'h95dc;
5681: douta=16'h8d1a;
5682: douta=16'h7cb8;
5683: douta=16'h8539;
5684: douta=16'h959b;
5685: douta=16'h84d8;
5686: douta=16'h6c16;
5687: douta=16'h7cb8;
5688: douta=16'h84d8;
5689: douta=16'h6415;
5690: douta=16'h6c56;
5691: douta=16'h63f5;
5692: douta=16'h7cf9;
5693: douta=16'h851a;
5694: douta=16'h853a;
5695: douta=16'h8d5a;
5696: douta=16'h8d7a;
5697: douta=16'h853a;
5698: douta=16'h851a;
5699: douta=16'h7cd9;
5700: douta=16'h853a;
5701: douta=16'h9ddc;
5702: douta=16'h8d5a;
5703: douta=16'h7cd9;
5704: douta=16'h8d3a;
5705: douta=16'h8d3a;
5706: douta=16'h8d5a;
5707: douta=16'h8d7b;
5708: douta=16'h8d3a;
5709: douta=16'h8d7b;
5710: douta=16'h8d3a;
5711: douta=16'h8d5b;
5712: douta=16'h959b;
5713: douta=16'h851a;
5714: douta=16'h851a;
5715: douta=16'h853a;
5716: douta=16'h8d7b;
5717: douta=16'h855a;
5718: douta=16'h855c;
5719: douta=16'h5417;
5720: douta=16'h8e1e;
5721: douta=16'h9e3e;
5722: douta=16'h5c58;
5723: douta=16'h6cfa;
5724: douta=16'h6cba;
5725: douta=16'h7d3b;
5726: douta=16'h857c;
5727: douta=16'h7d3b;
5728: douta=16'h7d1a;
5729: douta=16'h857b;
5730: douta=16'h857b;
5731: douta=16'h74ba;
5732: douta=16'h74fa;
5733: douta=16'h7d3a;
5734: douta=16'h6cb9;
5735: douta=16'h6458;
5736: douta=16'h74da;
5737: douta=16'h74f9;
5738: douta=16'h8d5b;
5739: douta=16'h7d3b;
5740: douta=16'h6cd9;
5741: douta=16'h6cfa;
5742: douta=16'h7d5c;
5743: douta=16'h5c58;
5744: douta=16'h74fa;
5745: douta=16'h7d3b;
5746: douta=16'h31ea;
5747: douta=16'h1906;
5748: douta=16'h2989;
5749: douta=16'h957a;
5750: douta=16'h5353;
5751: douta=16'h9559;
5752: douta=16'h9d7a;
5753: douta=16'h19cc;
5754: douta=16'h84d7;
5755: douta=16'h3290;
5756: douta=16'h4b51;
5757: douta=16'h7433;
5758: douta=16'ha597;
5759: douta=16'h42d0;
5760: douta=16'h3b53;
5761: douta=16'h32d1;
5762: douta=16'h74fa;
5763: douta=16'h5373;
5764: douta=16'h5bb4;
5765: douta=16'h6436;
5766: douta=16'h5373;
5767: douta=16'h5351;
5768: douta=16'h8cf8;
5769: douta=16'h7c96;
5770: douta=16'h9d16;
5771: douta=16'h9cf5;
5772: douta=16'h6392;
5773: douta=16'h8c94;
5774: douta=16'hbdf9;
5775: douta=16'h8454;
5776: douta=16'hce38;
5777: douta=16'hcdf6;
5778: douta=16'h8c53;
5779: douta=16'had55;
5780: douta=16'had34;
5781: douta=16'h9cd3;
5782: douta=16'hd637;
5783: douta=16'hee98;
5784: douta=16'hef39;
5785: douta=16'h83ef;
5786: douta=16'hc5d4;
5787: douta=16'hb593;
5788: douta=16'heed8;
5789: douta=16'hbd52;
5790: douta=16'he697;
5791: douta=16'h6269;
5792: douta=16'h8cd1;
5793: douta=16'hcdf3;
5794: douta=16'heef8;
5795: douta=16'hdeb7;
5796: douta=16'hc592;
5797: douta=16'hac91;
5798: douta=16'h94cf;
5799: douta=16'h736c;
5800: douta=16'h8b8c;
5801: douta=16'h8bac;
5802: douta=16'h838b;
5803: douta=16'h7b2a;
5804: douta=16'h62a9;
5805: douta=16'h4a49;
5806: douta=16'h4a6b;
5807: douta=16'h320a;
5808: douta=16'h29a8;
5809: douta=16'h1905;
5810: douta=16'h10e4;
5811: douta=16'h18e5;
5812: douta=16'h10c4;
5813: douta=16'h1105;
5814: douta=16'h10e4;
5815: douta=16'h4a8a;
5816: douta=16'h528a;
5817: douta=16'h8c70;
5818: douta=16'h63b1;
5819: douta=16'h63d2;
5820: douta=16'h5b6f;
5821: douta=16'h7bae;
5822: douta=16'h2189;
5823: douta=16'h73d0;
5824: douta=16'h2189;
5825: douta=16'h3209;
5826: douta=16'h528b;
5827: douta=16'h29aa;
5828: douta=16'h6bf1;
5829: douta=16'h2a2c;
5830: douta=16'h5371;
5831: douta=16'h6391;
5832: douta=16'h21cb;
5833: douta=16'h5330;
5834: douta=16'h63d2;
5835: douta=16'h53f6;
5836: douta=16'h2986;
5837: douta=16'h10a3;
5838: douta=16'h18e4;
5839: douta=16'h0841;
5840: douta=16'h0021;
5841: douta=16'h4aef;
5842: douta=16'h00a6;
5843: douta=16'h2a8f;
5844: douta=16'h4311;
5845: douta=16'h5bd5;
5846: douta=16'h3b32;
5847: douta=16'h00e9;
5848: douta=16'h4b32;
5849: douta=16'h3af1;
5850: douta=16'h6497;
5851: douta=16'h6436;
5852: douta=16'h5bd4;
5853: douta=16'h5228;
5854: douta=16'hacce;
5855: douta=16'h41e8;
5856: douta=16'h9ddd;
5857: douta=16'h8d5b;
5858: douta=16'h8d7b;
5859: douta=16'h7cd9;
5860: douta=16'h7498;
5861: douta=16'h959b;
5862: douta=16'h9ddc;
5863: douta=16'h6c36;
5864: douta=16'h5bd5;
5865: douta=16'h6c57;
5866: douta=16'h8d39;
5867: douta=16'h84f9;
5868: douta=16'h7cb8;
5869: douta=16'h84d8;
5870: douta=16'h8d19;
5871: douta=16'h7c98;
5872: douta=16'h6c36;
5873: douta=16'h9ddb;
5874: douta=16'ha61c;
5875: douta=16'h7cb8;
5876: douta=16'h84d9;
5877: douta=16'h8d5a;
5878: douta=16'h84d8;
5879: douta=16'h7cb8;
5880: douta=16'h7477;
5881: douta=16'h7cd8;
5882: douta=16'h7457;
5883: douta=16'h63f5;
5884: douta=16'h6416;
5885: douta=16'h6c57;
5886: douta=16'h8519;
5887: douta=16'h8519;
5888: douta=16'h8539;
5889: douta=16'h8519;
5890: douta=16'h8519;
5891: douta=16'h7cf9;
5892: douta=16'h7cf9;
5893: douta=16'h8d5b;
5894: douta=16'h9ddc;
5895: douta=16'h959b;
5896: douta=16'h851a;
5897: douta=16'h8519;
5898: douta=16'h957a;
5899: douta=16'h851a;
5900: douta=16'h957b;
5901: douta=16'h8d3a;
5902: douta=16'h8519;
5903: douta=16'h8d3a;
5904: douta=16'h8d7b;
5905: douta=16'h8d5b;
5906: douta=16'h851a;
5907: douta=16'h851a;
5908: douta=16'h8d5b;
5909: douta=16'h8d7c;
5910: douta=16'h959c;
5911: douta=16'h53d7;
5912: douta=16'h4bd6;
5913: douta=16'h751a;
5914: douta=16'h8d9c;
5915: douta=16'h6cfa;
5916: douta=16'h6cda;
5917: douta=16'h7d5b;
5918: douta=16'h859c;
5919: douta=16'h6cda;
5920: douta=16'h855b;
5921: douta=16'h857b;
5922: douta=16'h855b;
5923: douta=16'h6478;
5924: douta=16'h74b9;
5925: douta=16'h751a;
5926: douta=16'h74d9;
5927: douta=16'h74d9;
5928: douta=16'h74b9;
5929: douta=16'h8dbc;
5930: douta=16'h8dbc;
5931: douta=16'h8d9c;
5932: douta=16'h751a;
5933: douta=16'h6cd9;
5934: douta=16'h859b;
5935: douta=16'h74fb;
5936: douta=16'h6478;
5937: douta=16'h6457;
5938: douta=16'h7457;
5939: douta=16'h29a9;
5940: douta=16'h2189;
5941: douta=16'h2a8f;
5942: douta=16'h4b51;
5943: douta=16'h6c15;
5944: douta=16'hae1c;
5945: douta=16'h7435;
5946: douta=16'h84d7;
5947: douta=16'h5393;
5948: douta=16'h0969;
5949: douta=16'h3a8d;
5950: douta=16'h326e;
5951: douta=16'h6371;
5952: douta=16'h3312;
5953: douta=16'h2a4f;
5954: douta=16'h4312;
5955: douta=16'h5bf5;
5956: douta=16'h7cf9;
5957: douta=16'h4b53;
5958: douta=16'h5393;
5959: douta=16'h5b72;
5960: douta=16'h84d7;
5961: douta=16'h7c96;
5962: douta=16'h94b5;
5963: douta=16'h73f2;
5964: douta=16'h73f2;
5965: douta=16'h94d5;
5966: douta=16'hadb7;
5967: douta=16'h8c94;
5968: douta=16'hc5d6;
5969: douta=16'hb554;
5970: douta=16'h6b70;
5971: douta=16'hb535;
5972: douta=16'hbdd6;
5973: douta=16'h9cd3;
5974: douta=16'hce36;
5975: douta=16'hc574;
5976: douta=16'hf6d8;
5977: douta=16'h736e;
5978: douta=16'h83d0;
5979: douta=16'had32;
5980: douta=16'hd636;
5981: douta=16'ha4d1;
5982: douta=16'hc593;
5983: douta=16'h6aeb;
5984: douta=16'h532c;
5985: douta=16'hb551;
5986: douta=16'hf718;
5987: douta=16'hef39;
5988: douta=16'h9caf;
5989: douta=16'h7b8c;
5990: douta=16'h8b8c;
5991: douta=16'h838c;
5992: douta=16'h836b;
5993: douta=16'h8bcc;
5994: douta=16'h93cc;
5995: douta=16'h8bac;
5996: douta=16'h5248;
5997: douta=16'h31a7;
5998: douta=16'h18e5;
5999: douta=16'h2146;
6000: douta=16'h1906;
6001: douta=16'h3a08;
6002: douta=16'h10c5;
6003: douta=16'h10e5;
6004: douta=16'h10e5;
6005: douta=16'h10c4;
6006: douta=16'h10e5;
6007: douta=16'h39c8;
6008: douta=16'h2125;
6009: douta=16'h9c8f;
6010: douta=16'h5b72;
6011: douta=16'h5b71;
6012: douta=16'h9cb0;
6013: douta=16'h6b6e;
6014: douta=16'h1107;
6015: douta=16'h4acd;
6016: douta=16'h73cf;
6017: douta=16'h4aac;
6018: douta=16'h5aec;
6019: douta=16'h6b6e;
6020: douta=16'h29ca;
6021: douta=16'h52ac;
6022: douta=16'h4acd;
6023: douta=16'h426d;
6024: douta=16'h5b4f;
6025: douta=16'h5bb3;
6026: douta=16'h6c14;
6027: douta=16'h4373;
6028: douta=16'h4b11;
6029: douta=16'h2a2d;
6030: douta=16'h2a2e;
6031: douta=16'h1061;
6032: douta=16'h1082;
6033: douta=16'h0001;
6034: douta=16'h0000;
6035: douta=16'h5b50;
6036: douta=16'h4aef;
6037: douta=16'h224f;
6038: douta=16'h222d;
6039: douta=16'h5bb4;
6040: douta=16'h2a8f;
6041: douta=16'h326f;
6042: douta=16'h53f5;
6043: douta=16'h5b50;
6044: douta=16'h39e9;
6045: douta=16'h830a;
6046: douta=16'h9dfd;
6047: douta=16'h9ddc;
6048: douta=16'h8d7a;
6049: douta=16'h959b;
6050: douta=16'ha5dc;
6051: douta=16'ha5fc;
6052: douta=16'h8519;
6053: douta=16'h7cf9;
6054: douta=16'h853a;
6055: douta=16'h8d7b;
6056: douta=16'h957b;
6057: douta=16'h8d7b;
6058: douta=16'h8519;
6059: douta=16'h8d3a;
6060: douta=16'h8519;
6061: douta=16'h7497;
6062: douta=16'h84f8;
6063: douta=16'h8519;
6064: douta=16'h8d5a;
6065: douta=16'h74b8;
6066: douta=16'h855a;
6067: douta=16'h7cd9;
6068: douta=16'h853a;
6069: douta=16'h95bb;
6070: douta=16'h6c15;
6071: douta=16'h7476;
6072: douta=16'h8d5a;
6073: douta=16'h8519;
6074: douta=16'h7478;
6075: douta=16'h7498;
6076: douta=16'h8d5a;
6077: douta=16'h8d5a;
6078: douta=16'h7457;
6079: douta=16'h7cb8;
6080: douta=16'h7cf9;
6081: douta=16'h6c36;
6082: douta=16'h959b;
6083: douta=16'h8d7b;
6084: douta=16'h8d7b;
6085: douta=16'h8d7b;
6086: douta=16'h8d7b;
6087: douta=16'h8d7b;
6088: douta=16'h9ddc;
6089: douta=16'h95bb;
6090: douta=16'h8d7b;
6091: douta=16'h8d3a;
6092: douta=16'h957b;
6093: douta=16'h74b8;
6094: douta=16'h8519;
6095: douta=16'h8d5b;
6096: douta=16'h8d7b;
6097: douta=16'h8d5a;
6098: douta=16'h8d7b;
6099: douta=16'h959c;
6100: douta=16'h7d1a;
6101: douta=16'h855b;
6102: douta=16'h95bc;
6103: douta=16'h8d7b;
6104: douta=16'h855b;
6105: douta=16'h95bc;
6106: douta=16'h4b11;
6107: douta=16'h3b33;
6108: douta=16'h7d3b;
6109: douta=16'h6458;
6110: douta=16'h6438;
6111: douta=16'h53d6;
6112: douta=16'h6cd9;
6113: douta=16'h6cb9;
6114: douta=16'h74fa;
6115: douta=16'h855b;
6116: douta=16'h8dbc;
6117: douta=16'h751a;
6118: douta=16'h6c99;
6119: douta=16'h74d9;
6120: douta=16'h7d3a;
6121: douta=16'h7d1a;
6122: douta=16'h7d1a;
6123: douta=16'h855b;
6124: douta=16'h7d1a;
6125: douta=16'h6cb9;
6126: douta=16'h95bc;
6127: douta=16'h6cba;
6128: douta=16'h6478;
6129: douta=16'h6c98;
6130: douta=16'h6c97;
6131: douta=16'h6c77;
6132: douta=16'h4acf;
6133: douta=16'h2189;
6134: douta=16'h7cb7;
6135: douta=16'hcebd;
6136: douta=16'hc65b;
6137: douta=16'h5bd4;
6138: douta=16'h3aaf;
6139: douta=16'h63d2;
6140: douta=16'had77;
6141: douta=16'ha536;
6142: douta=16'h3ad0;
6143: douta=16'h4af0;
6144: douta=16'h4bb6;
6145: douta=16'h3b33;
6146: douta=16'h4333;
6147: douta=16'h5394;
6148: douta=16'h326f;
6149: douta=16'h322e;
6150: douta=16'h4311;
6151: douta=16'h5b93;
6152: douta=16'h84b7;
6153: douta=16'h8d39;
6154: douta=16'h6bf3;
6155: douta=16'h7c35;
6156: douta=16'h5b70;
6157: douta=16'hd659;
6158: douta=16'hd69b;
6159: douta=16'hb5f8;
6160: douta=16'h9472;
6161: douta=16'hbd95;
6162: douta=16'h8451;
6163: douta=16'hd637;
6164: douta=16'hde97;
6165: douta=16'had34;
6166: douta=16'ha512;
6167: douta=16'h5aed;
6168: douta=16'h83ae;
6169: douta=16'hc5f4;
6170: douta=16'hbd94;
6171: douta=16'hc5d4;
6172: douta=16'hacd1;
6173: douta=16'h8c4f;
6174: douta=16'hde56;
6175: douta=16'hc5b3;
6176: douta=16'hb530;
6177: douta=16'hff9b;
6178: douta=16'ha4b0;
6179: douta=16'hbd93;
6180: douta=16'h7bcd;
6181: douta=16'h836b;
6182: douta=16'h8bcc;
6183: douta=16'h93ec;
6184: douta=16'h8bab;
6185: douta=16'h9c0d;
6186: douta=16'h9c0d;
6187: douta=16'h9c0d;
6188: douta=16'h6aea;
6189: douta=16'h31a8;
6190: douta=16'h2967;
6191: douta=16'h2987;
6192: douta=16'h2106;
6193: douta=16'h39e9;
6194: douta=16'h1926;
6195: douta=16'h1105;
6196: douta=16'h18e5;
6197: douta=16'h18e5;
6198: douta=16'h18e5;
6199: douta=16'h41e8;
6200: douta=16'hacd0;
6201: douta=16'h5aeb;
6202: douta=16'h7c75;
6203: douta=16'h5b90;
6204: douta=16'h52cb;
6205: douta=16'h636f;
6206: douta=16'h634d;
6207: douta=16'h52cc;
6208: douta=16'h73cf;
6209: douta=16'h29a9;
6210: douta=16'h73d0;
6211: douta=16'h4acc;
6212: douta=16'h1106;
6213: douta=16'h426a;
6214: douta=16'h6b6f;
6215: douta=16'h29cb;
6216: douta=16'h6bd0;
6217: douta=16'h6435;
6218: douta=16'h3b10;
6219: douta=16'h19ac;
6220: douta=16'h324d;
6221: douta=16'h42f1;
6222: douta=16'h5b91;
6223: douta=16'h4b51;
6224: douta=16'h4acd;
6225: douta=16'h0800;
6226: douta=16'h1061;
6227: douta=16'h0820;
6228: douta=16'h0000;
6229: douta=16'h4b31;
6230: douta=16'h3a8f;
6231: douta=16'h198a;
6232: douta=16'h53f5;
6233: douta=16'h5c36;
6234: douta=16'h222e;
6235: douta=16'h4a29;
6236: douta=16'hd550;
6237: douta=16'h734b;
6238: douta=16'h5bd5;
6239: douta=16'h5375;
6240: douta=16'h6c78;
6241: douta=16'h84f9;
6242: douta=16'h853a;
6243: douta=16'h8519;
6244: douta=16'h95bb;
6245: douta=16'hae1c;
6246: douta=16'h957a;
6247: douta=16'h7cd9;
6248: douta=16'h853a;
6249: douta=16'h8519;
6250: douta=16'ha5fc;
6251: douta=16'ha5db;
6252: douta=16'h957a;
6253: douta=16'h6c57;
6254: douta=16'h7cb8;
6255: douta=16'h8d5a;
6256: douta=16'h8d5a;
6257: douta=16'h9dbb;
6258: douta=16'h8d5a;
6259: douta=16'h8d39;
6260: douta=16'h7cd9;
6261: douta=16'h6c37;
6262: douta=16'h9dbb;
6263: douta=16'h9ddb;
6264: douta=16'h8539;
6265: douta=16'h7497;
6266: douta=16'h957a;
6267: douta=16'h955a;
6268: douta=16'h7cb8;
6269: douta=16'h7cd8;
6270: douta=16'h95bb;
6271: douta=16'h957b;
6272: douta=16'h74b8;
6273: douta=16'h855a;
6274: douta=16'h7497;
6275: douta=16'h7cb8;
6276: douta=16'h7cf9;
6277: douta=16'h7498;
6278: douta=16'h6c36;
6279: douta=16'h84f9;
6280: douta=16'h84f9;
6281: douta=16'h8d5b;
6282: douta=16'h8d5b;
6283: douta=16'h95bc;
6284: douta=16'h95bc;
6285: douta=16'h8d5b;
6286: douta=16'h8d7b;
6287: douta=16'h959c;
6288: douta=16'h8d9b;
6289: douta=16'h851a;
6290: douta=16'h959b;
6291: douta=16'h95bb;
6292: douta=16'h8d5b;
6293: douta=16'h8d7b;
6294: douta=16'h8d7b;
6295: douta=16'h7cf9;
6296: douta=16'h857b;
6297: douta=16'h853a;
6298: douta=16'h8d5b;
6299: douta=16'h95bd;
6300: douta=16'h853b;
6301: douta=16'h855b;
6302: douta=16'h857b;
6303: douta=16'h74fa;
6304: douta=16'h6458;
6305: douta=16'h751b;
6306: douta=16'h74fa;
6307: douta=16'h6c99;
6308: douta=16'h751b;
6309: douta=16'h7d5b;
6310: douta=16'h8ddc;
6311: douta=16'h6cb9;
6312: douta=16'h7d1a;
6313: douta=16'h74b9;
6314: douta=16'h7d5a;
6315: douta=16'h7d5b;
6316: douta=16'h6cd9;
6317: douta=16'h8d7b;
6318: douta=16'h7d3a;
6319: douta=16'h7d5b;
6320: douta=16'h857b;
6321: douta=16'h7d5b;
6322: douta=16'h74d9;
6323: douta=16'h74fa;
6324: douta=16'h74f9;
6325: douta=16'h2127;
6326: douta=16'h2189;
6327: douta=16'h21ec;
6328: douta=16'h7413;
6329: douta=16'h8cf5;
6330: douta=16'h73f3;
6331: douta=16'h7c55;
6332: douta=16'h63b2;
6333: douta=16'h2a4f;
6334: douta=16'h63d3;
6335: douta=16'h8453;
6336: douta=16'h3b13;
6337: douta=16'h2270;
6338: douta=16'h53d4;
6339: douta=16'h4332;
6340: douta=16'h6416;
6341: douta=16'h6c36;
6342: douta=16'h6c77;
6343: douta=16'h42cf;
6344: douta=16'h6bd4;
6345: douta=16'h7435;
6346: douta=16'h9d17;
6347: douta=16'h8cb5;
6348: douta=16'h4b10;
6349: douta=16'hbe39;
6350: douta=16'h94b4;
6351: douta=16'ha576;
6352: douta=16'hc5d6;
6353: douta=16'heeb8;
6354: douta=16'h8c52;
6355: douta=16'hb596;
6356: douta=16'hb596;
6357: douta=16'h9492;
6358: douta=16'hbd94;
6359: douta=16'h8c10;
6360: douta=16'heeb7;
6361: douta=16'h9cd1;
6362: douta=16'hb574;
6363: douta=16'h83ef;
6364: douta=16'hde96;
6365: douta=16'hb512;
6366: douta=16'heed7;
6367: douta=16'h7b8d;
6368: douta=16'h948f;
6369: douta=16'heef8;
6370: douta=16'hf737;
6371: douta=16'hf718;
6372: douta=16'h734a;
6373: douta=16'h836b;
6374: douta=16'h93cc;
6375: douta=16'h940c;
6376: douta=16'h8bab;
6377: douta=16'h9c0c;
6378: douta=16'hac6d;
6379: douta=16'ha46d;
6380: douta=16'h9c0d;
6381: douta=16'h730b;
6382: douta=16'h41e7;
6383: douta=16'h2946;
6384: douta=16'h1906;
6385: douta=16'h2967;
6386: douta=16'h2968;
6387: douta=16'h1105;
6388: douta=16'h1905;
6389: douta=16'h10e5;
6390: douta=16'h1905;
6391: douta=16'h2125;
6392: douta=16'h840e;
6393: douta=16'h0001;
6394: douta=16'h84d6;
6395: douta=16'h7c33;
6396: douta=16'h8470;
6397: douta=16'h73ef;
6398: douta=16'h29a9;
6399: douta=16'h322a;
6400: douta=16'h3209;
6401: douta=16'h1947;
6402: douta=16'h840f;
6403: douta=16'h73d0;
6404: douta=16'h3a0a;
6405: douta=16'h530d;
6406: douta=16'h4acc;
6407: douta=16'h2148;
6408: douta=16'h5b4e;
6409: douta=16'h7cd6;
6410: douta=16'h3b12;
6411: douta=16'h4b10;
6412: douta=16'h32b0;
6413: douta=16'h21cc;
6414: douta=16'h42cf;
6415: douta=16'h5393;
6416: douta=16'h4b94;
6417: douta=16'h39c8;
6418: douta=16'h1061;
6419: douta=16'h18a2;
6420: douta=16'h10a3;
6421: douta=16'h18e4;
6422: douta=16'h7414;
6423: douta=16'h32af;
6424: douta=16'h3ad1;
6425: douta=16'h5416;
6426: douta=16'h4374;
6427: douta=16'h41a8;
6428: douta=16'h83cb;
6429: douta=16'h3967;
6430: douta=16'h8d7a;
6431: douta=16'h74b8;
6432: douta=16'h3af3;
6433: douta=16'h8d7a;
6434: douta=16'h74b9;
6435: douta=16'h7cf9;
6436: douta=16'h7d19;
6437: douta=16'hae3c;
6438: douta=16'hae3c;
6439: douta=16'h855a;
6440: douta=16'h95bb;
6441: douta=16'h7cd9;
6442: douta=16'h8519;
6443: douta=16'hae1c;
6444: douta=16'ha61c;
6445: douta=16'h7c97;
6446: douta=16'h7c77;
6447: douta=16'h7457;
6448: douta=16'h851a;
6449: douta=16'h8d3a;
6450: douta=16'h9ddc;
6451: douta=16'h851a;
6452: douta=16'h851a;
6453: douta=16'h7cd8;
6454: douta=16'h84f9;
6455: douta=16'h8d39;
6456: douta=16'h959a;
6457: douta=16'h6c36;
6458: douta=16'h7477;
6459: douta=16'h7cb8;
6460: douta=16'h7477;
6461: douta=16'h6c15;
6462: douta=16'h7cb8;
6463: douta=16'h8d7b;
6464: douta=16'h8d5b;
6465: douta=16'h7cd9;
6466: douta=16'h7cb9;
6467: douta=16'h7cd8;
6468: douta=16'h7478;
6469: douta=16'h853a;
6470: douta=16'h7cb8;
6471: douta=16'h7498;
6472: douta=16'h8d5b;
6473: douta=16'h8d5b;
6474: douta=16'h959b;
6475: douta=16'h7cd9;
6476: douta=16'h8d5a;
6477: douta=16'h9ddd;
6478: douta=16'h8d7b;
6479: douta=16'h853a;
6480: douta=16'h8d7b;
6481: douta=16'h95bc;
6482: douta=16'h853a;
6483: douta=16'h855a;
6484: douta=16'h855a;
6485: douta=16'h853a;
6486: douta=16'h855a;
6487: douta=16'h853a;
6488: douta=16'h7d3a;
6489: douta=16'h7d1a;
6490: douta=16'h7cfa;
6491: douta=16'h7d3b;
6492: douta=16'h95bc;
6493: douta=16'h8d5b;
6494: douta=16'h853a;
6495: douta=16'h6c98;
6496: douta=16'h53f6;
6497: douta=16'h6cb9;
6498: douta=16'h7d3b;
6499: douta=16'h6c99;
6500: douta=16'h751b;
6501: douta=16'h74fb;
6502: douta=16'h8d9c;
6503: douta=16'h7d5b;
6504: douta=16'h7d3a;
6505: douta=16'h74b9;
6506: douta=16'h74da;
6507: douta=16'h7d3b;
6508: douta=16'h74fa;
6509: douta=16'h7d1a;
6510: douta=16'h9dfd;
6511: douta=16'h74da;
6512: douta=16'h6cda;
6513: douta=16'h751a;
6514: douta=16'h7d1a;
6515: douta=16'h6c78;
6516: douta=16'h6cb8;
6517: douta=16'h1906;
6518: douta=16'h2168;
6519: douta=16'h3aad;
6520: douta=16'h5b92;
6521: douta=16'h5371;
6522: douta=16'h3a8e;
6523: douta=16'h7c54;
6524: douta=16'hc619;
6525: douta=16'h5373;
6526: douta=16'h4b11;
6527: douta=16'h7c54;
6528: douta=16'h2ad1;
6529: douta=16'h32d2;
6530: douta=16'h32f2;
6531: douta=16'h4311;
6532: douta=16'h7477;
6533: douta=16'h7477;
6534: douta=16'h7cd8;
6535: douta=16'h42f0;
6536: douta=16'h7c96;
6537: douta=16'h7435;
6538: douta=16'ha557;
6539: douta=16'h94d6;
6540: douta=16'h94b5;
6541: douta=16'hbdd8;
6542: douta=16'h8c93;
6543: douta=16'ha535;
6544: douta=16'hcdf6;
6545: douta=16'hc5d6;
6546: douta=16'h94b2;
6547: douta=16'hbdb5;
6548: douta=16'h9cd2;
6549: douta=16'h9470;
6550: douta=16'hcdf5;
6551: douta=16'h52ab;
6552: douta=16'had12;
6553: douta=16'hc5f4;
6554: douta=16'had11;
6555: douta=16'h7bad;
6556: douta=16'hf77a;
6557: douta=16'h630c;
6558: douta=16'hc594;
6559: douta=16'h8c2e;
6560: douta=16'hd614;
6561: douta=16'hbd72;
6562: douta=16'hc613;
6563: douta=16'h838b;
6564: douta=16'h838b;
6565: douta=16'h8b8b;
6566: douta=16'h9bec;
6567: douta=16'h9c0c;
6568: douta=16'ha44c;
6569: douta=16'ha46d;
6570: douta=16'hac8d;
6571: douta=16'hac8d;
6572: douta=16'h836c;
6573: douta=16'h836c;
6574: douta=16'h6b2b;
6575: douta=16'h6aea;
6576: douta=16'h2167;
6577: douta=16'h10c5;
6578: douta=16'h1105;
6579: douta=16'h2125;
6580: douta=16'h10e5;
6581: douta=16'h10e5;
6582: douta=16'h10e5;
6583: douta=16'h10c4;
6584: douta=16'h0021;
6585: douta=16'h0001;
6586: douta=16'h5b2f;
6587: douta=16'h63f3;
6588: douta=16'h6bf2;
6589: douta=16'h4aab;
6590: douta=16'h528a;
6591: douta=16'h10c5;
6592: douta=16'h29a9;
6593: douta=16'h2168;
6594: douta=16'h52cd;
6595: douta=16'h530d;
6596: douta=16'h6b8e;
6597: douta=16'h5b4f;
6598: douta=16'h3a2a;
6599: douta=16'h29a8;
6600: douta=16'h3a4c;
6601: douta=16'h42ef;
6602: douta=16'h324d;
6603: douta=16'h6370;
6604: douta=16'h5372;
6605: douta=16'h324d;
6606: douta=16'h5351;
6607: douta=16'h3ad0;
6608: douta=16'h2a6f;
6609: douta=16'h63f3;
6610: douta=16'h326d;
6611: douta=16'h2989;
6612: douta=16'h2124;
6613: douta=16'h1903;
6614: douta=16'h18e3;
6615: douta=16'h0841;
6616: douta=16'h5b93;
6617: douta=16'h4b31;
6618: douta=16'h4a28;
6619: douta=16'h7b8c;
6620: douta=16'hb63b;
6621: douta=16'h5c16;
6622: douta=16'h8d79;
6623: douta=16'h8d5a;
6624: douta=16'h8d5a;
6625: douta=16'h8519;
6626: douta=16'h7cf9;
6627: douta=16'h74b8;
6628: douta=16'h5bf6;
6629: douta=16'h6c77;
6630: douta=16'h6c57;
6631: douta=16'hae3c;
6632: douta=16'hae1c;
6633: douta=16'h9ddc;
6634: douta=16'h955a;
6635: douta=16'ha5db;
6636: douta=16'h9559;
6637: douta=16'h6c16;
6638: douta=16'h6c56;
6639: douta=16'h8d3a;
6640: douta=16'h8d5a;
6641: douta=16'h9dbb;
6642: douta=16'hae1c;
6643: douta=16'h8d5a;
6644: douta=16'h8539;
6645: douta=16'h8d5a;
6646: douta=16'h8d5a;
6647: douta=16'h8d5a;
6648: douta=16'h8d39;
6649: douta=16'h7cb8;
6650: douta=16'h6c36;
6651: douta=16'h7cb8;
6652: douta=16'h84f8;
6653: douta=16'h6c35;
6654: douta=16'h7456;
6655: douta=16'h9dfc;
6656: douta=16'h95bb;
6657: douta=16'h957a;
6658: douta=16'h8d7a;
6659: douta=16'h7cd9;
6660: douta=16'h7cb9;
6661: douta=16'h7cb8;
6662: douta=16'h7cb9;
6663: douta=16'h853a;
6664: douta=16'h84f9;
6665: douta=16'h7cf9;
6666: douta=16'h7c98;
6667: douta=16'h6416;
6668: douta=16'h957b;
6669: douta=16'h8d9c;
6670: douta=16'h7d1a;
6671: douta=16'h851a;
6672: douta=16'h8d5b;
6673: douta=16'h8d5a;
6674: douta=16'h7d1a;
6675: douta=16'h855b;
6676: douta=16'h853a;
6677: douta=16'h7d1a;
6678: douta=16'h853a;
6679: douta=16'h959b;
6680: douta=16'h853a;
6681: douta=16'h853b;
6682: douta=16'h7d1a;
6683: douta=16'h8d9c;
6684: douta=16'h7cda;
6685: douta=16'h855a;
6686: douta=16'h855a;
6687: douta=16'h8d7b;
6688: douta=16'h855a;
6689: douta=16'h7cf9;
6690: douta=16'h5c37;
6691: douta=16'h74fa;
6692: douta=16'h751a;
6693: douta=16'h74f9;
6694: douta=16'h6cba;
6695: douta=16'h5c38;
6696: douta=16'h6479;
6697: douta=16'h85bc;
6698: douta=16'h74fa;
6699: douta=16'h857c;
6700: douta=16'h7d1b;
6701: douta=16'h6cb9;
6702: douta=16'h7d5b;
6703: douta=16'h7d3b;
6704: douta=16'h855b;
6705: douta=16'h8ddc;
6706: douta=16'h6c78;
6707: douta=16'h74da;
6708: douta=16'h857b;
6709: douta=16'h74b8;
6710: douta=16'h1906;
6711: douta=16'h2988;
6712: douta=16'h4310;
6713: douta=16'h4b31;
6714: douta=16'h8cd6;
6715: douta=16'h7cb8;
6716: douta=16'h5bb4;
6717: douta=16'h3290;
6718: douta=16'h7c33;
6719: douta=16'h7c75;
6720: douta=16'h4b94;
6721: douta=16'h3b32;
6722: douta=16'h4b95;
6723: douta=16'h3290;
6724: douta=16'h3af1;
6725: douta=16'h2a2e;
6726: douta=16'h3ab0;
6727: douta=16'h5351;
6728: douta=16'h7c76;
6729: douta=16'h9539;
6730: douta=16'h7c33;
6731: douta=16'h8cb5;
6732: douta=16'h6c13;
6733: douta=16'h9d15;
6734: douta=16'h9c93;
6735: douta=16'hc5f7;
6736: douta=16'h9c92;
6737: douta=16'h39eb;
6738: douta=16'h6bb0;
6739: douta=16'ha4b1;
6740: douta=16'h9470;
6741: douta=16'hcdf6;
6742: douta=16'ha4f2;
6743: douta=16'h9450;
6744: douta=16'hc5b3;
6745: douta=16'ha4b0;
6746: douta=16'ha4d0;
6747: douta=16'he6b6;
6748: douta=16'hde96;
6749: douta=16'hb572;
6750: douta=16'hce14;
6751: douta=16'hb50f;
6752: douta=16'hce34;
6753: douta=16'heed7;
6754: douta=16'h8bab;
6755: douta=16'h8bac;
6756: douta=16'h8bac;
6757: douta=16'h9c0c;
6758: douta=16'h9c0c;
6759: douta=16'ha40c;
6760: douta=16'hb48d;
6761: douta=16'hb4ad;
6762: douta=16'hac6d;
6763: douta=16'hb48e;
6764: douta=16'hac6d;
6765: douta=16'h93cc;
6766: douta=16'h6aea;
6767: douta=16'h6b0a;
6768: douta=16'h524a;
6769: douta=16'h18e5;
6770: douta=16'h18e5;
6771: douta=16'h10e5;
6772: douta=16'h18e5;
6773: douta=16'h1905;
6774: douta=16'h1905;
6775: douta=16'h1905;
6776: douta=16'h0883;
6777: douta=16'h0000;
6778: douta=16'h3125;
6779: douta=16'h84b6;
6780: douta=16'h7cb6;
6781: douta=16'h29a7;
6782: douta=16'h4229;
6783: douta=16'h10c5;
6784: douta=16'h29a9;
6785: douta=16'h632d;
6786: douta=16'h42ac;
6787: douta=16'h3a6b;
6788: douta=16'h428c;
6789: douta=16'h5b4e;
6790: douta=16'h322b;
6791: douta=16'h6b6f;
6792: douta=16'h322b;
6793: douta=16'h326d;
6794: douta=16'h1927;
6795: douta=16'h21cb;
6796: douta=16'h21ca;
6797: douta=16'h6bd2;
6798: douta=16'h4b31;
6799: douta=16'h4353;
6800: douta=16'h328f;
6801: douta=16'h326e;
6802: douta=16'h320a;
6803: douta=16'h3a4b;
6804: douta=16'h5b50;
6805: douta=16'h31a8;
6806: douta=16'h18c3;
6807: douta=16'h18e3;
6808: douta=16'h0840;
6809: douta=16'h0860;
6810: douta=16'h6a49;
6811: douta=16'h73d2;
6812: douta=16'h9579;
6813: douta=16'h7498;
6814: douta=16'h8d19;
6815: douta=16'h7cd7;
6816: douta=16'h84f9;
6817: douta=16'h7cb8;
6818: douta=16'h8d5a;
6819: douta=16'h8d5a;
6820: douta=16'h5394;
6821: douta=16'h84f9;
6822: douta=16'h7cb8;
6823: douta=16'h5c16;
6824: douta=16'h7cd9;
6825: douta=16'h95bc;
6826: douta=16'h959a;
6827: douta=16'h8519;
6828: douta=16'h84d8;
6829: douta=16'h8d39;
6830: douta=16'h84b8;
6831: douta=16'hadfb;
6832: douta=16'h6cb9;
6833: douta=16'ha5fc;
6834: douta=16'h9ddb;
6835: douta=16'hb65c;
6836: douta=16'h957a;
6837: douta=16'h9dbb;
6838: douta=16'h8519;
6839: douta=16'h84f9;
6840: douta=16'h8d5a;
6841: douta=16'h851a;
6842: douta=16'h8d5a;
6843: douta=16'h8d39;
6844: douta=16'h851a;
6845: douta=16'h8d3a;
6846: douta=16'h8d5a;
6847: douta=16'h7cb8;
6848: douta=16'h7477;
6849: douta=16'h7477;
6850: douta=16'h8d79;
6851: douta=16'h8d5a;
6852: douta=16'h853a;
6853: douta=16'h7456;
6854: douta=16'h6c15;
6855: douta=16'h5bd5;
6856: douta=16'h7cd9;
6857: douta=16'h8d3a;
6858: douta=16'h7cd8;
6859: douta=16'h9ddc;
6860: douta=16'h853a;
6861: douta=16'h6c36;
6862: douta=16'h7cf9;
6863: douta=16'h7cf9;
6864: douta=16'h851a;
6865: douta=16'h853a;
6866: douta=16'h957b;
6867: douta=16'h959c;
6868: douta=16'h853a;
6869: douta=16'h851a;
6870: douta=16'h8d9c;
6871: douta=16'h7d3a;
6872: douta=16'h7d3a;
6873: douta=16'h8d7b;
6874: douta=16'h95dc;
6875: douta=16'h7d1b;
6876: douta=16'h853a;
6877: douta=16'h853a;
6878: douta=16'h7d1a;
6879: douta=16'h8d7b;
6880: douta=16'h855b;
6881: douta=16'h7cfa;
6882: douta=16'h8d9c;
6883: douta=16'h6c37;
6884: douta=16'h53b5;
6885: douta=16'h53b6;
6886: douta=16'h74da;
6887: douta=16'h8dfd;
6888: douta=16'h7d5b;
6889: douta=16'h6cda;
6890: douta=16'h6cba;
6891: douta=16'h859c;
6892: douta=16'h7d5b;
6893: douta=16'h859c;
6894: douta=16'h74fa;
6895: douta=16'h74d9;
6896: douta=16'h8dbc;
6897: douta=16'h857b;
6898: douta=16'h857b;
6899: douta=16'h7d1a;
6900: douta=16'h855b;
6901: douta=16'h6c77;
6902: douta=16'h5b72;
6903: douta=16'h18a4;
6904: douta=16'h8cf6;
6905: douta=16'h8496;
6906: douta=16'h5b72;
6907: douta=16'h42f1;
6908: douta=16'h6c13;
6909: douta=16'h9d37;
6910: douta=16'h8cd6;
6911: douta=16'h5331;
6912: douta=16'h4353;
6913: douta=16'h220e;
6914: douta=16'h6479;
6915: douta=16'h4b73;
6916: douta=16'h6c36;
6917: douta=16'h7497;
6918: douta=16'h5373;
6919: douta=16'h3a6e;
6920: douta=16'h5b72;
6921: douta=16'h5372;
6922: douta=16'h8c74;
6923: douta=16'ha538;
6924: douta=16'hb5b9;
6925: douta=16'h9d35;
6926: douta=16'h3a4d;
6927: douta=16'h7413;
6928: douta=16'hc5f6;
6929: douta=16'hbd55;
6930: douta=16'hbdd6;
6931: douta=16'h8431;
6932: douta=16'h428d;
6933: douta=16'h6b6e;
6934: douta=16'hbd74;
6935: douta=16'hb512;
6936: douta=16'hde76;
6937: douta=16'hbdd3;
6938: douta=16'h842f;
6939: douta=16'h944e;
6940: douta=16'he6d9;
6941: douta=16'hce14;
6942: douta=16'hde96;
6943: douta=16'h942d;
6944: douta=16'had11;
6945: douta=16'had10;
6946: douta=16'h8bab;
6947: douta=16'h8bac;
6948: douta=16'h8bec;
6949: douta=16'ha42c;
6950: douta=16'ha44c;
6951: douta=16'hac6d;
6952: douta=16'hb4ad;
6953: douta=16'hbcce;
6954: douta=16'ha44c;
6955: douta=16'hb48d;
6956: douta=16'hb4ae;
6957: douta=16'h9c0c;
6958: douta=16'h62ca;
6959: douta=16'h62a9;
6960: douta=16'h4a29;
6961: douta=16'h2167;
6962: douta=16'h10e5;
6963: douta=16'h1926;
6964: douta=16'h18e5;
6965: douta=16'h1905;
6966: douta=16'h2106;
6967: douta=16'h1925;
6968: douta=16'h1905;
6969: douta=16'h0000;
6970: douta=16'h0000;
6971: douta=16'h7c95;
6972: douta=16'h63f2;
6973: douta=16'h2187;
6974: douta=16'h630b;
6975: douta=16'h31a7;
6976: douta=16'h18e5;
6977: douta=16'h31a7;
6978: douta=16'h322a;
6979: douta=16'h322a;
6980: douta=16'h6bb0;
6981: douta=16'h2a2b;
6982: douta=16'h2188;
6983: douta=16'h424b;
6984: douta=16'h4a8c;
6985: douta=16'h2a4d;
6986: douta=16'h52ee;
6987: douta=16'h3a8d;
6988: douta=16'h1989;
6989: douta=16'h5351;
6990: douta=16'h4b31;
6991: douta=16'h3aaf;
6992: douta=16'h5b72;
6993: douta=16'h3b11;
6994: douta=16'h3a6d;
6995: douta=16'h428c;
6996: douta=16'h5b50;
6997: douta=16'h6bb2;
6998: douta=16'h10e3;
6999: douta=16'h1082;
7000: douta=16'h1062;
7001: douta=16'h2924;
7002: douta=16'hac2c;
7003: douta=16'hb5da;
7004: douta=16'h84d8;
7005: douta=16'h955a;
7006: douta=16'h84d8;
7007: douta=16'h8d3a;
7008: douta=16'h957a;
7009: douta=16'h7cd8;
7010: douta=16'h6c57;
7011: douta=16'h7457;
7012: douta=16'h6c77;
7013: douta=16'h6415;
7014: douta=16'h84d8;
7015: douta=16'h6c77;
7016: douta=16'h6c36;
7017: douta=16'h84f9;
7018: douta=16'h8d19;
7019: douta=16'h9d9a;
7020: douta=16'h9d9a;
7021: douta=16'h84f8;
7022: douta=16'h63f4;
7023: douta=16'h8d5a;
7024: douta=16'h957b;
7025: douta=16'hb67d;
7026: douta=16'hae3c;
7027: douta=16'ha61c;
7028: douta=16'h8d7a;
7029: douta=16'ha61c;
7030: douta=16'h9dfb;
7031: douta=16'h957b;
7032: douta=16'h8d3a;
7033: douta=16'h8519;
7034: douta=16'h851a;
7035: douta=16'h959a;
7036: douta=16'h7cf9;
7037: douta=16'h8d3a;
7038: douta=16'h8519;
7039: douta=16'h84d9;
7040: douta=16'h8d3a;
7041: douta=16'h8d7a;
7042: douta=16'h7477;
7043: douta=16'h853a;
7044: douta=16'h7cf9;
7045: douta=16'h95bc;
7046: douta=16'h7d19;
7047: douta=16'h7457;
7048: douta=16'h7cd9;
7049: douta=16'h8539;
7050: douta=16'h8519;
7051: douta=16'h74b8;
7052: douta=16'h8d7b;
7053: douta=16'h855a;
7054: douta=16'h7498;
7055: douta=16'h6456;
7056: douta=16'h7477;
7057: douta=16'h95bc;
7058: douta=16'h74b8;
7059: douta=16'h7d1a;
7060: douta=16'h8d7b;
7061: douta=16'h8d7b;
7062: douta=16'h853a;
7063: douta=16'h95bc;
7064: douta=16'h7d1a;
7065: douta=16'h7cd9;
7066: douta=16'h8d5b;
7067: douta=16'h95bc;
7068: douta=16'h8d7b;
7069: douta=16'h74b8;
7070: douta=16'h7d1a;
7071: douta=16'h7d1a;
7072: douta=16'h855b;
7073: douta=16'h851b;
7074: douta=16'h855b;
7075: douta=16'h95dd;
7076: douta=16'h8dbc;
7077: douta=16'h5394;
7078: douta=16'h53f6;
7079: douta=16'h7d7c;
7080: douta=16'h8ddd;
7081: douta=16'h7d7c;
7082: douta=16'h5c78;
7083: douta=16'h859c;
7084: douta=16'h7d3b;
7085: douta=16'h751a;
7086: douta=16'h751a;
7087: douta=16'h74fa;
7088: douta=16'h74d9;
7089: douta=16'h8dbc;
7090: douta=16'h7d5b;
7091: douta=16'h859b;
7092: douta=16'h857b;
7093: douta=16'h7d19;
7094: douta=16'h6416;
7095: douta=16'h31c9;
7096: douta=16'h5351;
7097: douta=16'h9d36;
7098: douta=16'h7c76;
7099: douta=16'h7c55;
7100: douta=16'h326e;
7101: douta=16'h6c14;
7102: douta=16'h8cd6;
7103: douta=16'hadb8;
7104: douta=16'h220d;
7105: douta=16'h2ab0;
7106: douta=16'h224f;
7107: douta=16'h6457;
7108: douta=16'h7436;
7109: douta=16'h7456;
7110: douta=16'h6436;
7111: douta=16'h4b11;
7112: douta=16'h7435;
7113: douta=16'h8496;
7114: douta=16'h9d37;
7115: douta=16'hadba;
7116: douta=16'h9d16;
7117: douta=16'h9493;
7118: douta=16'h4aef;
7119: douta=16'h6370;
7120: douta=16'hbdb5;
7121: douta=16'hcdd6;
7122: douta=16'hb573;
7123: douta=16'h9c91;
7124: douta=16'h9cf2;
7125: douta=16'h7c10;
7126: douta=16'h736d;
7127: douta=16'hbd72;
7128: douta=16'hf737;
7129: douta=16'h9cb0;
7130: douta=16'h840e;
7131: douta=16'h83ee;
7132: douta=16'hde56;
7133: douta=16'hd655;
7134: douta=16'heef8;
7135: douta=16'h8bed;
7136: douta=16'had32;
7137: douta=16'h838b;
7138: douta=16'h93cb;
7139: douta=16'h940c;
7140: douta=16'ha42c;
7141: douta=16'ha42c;
7142: douta=16'hac6c;
7143: douta=16'hb48c;
7144: douta=16'hbcee;
7145: douta=16'hbccd;
7146: douta=16'hc50e;
7147: douta=16'hac4d;
7148: douta=16'h9bec;
7149: douta=16'h8bab;
7150: douta=16'h8b8d;
7151: douta=16'h838b;
7152: douta=16'h5a69;
7153: douta=16'h41e9;
7154: douta=16'h29a8;
7155: douta=16'h2946;
7156: douta=16'h18e5;
7157: douta=16'h2126;
7158: douta=16'h18e5;
7159: douta=16'h18e5;
7160: douta=16'h1104;
7161: douta=16'h10a4;
7162: douta=16'h0022;
7163: douta=16'h2125;
7164: douta=16'h6370;
7165: douta=16'h426c;
7166: douta=16'h3a08;
7167: douta=16'h4269;
7168: douta=16'h10e4;
7169: douta=16'h39a8;
7170: douta=16'h2987;
7171: douta=16'h3a2a;
7172: douta=16'h42ce;
7173: douta=16'h1107;
7174: douta=16'h1968;
7175: douta=16'h4a8b;
7176: douta=16'h1126;
7177: douta=16'h08e6;
7178: douta=16'h4aac;
7179: douta=16'h42ad;
7180: douta=16'h1927;
7181: douta=16'h3a6d;
7182: douta=16'h322b;
7183: douta=16'h6390;
7184: douta=16'h6bd2;
7185: douta=16'h42cf;
7186: douta=16'h2a0c;
7187: douta=16'h3aae;
7188: douta=16'h2a2c;
7189: douta=16'h1128;
7190: douta=16'h6391;
7191: douta=16'h3a4c;
7192: douta=16'h39e8;
7193: douta=16'h6227;
7194: douta=16'h4a29;
7195: douta=16'h7cd7;
7196: douta=16'h7cb7;
7197: douta=16'h7477;
7198: douta=16'h8d5a;
7199: douta=16'h8d39;
7200: douta=16'h6c57;
7201: douta=16'h74b8;
7202: douta=16'h7cd8;
7203: douta=16'h84d8;
7204: douta=16'h7477;
7205: douta=16'h8539;
7206: douta=16'h8d5a;
7207: douta=16'h6c35;
7208: douta=16'h5bd5;
7209: douta=16'h7457;
7210: douta=16'h8d19;
7211: douta=16'h6416;
7212: douta=16'h7c98;
7213: douta=16'h7c96;
7214: douta=16'h9559;
7215: douta=16'h9d7a;
7216: douta=16'h9d9a;
7217: douta=16'hb67d;
7218: douta=16'hae3d;
7219: douta=16'hae3d;
7220: douta=16'h7d1a;
7221: douta=16'h9ddc;
7222: douta=16'hae3d;
7223: douta=16'ha61c;
7224: douta=16'h959b;
7225: douta=16'h95bb;
7226: douta=16'h8519;
7227: douta=16'h7cd8;
7228: douta=16'h8d3a;
7229: douta=16'h853a;
7230: douta=16'h8d5a;
7231: douta=16'h8519;
7232: douta=16'h8d5a;
7233: douta=16'h8d3a;
7234: douta=16'h8519;
7235: douta=16'h8d3a;
7236: douta=16'h957b;
7237: douta=16'h84f9;
7238: douta=16'h7457;
7239: douta=16'h5bf5;
7240: douta=16'h6c56;
7241: douta=16'h853a;
7242: douta=16'h74b8;
7243: douta=16'h851a;
7244: douta=16'h6c37;
7245: douta=16'h74b8;
7246: douta=16'h7498;
7247: douta=16'h7cf9;
7248: douta=16'h851a;
7249: douta=16'h7cd9;
7250: douta=16'h74b8;
7251: douta=16'h6c57;
7252: douta=16'h6c57;
7253: douta=16'h6c77;
7254: douta=16'h7cfa;
7255: douta=16'h8d5a;
7256: douta=16'h8d5a;
7257: douta=16'h7cf9;
7258: douta=16'h855b;
7259: douta=16'h853b;
7260: douta=16'h851a;
7261: douta=16'h855b;
7262: douta=16'h8d9b;
7263: douta=16'h8d7b;
7264: douta=16'h853b;
7265: douta=16'h7d1a;
7266: douta=16'h74b9;
7267: douta=16'h7d3b;
7268: douta=16'h855b;
7269: douta=16'h7d1a;
7270: douta=16'h7d3b;
7271: douta=16'h857c;
7272: douta=16'h7d3a;
7273: douta=16'h6cba;
7274: douta=16'h7d1b;
7275: douta=16'h751a;
7276: douta=16'h6cba;
7277: douta=16'h6cba;
7278: douta=16'h6c99;
7279: douta=16'h7d3b;
7280: douta=16'h8ddc;
7281: douta=16'h74d9;
7282: douta=16'h859c;
7283: douta=16'h8d9b;
7284: douta=16'h8dbc;
7285: douta=16'h74f9;
7286: douta=16'h74d9;
7287: douta=16'h74d8;
7288: douta=16'h4ace;
7289: douta=16'h42cf;
7290: douta=16'hadd9;
7291: douta=16'h8495;
7292: douta=16'h5b92;
7293: douta=16'h7c54;
7294: douta=16'had78;
7295: douta=16'h6371;
7296: douta=16'h2ab0;
7297: douta=16'h32f2;
7298: douta=16'h4312;
7299: douta=16'h5c36;
7300: douta=16'h7c76;
7301: douta=16'h7477;
7302: douta=16'h63f4;
7303: douta=16'h7cb8;
7304: douta=16'h6bf3;
7305: douta=16'h84b7;
7306: douta=16'h7413;
7307: douta=16'h8cb5;
7308: douta=16'h7c13;
7309: douta=16'ha514;
7310: douta=16'hb535;
7311: douta=16'hdeb9;
7312: douta=16'had14;
7313: douta=16'h7b90;
7314: douta=16'h8451;
7315: douta=16'ha4d1;
7316: douta=16'ha4f2;
7317: douta=16'h9cd1;
7318: douta=16'he696;
7319: douta=16'h944f;
7320: douta=16'h9c6f;
7321: douta=16'hce34;
7322: douta=16'hbd92;
7323: douta=16'h7c0d;
7324: douta=16'he6b7;
7325: douta=16'hb531;
7326: douta=16'hbdb2;
7327: douta=16'hb571;
7328: douta=16'h7309;
7329: douta=16'h93ec;
7330: douta=16'h9c0c;
7331: douta=16'h9c0d;
7332: douta=16'hac4d;
7333: douta=16'hb48d;
7334: douta=16'hb4cd;
7335: douta=16'hbced;
7336: douta=16'hcd4f;
7337: douta=16'hd570;
7338: douta=16'hcd4f;
7339: douta=16'hc50f;
7340: douta=16'hac4d;
7341: douta=16'h9c0d;
7342: douta=16'h72ca;
7343: douta=16'h5a68;
7344: douta=16'h62ca;
7345: douta=16'h31c8;
7346: douta=16'h2967;
7347: douta=16'h2146;
7348: douta=16'h630c;
7349: douta=16'h08a4;
7350: douta=16'h18e4;
7351: douta=16'h10e4;
7352: douta=16'h10e4;
7353: douta=16'h1905;
7354: douta=16'h0000;
7355: douta=16'h0000;
7356: douta=16'h0020;
7357: douta=16'h6bf1;
7358: douta=16'h428b;
7359: douta=16'h732b;
7360: douta=16'h940e;
7361: douta=16'h6b4d;
7362: douta=16'h2966;
7363: douta=16'h29a9;
7364: douta=16'h29ea;
7365: douta=16'h422b;
7366: douta=16'h320a;
7367: douta=16'h73ae;
7368: douta=16'h632e;
7369: douta=16'h424b;
7370: douta=16'h42ce;
7371: douta=16'h1968;
7372: douta=16'h1106;
7373: douta=16'h29c9;
7374: douta=16'h4a8c;
7375: douta=16'h4aee;
7376: douta=16'h32ae;
7377: douta=16'h3a4d;
7378: douta=16'h21ca;
7379: douta=16'h3a4c;
7380: douta=16'h322c;
7381: douta=16'h4ad0;
7382: douta=16'h5371;
7383: douta=16'h428d;
7384: douta=16'h49a7;
7385: douta=16'hb48d;
7386: douta=16'h9cb5;
7387: douta=16'h7c97;
7388: douta=16'h84d8;
7389: douta=16'h84d8;
7390: douta=16'h7497;
7391: douta=16'h7477;
7392: douta=16'h7cb7;
7393: douta=16'h84b7;
7394: douta=16'h7477;
7395: douta=16'h8d19;
7396: douta=16'h8519;
7397: douta=16'h8cf8;
7398: douta=16'h8519;
7399: douta=16'h8519;
7400: douta=16'h8d3a;
7401: douta=16'h84d8;
7402: douta=16'h6c57;
7403: douta=16'h7cb7;
7404: douta=16'h8d19;
7405: douta=16'h955a;
7406: douta=16'h84f8;
7407: douta=16'hb61b;
7408: douta=16'h7cd8;
7409: douta=16'h957b;
7410: douta=16'h7498;
7411: douta=16'h9dbc;
7412: douta=16'h7d19;
7413: douta=16'h8d5a;
7414: douta=16'h8d5a;
7415: douta=16'h95db;
7416: douta=16'h959b;
7417: douta=16'h7498;
7418: douta=16'h7cd9;
7419: douta=16'h957b;
7420: douta=16'h9ddc;
7421: douta=16'h8d7a;
7422: douta=16'h7cd9;
7423: douta=16'h8d5a;
7424: douta=16'h8d39;
7425: douta=16'h8d3a;
7426: douta=16'h8d7a;
7427: douta=16'h8d5a;
7428: douta=16'h853a;
7429: douta=16'h6c57;
7430: douta=16'h853a;
7431: douta=16'h851a;
7432: douta=16'h8519;
7433: douta=16'h7477;
7434: douta=16'h6c16;
7435: douta=16'h7498;
7436: douta=16'h8d3a;
7437: douta=16'h853a;
7438: douta=16'h7cd9;
7439: douta=16'h851a;
7440: douta=16'h5bf6;
7441: douta=16'h853a;
7442: douta=16'h74b8;
7443: douta=16'h851a;
7444: douta=16'h7498;
7445: douta=16'h6c77;
7446: douta=16'h6c57;
7447: douta=16'h6437;
7448: douta=16'h6436;
7449: douta=16'h6436;
7450: douta=16'h95bc;
7451: douta=16'h855b;
7452: douta=16'h7cb9;
7453: douta=16'h857b;
7454: douta=16'h7d1a;
7455: douta=16'h7d3a;
7456: douta=16'h95bc;
7457: douta=16'h95dc;
7458: douta=16'h853b;
7459: douta=16'h7d1b;
7460: douta=16'h7cfa;
7461: douta=16'h7d1b;
7462: douta=16'h7d1b;
7463: douta=16'h857c;
7464: douta=16'h7d3a;
7465: douta=16'h74f9;
7466: douta=16'h8d9c;
7467: douta=16'h6c99;
7468: douta=16'h751a;
7469: douta=16'h7d3b;
7470: douta=16'h74fa;
7471: douta=16'h7d5b;
7472: douta=16'h7d5a;
7473: douta=16'h7d5a;
7474: douta=16'h6cb8;
7475: douta=16'h7cf9;
7476: douta=16'h7d5b;
7477: douta=16'h855b;
7478: douta=16'h7d3a;
7479: douta=16'h7cf9;
7480: douta=16'h1928;
7481: douta=16'hb5d9;
7482: douta=16'h2a0c;
7483: douta=16'h5b71;
7484: douta=16'h8474;
7485: douta=16'h7c33;
7486: douta=16'h3a4c;
7487: douta=16'h73b0;
7488: douta=16'h2a6f;
7489: douta=16'h19ee;
7490: douta=16'h32f1;
7491: douta=16'h4b74;
7492: douta=16'h7c96;
7493: douta=16'h7cb8;
7494: douta=16'h6c16;
7495: douta=16'h5bb3;
7496: douta=16'h5310;
7497: douta=16'h6c14;
7498: douta=16'h8433;
7499: douta=16'h9d16;
7500: douta=16'h9cd6;
7501: douta=16'ha4f3;
7502: douta=16'had75;
7503: douta=16'hb555;
7504: douta=16'hbd75;
7505: douta=16'had33;
7506: douta=16'hce35;
7507: douta=16'had13;
7508: douta=16'h8c70;
7509: douta=16'h8c50;
7510: douta=16'h8c30;
7511: douta=16'ha4b0;
7512: douta=16'hc5d4;
7513: douta=16'hde56;
7514: douta=16'had11;
7515: douta=16'h9c8f;
7516: douta=16'hd655;
7517: douta=16'hd635;
7518: douta=16'hd676;
7519: douta=16'h732a;
7520: douta=16'h7b4b;
7521: douta=16'h9bec;
7522: douta=16'ha44d;
7523: douta=16'h9c0c;
7524: douta=16'ha44c;
7525: douta=16'hbcce;
7526: douta=16'hbcee;
7527: douta=16'hc50e;
7528: douta=16'hd590;
7529: douta=16'hd590;
7530: douta=16'hcd70;
7531: douta=16'hd591;
7532: douta=16'hbcee;
7533: douta=16'hac6d;
7534: douta=16'h93ed;
7535: douta=16'h6aa9;
7536: douta=16'h5a69;
7537: douta=16'h526b;
7538: douta=16'h39c8;
7539: douta=16'h2987;
7540: douta=16'h5aaa;
7541: douta=16'h2125;
7542: douta=16'h10a4;
7543: douta=16'h10e4;
7544: douta=16'h18e5;
7545: douta=16'h18e5;
7546: douta=16'h0000;
7547: douta=16'h0001;
7548: douta=16'h0000;
7549: douta=16'h7412;
7550: douta=16'h4a8c;
7551: douta=16'h52a9;
7552: douta=16'h5aaa;
7553: douta=16'h8c2e;
7554: douta=16'h734d;
7555: douta=16'h4a8b;
7556: douta=16'h3a4c;
7557: douta=16'h424b;
7558: douta=16'h31ea;
7559: douta=16'h320a;
7560: douta=16'h73cf;
7561: douta=16'h6b4e;
7562: douta=16'h73b0;
7563: douta=16'h3a2b;
7564: douta=16'h29ca;
7565: douta=16'h1148;
7566: douta=16'h2168;
7567: douta=16'h532f;
7568: douta=16'h21aa;
7569: douta=16'h3a2b;
7570: douta=16'h326d;
7571: douta=16'h19aa;
7572: douta=16'h1969;
7573: douta=16'h0908;
7574: douta=16'h4b2f;
7575: douta=16'h630d;
7576: douta=16'h9b8d;
7577: douta=16'h9c0c;
7578: douta=16'hb63c;
7579: douta=16'ha5db;
7580: douta=16'h8d39;
7581: douta=16'h7cb8;
7582: douta=16'h959a;
7583: douta=16'h9559;
7584: douta=16'h6c37;
7585: douta=16'h7497;
7586: douta=16'h84d8;
7587: douta=16'h7c97;
7588: douta=16'h9dba;
7589: douta=16'h7cb8;
7590: douta=16'h7cf8;
7591: douta=16'h957a;
7592: douta=16'h955a;
7593: douta=16'h8d3a;
7594: douta=16'h6c57;
7595: douta=16'h7456;
7596: douta=16'h7497;
7597: douta=16'h84f9;
7598: douta=16'h8d19;
7599: douta=16'hbe7c;
7600: douta=16'h84f9;
7601: douta=16'h9dbb;
7602: douta=16'h9d9a;
7603: douta=16'h959a;
7604: douta=16'h8d7b;
7605: douta=16'h7cb8;
7606: douta=16'h853a;
7607: douta=16'h851a;
7608: douta=16'h855a;
7609: douta=16'h7d19;
7610: douta=16'h6c57;
7611: douta=16'h6c98;
7612: douta=16'h8d7b;
7613: douta=16'h959b;
7614: douta=16'h8539;
7615: douta=16'h84f9;
7616: douta=16'h84f9;
7617: douta=16'h7cd8;
7618: douta=16'h853a;
7619: douta=16'h8d7b;
7620: douta=16'h959b;
7621: douta=16'h63f5;
7622: douta=16'h5b94;
7623: douta=16'h7cb8;
7624: douta=16'h7477;
7625: douta=16'h84f9;
7626: douta=16'h84f9;
7627: douta=16'h6457;
7628: douta=16'h7cf9;
7629: douta=16'h7cf9;
7630: douta=16'h7498;
7631: douta=16'h7cd9;
7632: douta=16'h853a;
7633: douta=16'h6c57;
7634: douta=16'h7cd9;
7635: douta=16'h7cd9;
7636: douta=16'h7cfa;
7637: douta=16'h7d1a;
7638: douta=16'h6436;
7639: douta=16'h7498;
7640: douta=16'h6c57;
7641: douta=16'h6416;
7642: douta=16'h7498;
7643: douta=16'h857b;
7644: douta=16'h8d9b;
7645: douta=16'h7cd9;
7646: douta=16'h7cfa;
7647: douta=16'h7d3a;
7648: douta=16'h7d3a;
7649: douta=16'h8d9c;
7650: douta=16'h95dd;
7651: douta=16'h857c;
7652: douta=16'h7cfa;
7653: douta=16'h7d1a;
7654: douta=16'h7d3b;
7655: douta=16'h855b;
7656: douta=16'h8dbc;
7657: douta=16'h74fa;
7658: douta=16'h857b;
7659: douta=16'h857c;
7660: douta=16'h6458;
7661: douta=16'h6478;
7662: douta=16'h7d3b;
7663: douta=16'h6cd9;
7664: douta=16'h8dbc;
7665: douta=16'h857b;
7666: douta=16'h857b;
7667: douta=16'h7d1b;
7668: douta=16'h74d9;
7669: douta=16'h7d3b;
7670: douta=16'h7d3a;
7671: douta=16'h74d9;
7672: douta=16'h08a4;
7673: douta=16'h7c54;
7674: douta=16'h9cf6;
7675: douta=16'h8cd6;
7676: douta=16'h6bd3;
7677: douta=16'h6bd3;
7678: douta=16'h8433;
7679: douta=16'ha4f4;
7680: douta=16'h3312;
7681: douta=16'h4b95;
7682: douta=16'h220d;
7683: douta=16'h4b73;
7684: douta=16'h5bb3;
7685: douta=16'h7477;
7686: douta=16'h63f4;
7687: douta=16'h428f;
7688: douta=16'h5310;
7689: douta=16'h42af;
7690: douta=16'h6392;
7691: douta=16'h6bb2;
7692: douta=16'ha557;
7693: douta=16'hbd96;
7694: douta=16'hb556;
7695: douta=16'hbdb6;
7696: douta=16'h9450;
7697: douta=16'hacf2;
7698: douta=16'hbdb4;
7699: douta=16'ha4f2;
7700: douta=16'hb533;
7701: douta=16'h8c2f;
7702: douta=16'h9c91;
7703: douta=16'hb532;
7704: douta=16'hbd73;
7705: douta=16'he6b7;
7706: douta=16'hcdf4;
7707: douta=16'h9cb0;
7708: douta=16'hbdb3;
7709: douta=16'he6b6;
7710: douta=16'hb592;
7711: douta=16'h7b4a;
7712: douta=16'h93cb;
7713: douta=16'h93cb;
7714: douta=16'hac6c;
7715: douta=16'hac8d;
7716: douta=16'hb4ad;
7717: douta=16'hcd6f;
7718: douta=16'hd5b1;
7719: douta=16'hd591;
7720: douta=16'hddf2;
7721: douta=16'hddd2;
7722: douta=16'hddf2;
7723: douta=16'hddd1;
7724: douta=16'he613;
7725: douta=16'he654;
7726: douta=16'hc50f;
7727: douta=16'h8c0f;
7728: douta=16'h4a08;
7729: douta=16'h7bce;
7730: douta=16'h4a6b;
7731: douta=16'h31a8;
7732: douta=16'h4a4a;
7733: douta=16'h2166;
7734: douta=16'h2126;
7735: douta=16'h2125;
7736: douta=16'h1905;
7737: douta=16'h10e4;
7738: douta=16'h2125;
7739: douta=16'h0000;
7740: douta=16'h0000;
7741: douta=16'h0062;
7742: douta=16'h5b2f;
7743: douta=16'h29c9;
7744: douta=16'h2126;
7745: douta=16'h83cd;
7746: douta=16'h5269;
7747: douta=16'h632c;
7748: douta=16'h2146;
7749: douta=16'h31c9;
7750: douta=16'h21a8;
7751: douta=16'h2147;
7752: douta=16'h324a;
7753: douta=16'h73b0;
7754: douta=16'h4aad;
7755: douta=16'h322c;
7756: douta=16'h324c;
7757: douta=16'h1968;
7758: douta=16'h29a9;
7759: douta=16'h2189;
7760: douta=16'h3a09;
7761: douta=16'h320b;
7762: douta=16'h1969;
7763: douta=16'h2189;
7764: douta=16'h29ec;
7765: douta=16'h0908;
7766: douta=16'h198a;
7767: douta=16'h322c;
7768: douta=16'h8bab;
7769: douta=16'h52cd;
7770: douta=16'h957a;
7771: douta=16'h7497;
7772: douta=16'h84d8;
7773: douta=16'h8d19;
7774: douta=16'h7cb8;
7775: douta=16'h959b;
7776: douta=16'h6c36;
7777: douta=16'h84f9;
7778: douta=16'h957a;
7779: douta=16'h8518;
7780: douta=16'h7457;
7781: douta=16'h84f9;
7782: douta=16'h84f9;
7783: douta=16'h853a;
7784: douta=16'h7497;
7785: douta=16'h84f9;
7786: douta=16'h8d79;
7787: douta=16'h7cd8;
7788: douta=16'h7cb8;
7789: douta=16'h8519;
7790: douta=16'h9d9b;
7791: douta=16'h9ddc;
7792: douta=16'h7cd9;
7793: douta=16'h8d7a;
7794: douta=16'h8519;
7795: douta=16'h9ddb;
7796: douta=16'h8519;
7797: douta=16'h84f8;
7798: douta=16'h8539;
7799: douta=16'h959b;
7800: douta=16'h7498;
7801: douta=16'h6437;
7802: douta=16'h6c77;
7803: douta=16'h5c37;
7804: douta=16'h959b;
7805: douta=16'h8d5a;
7806: douta=16'h74b8;
7807: douta=16'h5bd5;
7808: douta=16'h6416;
7809: douta=16'h9dbb;
7810: douta=16'h84f9;
7811: douta=16'h8d5b;
7812: douta=16'h855a;
7813: douta=16'h7cd9;
7814: douta=16'h7cd9;
7815: douta=16'h8d7b;
7816: douta=16'h74b8;
7817: douta=16'h5bd4;
7818: douta=16'h6c36;
7819: douta=16'h7cf9;
7820: douta=16'h5bb4;
7821: douta=16'h7cd9;
7822: douta=16'h6c57;
7823: douta=16'h5bb4;
7824: douta=16'h7cf9;
7825: douta=16'h855b;
7826: douta=16'h7477;
7827: douta=16'h7457;
7828: douta=16'h5bd4;
7829: douta=16'h6c97;
7830: douta=16'h6415;
7831: douta=16'h6415;
7832: douta=16'h7498;
7833: douta=16'h74b8;
7834: douta=16'h6416;
7835: douta=16'h7cd9;
7836: douta=16'h74f9;
7837: douta=16'h7d1a;
7838: douta=16'h7cfa;
7839: douta=16'h855b;
7840: douta=16'h857b;
7841: douta=16'h853c;
7842: douta=16'h7d1a;
7843: douta=16'h74da;
7844: douta=16'h7cfb;
7845: douta=16'h8dbd;
7846: douta=16'h8d7c;
7847: douta=16'h74b9;
7848: douta=16'h7cfa;
7849: douta=16'h6cb9;
7850: douta=16'h74fa;
7851: douta=16'h7d3a;
7852: douta=16'h7cfa;
7853: douta=16'h7d1a;
7854: douta=16'h7d3a;
7855: douta=16'h74fa;
7856: douta=16'h6458;
7857: douta=16'h5c37;
7858: douta=16'h857b;
7859: douta=16'h857b;
7860: douta=16'h855b;
7861: douta=16'h8dbc;
7862: douta=16'h751a;
7863: douta=16'h74d9;
7864: douta=16'h3a4c;
7865: douta=16'h7474;
7866: douta=16'h8cb5;
7867: douta=16'h4b0f;
7868: douta=16'h42ae;
7869: douta=16'h6391;
7870: douta=16'h9d15;
7871: douta=16'h3a8d;
7872: douta=16'h222f;
7873: douta=16'h32d1;
7874: douta=16'h2a2e;
7875: douta=16'h4333;
7876: douta=16'h5393;
7877: douta=16'h84b8;
7878: douta=16'h4b10;
7879: douta=16'h42af;
7880: douta=16'h7c75;
7881: douta=16'h7454;
7882: douta=16'h94d6;
7883: douta=16'h9d16;
7884: douta=16'h8c95;
7885: douta=16'h5b2f;
7886: douta=16'h7bf1;
7887: douta=16'h9cf3;
7888: douta=16'hcdd6;
7889: douta=16'hc5f5;
7890: douta=16'h9cd2;
7891: douta=16'h62cb;
7892: douta=16'h8bee;
7893: douta=16'h83ee;
7894: douta=16'hce36;
7895: douta=16'heef8;
7896: douta=16'hd677;
7897: douta=16'hbd92;
7898: douta=16'hb531;
7899: douta=16'hbdb3;
7900: douta=16'hff7a;
7901: douta=16'h6ae9;
7902: douta=16'h7b0a;
7903: douta=16'h8b8b;
7904: douta=16'h93eb;
7905: douta=16'h9bec;
7906: douta=16'hac6c;
7907: douta=16'hb48d;
7908: douta=16'hbccd;
7909: douta=16'hcd70;
7910: douta=16'hddf3;
7911: douta=16'he613;
7912: douta=16'hde13;
7913: douta=16'he634;
7914: douta=16'hddf3;
7915: douta=16'he633;
7916: douta=16'hcd6f;
7917: douta=16'hcd90;
7918: douta=16'hb4f0;
7919: douta=16'h3165;
7920: douta=16'ha46f;
7921: douta=16'h62eb;
7922: douta=16'h39e9;
7923: douta=16'h4209;
7924: douta=16'h39e9;
7925: douta=16'h29a8;
7926: douta=16'h29a8;
7927: douta=16'h2946;
7928: douta=16'h10a3;
7929: douta=16'h1905;
7930: douta=16'h18e4;
7931: douta=16'h2145;
7932: douta=16'h0883;
7933: douta=16'h0022;
7934: douta=16'h1106;
7935: douta=16'h1968;
7936: douta=16'h1926;
7937: douta=16'h10e5;
7938: douta=16'h08c4;
7939: douta=16'h4a48;
7940: douta=16'h4208;
7941: douta=16'h2966;
7942: douta=16'h8c0e;
7943: douta=16'h630d;
7944: douta=16'h324d;
7945: douta=16'h21cb;
7946: douta=16'h1948;
7947: douta=16'h29a9;
7948: douta=16'h320a;
7949: douta=16'h4aab;
7950: douta=16'h29ca;
7951: douta=16'h29a9;
7952: douta=16'h3a09;
7953: douta=16'h29a8;
7954: douta=16'h4acc;
7955: douta=16'h29ca;
7956: douta=16'h322a;
7957: douta=16'h8452;
7958: douta=16'h530f;
7959: douta=16'h32af;
7960: douta=16'h5aed;
7961: douta=16'ha598;
7962: douta=16'h959b;
7963: douta=16'h8519;
7964: douta=16'h9dbb;
7965: douta=16'h8d38;
7966: douta=16'h8d5a;
7967: douta=16'h8519;
7968: douta=16'haddc;
7969: douta=16'h7477;
7970: douta=16'h7cd8;
7971: douta=16'h84f9;
7972: douta=16'h8d19;
7973: douta=16'ha5dc;
7974: douta=16'h5bb4;
7975: douta=16'h8519;
7976: douta=16'h9dbb;
7977: douta=16'h8539;
7978: douta=16'h84d9;
7979: douta=16'h9559;
7980: douta=16'h8d7a;
7981: douta=16'h959b;
7982: douta=16'h8d3a;
7983: douta=16'h957a;
7984: douta=16'ha5db;
7985: douta=16'h853a;
7986: douta=16'h8519;
7987: douta=16'h8d3a;
7988: douta=16'h959a;
7989: douta=16'h84d8;
7990: douta=16'h84f9;
7991: douta=16'h7cd9;
7992: douta=16'h853a;
7993: douta=16'h957a;
7994: douta=16'h6417;
7995: douta=16'h74b8;
7996: douta=16'h74b8;
7997: douta=16'h959b;
7998: douta=16'h9d9c;
7999: douta=16'h7cd8;
8000: douta=16'h955a;
8001: douta=16'h5bd5;
8002: douta=16'h5c16;
8003: douta=16'h853a;
8004: douta=16'h7d3a;
8005: douta=16'h7d1a;
8006: douta=16'h7d3b;
8007: douta=16'h7498;
8008: douta=16'h74d9;
8009: douta=16'h7d1a;
8010: douta=16'h7cf9;
8011: douta=16'h5bf5;
8012: douta=16'h6c57;
8013: douta=16'h8d39;
8014: douta=16'h6c56;
8015: douta=16'h6c77;
8016: douta=16'h7cd9;
8017: douta=16'h5b94;
8018: douta=16'h6436;
8019: douta=16'h6cb8;
8020: douta=16'h7456;
8021: douta=16'h6c15;
8022: douta=16'h63f5;
8023: douta=16'h6c77;
8024: douta=16'h6415;
8025: douta=16'h63f4;
8026: douta=16'h5bd5;
8027: douta=16'h6c78;
8028: douta=16'h6c98;
8029: douta=16'h74d9;
8030: douta=16'h6c78;
8031: douta=16'h6c78;
8032: douta=16'h855b;
8033: douta=16'h855c;
8034: douta=16'h857c;
8035: douta=16'h855c;
8036: douta=16'h859c;
8037: douta=16'h7cfa;
8038: douta=16'h855b;
8039: douta=16'h7cfa;
8040: douta=16'h7d3b;
8041: douta=16'h855b;
8042: douta=16'h857b;
8043: douta=16'h6c98;
8044: douta=16'h7d1a;
8045: douta=16'h7d1a;
8046: douta=16'h8d9c;
8047: douta=16'h6478;
8048: douta=16'h857c;
8049: douta=16'h8dbc;
8050: douta=16'h6458;
8051: douta=16'h7d3a;
8052: douta=16'h7d5b;
8053: douta=16'h74d9;
8054: douta=16'h8dbc;
8055: douta=16'h857c;
8056: douta=16'h5b73;
8057: douta=16'h52cd;
8058: douta=16'h5350;
8059: douta=16'h8cb5;
8060: douta=16'h63b2;
8061: douta=16'h8c73;
8062: douta=16'h21aa;
8063: douta=16'h73d2;
8064: douta=16'h3b33;
8065: douta=16'h4bd6;
8066: douta=16'h198b;
8067: douta=16'h3b12;
8068: douta=16'h42d0;
8069: douta=16'h5352;
8070: douta=16'h6c35;
8071: douta=16'h6bf4;
8072: douta=16'h5b51;
8073: douta=16'h6bf3;
8074: douta=16'h7413;
8075: douta=16'h9d17;
8076: douta=16'h9d36;
8077: douta=16'h9493;
8078: douta=16'h7c11;
8079: douta=16'h73b0;
8080: douta=16'h9c71;
8081: douta=16'hb574;
8082: douta=16'he677;
8083: douta=16'hb553;
8084: douta=16'ha4d1;
8085: douta=16'h730c;
8086: douta=16'h8c30;
8087: douta=16'had12;
8088: douta=16'he696;
8089: douta=16'heef8;
8090: douta=16'hc5d3;
8091: douta=16'h8c4f;
8092: douta=16'hce14;
8093: douta=16'h6ac9;
8094: douta=16'h732a;
8095: douta=16'h93ab;
8096: douta=16'h93eb;
8097: douta=16'h9c0c;
8098: douta=16'hb48d;
8099: douta=16'hbccd;
8100: douta=16'hbced;
8101: douta=16'hd5b1;
8102: douta=16'hddf2;
8103: douta=16'hde33;
8104: douta=16'hddf2;
8105: douta=16'hddf3;
8106: douta=16'he613;
8107: douta=16'hde12;
8108: douta=16'hc56f;
8109: douta=16'hc50f;
8110: douta=16'hc531;
8111: douta=16'h6aa9;
8112: douta=16'h9c2e;
8113: douta=16'h5acb;
8114: douta=16'h29a9;
8115: douta=16'h62cb;
8116: douta=16'h4229;
8117: douta=16'h31a8;
8118: douta=16'h2967;
8119: douta=16'h4229;
8120: douta=16'h2966;
8121: douta=16'h1904;
8122: douta=16'h10e4;
8123: douta=16'h18c4;
8124: douta=16'h1905;
8125: douta=16'h0001;
8126: douta=16'h10a5;
8127: douta=16'h2a0b;
8128: douta=16'h10e5;
8129: douta=16'h10e5;
8130: douta=16'h1946;
8131: douta=16'h630a;
8132: douta=16'h62ea;
8133: douta=16'h41e7;
8134: douta=16'h4249;
8135: douta=16'h6b2b;
8136: douta=16'h320b;
8137: douta=16'h4aee;
8138: douta=16'h29ea;
8139: douta=16'h3a2b;
8140: douta=16'h1148;
8141: douta=16'h1127;
8142: douta=16'h0084;
8143: douta=16'h426b;
8144: douta=16'h52ac;
8145: douta=16'h29a9;
8146: douta=16'h29ea;
8147: douta=16'h3a2c;
8148: douta=16'h1148;
8149: douta=16'h29ea;
8150: douta=16'h31a9;
8151: douta=16'h21cb;
8152: douta=16'h5b0d;
8153: douta=16'h9dba;
8154: douta=16'h6c77;
8155: douta=16'h84f9;
8156: douta=16'h9d9a;
8157: douta=16'h9d9a;
8158: douta=16'h7cd8;
8159: douta=16'h8d19;
8160: douta=16'ha5bb;
8161: douta=16'h957a;
8162: douta=16'h8d19;
8163: douta=16'h7477;
8164: douta=16'h8519;
8165: douta=16'h7477;
8166: douta=16'h959b;
8167: douta=16'h6c36;
8168: douta=16'h6c36;
8169: douta=16'h7498;
8170: douta=16'h84d8;
8171: douta=16'h8519;
8172: douta=16'h8d39;
8173: douta=16'h8d39;
8174: douta=16'h8d39;
8175: douta=16'ha5fb;
8176: douta=16'h957a;
8177: douta=16'h6c77;
8178: douta=16'h8d59;
8179: douta=16'h959a;
8180: douta=16'h8d19;
8181: douta=16'h9d9a;
8182: douta=16'h7cd8;
8183: douta=16'h7477;
8184: douta=16'h7cf9;
8185: douta=16'ha5fc;
8186: douta=16'h8d59;
8187: douta=16'h6c56;
8188: douta=16'h6416;
8189: douta=16'h6c77;
8190: douta=16'h7cb8;
8191: douta=16'h8d39;
8192: douta=16'h8d3a;
8193: douta=16'h853a;
8194: douta=16'h5394;
8195: douta=16'h6cda;
8196: douta=16'h6cb9;
8197: douta=16'h6457;
8198: douta=16'h6c98;
8199: douta=16'h7d3a;
8200: douta=16'h74b8;
8201: douta=16'h74b8;
8202: douta=16'h6c77;
8203: douta=16'h7cb8;
8204: douta=16'h6c15;
8205: douta=16'h7477;
8206: douta=16'h84d8;
8207: douta=16'h7476;
8208: douta=16'h6c14;
8209: douta=16'h84d9;
8210: douta=16'h5b73;
8211: douta=16'h5b73;
8212: douta=16'h7cf8;
8213: douta=16'h7cb8;
8214: douta=16'h4b31;
8215: douta=16'h7cb8;
8216: douta=16'h6c56;
8217: douta=16'h7497;
8218: douta=16'h5bf5;
8219: douta=16'h4b94;
8220: douta=16'h6417;
8221: douta=16'h855b;
8222: douta=16'h7d1a;
8223: douta=16'h74fa;
8224: douta=16'h857c;
8225: douta=16'h7d3b;
8226: douta=16'h7cfb;
8227: douta=16'h7d3b;
8228: douta=16'h751b;
8229: douta=16'h7d1b;
8230: douta=16'h7cfa;
8231: douta=16'h7d1a;
8232: douta=16'h6c98;
8233: douta=16'h7d3a;
8234: douta=16'h857b;
8235: douta=16'h7cfa;
8236: douta=16'h74b9;
8237: douta=16'h7cfa;
8238: douta=16'h74d9;
8239: douta=16'h855b;
8240: douta=16'h74d9;
8241: douta=16'h7d1a;
8242: douta=16'h6437;
8243: douta=16'h7499;
8244: douta=16'h855b;
8245: douta=16'h855b;
8246: douta=16'h7d5b;
8247: douta=16'h7d3b;
8248: douta=16'h6c77;
8249: douta=16'h532f;
8250: douta=16'h7412;
8251: douta=16'h5330;
8252: douta=16'h6bd2;
8253: douta=16'h9493;
8254: douta=16'h6391;
8255: douta=16'h7c53;
8256: douta=16'h32b1;
8257: douta=16'h4b94;
8258: douta=16'h3b12;
8259: douta=16'h4b95;
8260: douta=16'h3ab0;
8261: douta=16'h5b73;
8262: douta=16'h63d4;
8263: douta=16'h6c35;
8264: douta=16'h73f4;
8265: douta=16'h7c76;
8266: douta=16'h424b;
8267: douta=16'h6350;
8268: douta=16'h73f1;
8269: douta=16'h9cb4;
8270: douta=16'h9cd4;
8271: douta=16'hbd96;
8272: douta=16'h8410;
8273: douta=16'ha4b1;
8274: douta=16'hd615;
8275: douta=16'hb532;
8276: douta=16'hcdf5;
8277: douta=16'hb511;
8278: douta=16'h6b2c;
8279: douta=16'had10;
8280: douta=16'hd5f5;
8281: douta=16'hde76;
8282: douta=16'hbdd4;
8283: douta=16'ha4d0;
8284: douta=16'h732a;
8285: douta=16'h7b2a;
8286: douta=16'h8b8b;
8287: douta=16'h8b6a;
8288: douta=16'hb48c;
8289: douta=16'hac6c;
8290: douta=16'hbccd;
8291: douta=16'hc50e;
8292: douta=16'hd5d2;
8293: douta=16'hde33;
8294: douta=16'he654;
8295: douta=16'he634;
8296: douta=16'hddf2;
8297: douta=16'hd5b1;
8298: douta=16'hddd1;
8299: douta=16'hcd71;
8300: douta=16'hc50f;
8301: douta=16'hac8f;
8302: douta=16'hac6e;
8303: douta=16'hb4cf;
8304: douta=16'h9c4d;
8305: douta=16'h5acb;
8306: douta=16'h4a4a;
8307: douta=16'h8bed;
8308: douta=16'h62eb;
8309: douta=16'h424b;
8310: douta=16'h31ea;
8311: douta=16'h29c8;
8312: douta=16'h1947;
8313: douta=16'h31c8;
8314: douta=16'h10a4;
8315: douta=16'h18c4;
8316: douta=16'h10e4;
8317: douta=16'h10e4;
8318: douta=16'h0000;
8319: douta=16'h0042;
8320: douta=16'h29ca;
8321: douta=16'h2168;
8322: douta=16'h10e5;
8323: douta=16'h1906;
8324: douta=16'h5a89;
8325: douta=16'h2125;
8326: douta=16'h39e7;
8327: douta=16'h6b2b;
8328: douta=16'h4a28;
8329: douta=16'h7bef;
8330: douta=16'h1969;
8331: douta=16'h29c9;
8332: douta=16'h00c7;
8333: douta=16'h1127;
8334: douta=16'h1127;
8335: douta=16'h4a6a;
8336: douta=16'h29c9;
8337: douta=16'h73af;
8338: douta=16'h428b;
8339: douta=16'h29eb;
8340: douta=16'h424b;
8341: douta=16'h29c9;
8342: douta=16'h1906;
8343: douta=16'h3146;
8344: douta=16'h8475;
8345: douta=16'h8d7a;
8346: douta=16'h8518;
8347: douta=16'h8d59;
8348: douta=16'h8d59;
8349: douta=16'h7cd8;
8350: douta=16'h3ab0;
8351: douta=16'h4b53;
8352: douta=16'h8519;
8353: douta=16'h7456;
8354: douta=16'h9d9b;
8355: douta=16'ha5db;
8356: douta=16'h7498;
8357: douta=16'h84f9;
8358: douta=16'ha5db;
8359: douta=16'h7cb8;
8360: douta=16'h957a;
8361: douta=16'h7cd8;
8362: douta=16'h8d7a;
8363: douta=16'h84f9;
8364: douta=16'h8d5a;
8365: douta=16'h8d7a;
8366: douta=16'h7cd9;
8367: douta=16'h9d9a;
8368: douta=16'h8d5a;
8369: douta=16'h8519;
8370: douta=16'h8539;
8371: douta=16'h9ddc;
8372: douta=16'ha5db;
8373: douta=16'h84f9;
8374: douta=16'h63d5;
8375: douta=16'h7c98;
8376: douta=16'h8d7a;
8377: douta=16'h7cd7;
8378: douta=16'h84f8;
8379: douta=16'h84b8;
8380: douta=16'h7497;
8381: douta=16'h6415;
8382: douta=16'h7cb8;
8383: douta=16'h3af1;
8384: douta=16'h4b53;
8385: douta=16'h7d3b;
8386: douta=16'h751b;
8387: douta=16'h74d9;
8388: douta=16'h6457;
8389: douta=16'h5bd5;
8390: douta=16'h6416;
8391: douta=16'h3ab0;
8392: douta=16'h7c98;
8393: douta=16'h74b8;
8394: douta=16'h6c56;
8395: douta=16'h7497;
8396: douta=16'h7477;
8397: douta=16'h6c36;
8398: douta=16'h7476;
8399: douta=16'h7c97;
8400: douta=16'h63f4;
8401: douta=16'h6c14;
8402: douta=16'h63f4;
8403: douta=16'h7476;
8404: douta=16'h7477;
8405: douta=16'h7476;
8406: douta=16'h6c57;
8407: douta=16'h63f5;
8408: douta=16'h6c35;
8409: douta=16'h5bd4;
8410: douta=16'h5bd4;
8411: douta=16'h7d1b;
8412: douta=16'h6c99;
8413: douta=16'h53f6;
8414: douta=16'h6499;
8415: douta=16'h4b94;
8416: douta=16'h74fa;
8417: douta=16'h855b;
8418: douta=16'h855b;
8419: douta=16'h8d9c;
8420: douta=16'h7d5b;
8421: douta=16'h7d1a;
8422: douta=16'h6c98;
8423: douta=16'h853b;
8424: douta=16'h7d1a;
8425: douta=16'h857c;
8426: douta=16'h7d5b;
8427: douta=16'h7d1a;
8428: douta=16'h8d7b;
8429: douta=16'h855b;
8430: douta=16'h857b;
8431: douta=16'h8dbc;
8432: douta=16'h855b;
8433: douta=16'h857b;
8434: douta=16'h855a;
8435: douta=16'h7d3b;
8436: douta=16'h7d3a;
8437: douta=16'h7d1a;
8438: douta=16'h7cf9;
8439: douta=16'h74f9;
8440: douta=16'h6c98;
8441: douta=16'h31a8;
8442: douta=16'h326d;
8443: douta=16'h73f1;
8444: douta=16'h7c33;
8445: douta=16'h5b50;
8446: douta=16'h7c33;
8447: douta=16'h42d0;
8448: douta=16'h32b0;
8449: douta=16'h3312;
8450: douta=16'h2a90;
8451: douta=16'h222f;
8452: douta=16'h3290;
8453: douta=16'h5352;
8454: douta=16'h63d4;
8455: douta=16'h63f5;
8456: douta=16'h3a4e;
8457: douta=16'h3a8e;
8458: douta=16'h6350;
8459: douta=16'h7c33;
8460: douta=16'h73d2;
8461: douta=16'h8414;
8462: douta=16'h94d3;
8463: douta=16'h5b4f;
8464: douta=16'had55;
8465: douta=16'hbd74;
8466: douta=16'hde96;
8467: douta=16'h9c90;
8468: douta=16'ha4b1;
8469: douta=16'he697;
8470: douta=16'h7b6d;
8471: douta=16'ha4d1;
8472: douta=16'hcdf4;
8473: douta=16'hce14;
8474: douta=16'h8c0e;
8475: douta=16'h838b;
8476: douta=16'h7b2a;
8477: douta=16'h836a;
8478: douta=16'h93ec;
8479: douta=16'h8b8a;
8480: douta=16'hb4ad;
8481: douta=16'hb48b;
8482: douta=16'hc54f;
8483: douta=16'hcd90;
8484: douta=16'hddf3;
8485: douta=16'he654;
8486: douta=16'he654;
8487: douta=16'hde13;
8488: douta=16'hddf2;
8489: douta=16'hd5b1;
8490: douta=16'hcd50;
8491: douta=16'hbcef;
8492: douta=16'hb48e;
8493: douta=16'h8b69;
8494: douta=16'hc550;
8495: douta=16'hbd30;
8496: douta=16'hac8f;
8497: douta=16'h734c;
8498: douta=16'h6aec;
8499: douta=16'h940e;
8500: douta=16'h7bae;
8501: douta=16'h422a;
8502: douta=16'h29a9;
8503: douta=16'h31c9;
8504: douta=16'h1926;
8505: douta=16'h10e5;
8506: douta=16'h10c4;
8507: douta=16'h1905;
8508: douta=16'h10c4;
8509: douta=16'h10c3;
8510: douta=16'h10c4;
8511: douta=16'h0000;
8512: douta=16'h0062;
8513: douta=16'h1106;
8514: douta=16'h2169;
8515: douta=16'h0063;
8516: douta=16'h29a7;
8517: douta=16'h0000;
8518: douta=16'h3186;
8519: douta=16'h734c;
8520: douta=16'h83ad;
8521: douta=16'h630b;
8522: douta=16'h5aec;
8523: douta=16'h39e9;
8524: douta=16'h4aac;
8525: douta=16'h1147;
8526: douta=16'h7bce;
8527: douta=16'h634e;
8528: douta=16'h426c;
8529: douta=16'h426b;
8530: douta=16'h1128;
8531: douta=16'h0044;
8532: douta=16'h08e6;
8533: douta=16'h31c8;
8534: douta=16'h2167;
8535: douta=16'ha44e;
8536: douta=16'ha5dc;
8537: douta=16'h8d39;
8538: douta=16'h8d59;
8539: douta=16'h957a;
8540: douta=16'h9d9a;
8541: douta=16'h9579;
8542: douta=16'h9dbb;
8543: douta=16'hadfc;
8544: douta=16'h6c14;
8545: douta=16'h53b4;
8546: douta=16'h6435;
8547: douta=16'h6cb7;
8548: douta=16'hae1c;
8549: douta=16'h957a;
8550: douta=16'h9d7a;
8551: douta=16'h959b;
8552: douta=16'h957b;
8553: douta=16'h8d5a;
8554: douta=16'h95bb;
8555: douta=16'h8d5a;
8556: douta=16'h955b;
8557: douta=16'h957a;
8558: douta=16'h959b;
8559: douta=16'h74b8;
8560: douta=16'h955a;
8561: douta=16'h7cd9;
8562: douta=16'h84f9;
8563: douta=16'h8d5a;
8564: douta=16'h6c77;
8565: douta=16'h955a;
8566: douta=16'h9ddb;
8567: douta=16'hbe9e;
8568: douta=16'h7c76;
8569: douta=16'h6c36;
8570: douta=16'h6c56;
8571: douta=16'h5bd5;
8572: douta=16'h6c76;
8573: douta=16'h6436;
8574: douta=16'h5393;
8575: douta=16'h5394;
8576: douta=16'h6416;
8577: douta=16'h4b32;
8578: douta=16'h42d0;
8579: douta=16'h6cb9;
8580: douta=16'h753b;
8581: douta=16'h6458;
8582: douta=16'h6457;
8583: douta=16'h855b;
8584: douta=16'h5393;
8585: douta=16'h4b53;
8586: douta=16'h5bd4;
8587: douta=16'h7cd9;
8588: douta=16'h7497;
8589: douta=16'h7477;
8590: douta=16'h84d8;
8591: douta=16'h7c77;
8592: douta=16'h63f5;
8593: douta=16'h7c97;
8594: douta=16'h7c96;
8595: douta=16'h84b7;
8596: douta=16'h6bf4;
8597: douta=16'h6c35;
8598: douta=16'h7434;
8599: douta=16'h5bf5;
8600: douta=16'h5373;
8601: douta=16'h4b93;
8602: douta=16'h3a90;
8603: douta=16'h3b13;
8604: douta=16'h5c78;
8605: douta=16'h5c38;
8606: douta=16'h5c58;
8607: douta=16'h751b;
8608: douta=16'h6458;
8609: douta=16'h6458;
8610: douta=16'h6478;
8611: douta=16'h74fa;
8612: douta=16'h74da;
8613: douta=16'h7d1a;
8614: douta=16'h855b;
8615: douta=16'h74d9;
8616: douta=16'h74fa;
8617: douta=16'h7cfa;
8618: douta=16'h7d3a;
8619: douta=16'h7d3a;
8620: douta=16'h7d1a;
8621: douta=16'h7d3b;
8622: douta=16'h7d3a;
8623: douta=16'h7d3a;
8624: douta=16'h7499;
8625: douta=16'h7cfa;
8626: douta=16'h6cb9;
8627: douta=16'h7cd9;
8628: douta=16'h853b;
8629: douta=16'h7d1a;
8630: douta=16'h7d1a;
8631: douta=16'h7d3b;
8632: douta=16'h5bf5;
8633: douta=16'h1906;
8634: douta=16'h9d35;
8635: douta=16'h9518;
8636: douta=16'h63d3;
8637: douta=16'h8cf6;
8638: douta=16'h5b50;
8639: douta=16'h6bb1;
8640: douta=16'h4353;
8641: douta=16'h3b53;
8642: douta=16'h3291;
8643: douta=16'h3b12;
8644: douta=16'h5bd4;
8645: douta=16'h5b93;
8646: douta=16'h5bb4;
8647: douta=16'h5372;
8648: douta=16'h6392;
8649: douta=16'h6bf3;
8650: douta=16'h6370;
8651: douta=16'h7412;
8652: douta=16'h6bb1;
8653: douta=16'h634f;
8654: douta=16'hc5f7;
8655: douta=16'ha515;
8656: douta=16'h7390;
8657: douta=16'hb553;
8658: douta=16'hc5b4;
8659: douta=16'hcdf4;
8660: douta=16'hc5d5;
8661: douta=16'hde76;
8662: douta=16'h6aea;
8663: douta=16'h738c;
8664: douta=16'hacd1;
8665: douta=16'hf77a;
8666: douta=16'hbd94;
8667: douta=16'h838a;
8668: douta=16'h8b6a;
8669: douta=16'h8b6a;
8670: douta=16'h93cb;
8671: douta=16'h93cb;
8672: douta=16'hb4ac;
8673: douta=16'hb4ac;
8674: douta=16'hcd6f;
8675: douta=16'hd5b1;
8676: douta=16'he613;
8677: douta=16'he655;
8678: douta=16'he654;
8679: douta=16'hddf2;
8680: douta=16'hddf2;
8681: douta=16'hcd90;
8682: douta=16'hbcee;
8683: douta=16'hb48e;
8684: douta=16'h9bcb;
8685: douta=16'h8348;
8686: douta=16'hac8e;
8687: douta=16'hbd10;
8688: douta=16'hacaf;
8689: douta=16'h83cd;
8690: douta=16'h7b4c;
8691: douta=16'h9c4f;
8692: douta=16'h8bee;
8693: douta=16'h3a0a;
8694: douta=16'h2168;
8695: douta=16'h31a9;
8696: douta=16'h2168;
8697: douta=16'h1905;
8698: douta=16'h2966;
8699: douta=16'h18e5;
8700: douta=16'h18e5;
8701: douta=16'h10c4;
8702: douta=16'h1905;
8703: douta=16'h10c4;
8704: douta=16'h0000;
8705: douta=16'h0062;
8706: douta=16'h21ca;
8707: douta=16'h424a;
8708: douta=16'h2987;
8709: douta=16'h39c6;
8710: douta=16'h0883;
8711: douta=16'h5aaa;
8712: douta=16'h83cd;
8713: douta=16'h736d;
8714: douta=16'h2967;
8715: douta=16'h83ce;
8716: douta=16'h1128;
8717: douta=16'h0064;
8718: douta=16'h29ca;
8719: douta=16'h320a;
8720: douta=16'h31c9;
8721: douta=16'ha4f1;
8722: douta=16'h73d0;
8723: douta=16'h426b;
8724: douta=16'h4a8b;
8725: douta=16'h1968;
8726: douta=16'h08a5;
8727: douta=16'h6289;
8728: douta=16'h9d9a;
8729: douta=16'h8d19;
8730: douta=16'h8d59;
8731: douta=16'h9559;
8732: douta=16'h9dba;
8733: douta=16'ha59a;
8734: douta=16'h957a;
8735: douta=16'h9d9a;
8736: douta=16'hae1c;
8737: douta=16'h7476;
8738: douta=16'h5394;
8739: douta=16'h4b53;
8740: douta=16'h9dbb;
8741: douta=16'h959b;
8742: douta=16'ha5db;
8743: douta=16'h959a;
8744: douta=16'h8d5a;
8745: douta=16'h9ddb;
8746: douta=16'h8d3a;
8747: douta=16'h9ddc;
8748: douta=16'h9ddc;
8749: douta=16'h957b;
8750: douta=16'h957a;
8751: douta=16'h957a;
8752: douta=16'h7cb8;
8753: douta=16'h7cf8;
8754: douta=16'h74b8;
8755: douta=16'h8519;
8756: douta=16'h8d5a;
8757: douta=16'h959b;
8758: douta=16'h53b4;
8759: douta=16'h6c77;
8760: douta=16'hbebe;
8761: douta=16'h52ce;
8762: douta=16'h324c;
8763: douta=16'h21cb;
8764: douta=16'h4bd4;
8765: douta=16'h4353;
8766: douta=16'h4b74;
8767: douta=16'h4b53;
8768: douta=16'h3af2;
8769: douta=16'h5373;
8770: douta=16'h63d4;
8771: douta=16'h42b0;
8772: douta=16'h5b93;
8773: douta=16'h53d4;
8774: douta=16'h42f2;
8775: douta=16'h6c78;
8776: douta=16'h6416;
8777: douta=16'h6416;
8778: douta=16'h5bd4;
8779: douta=16'h7cf9;
8780: douta=16'h7d3a;
8781: douta=16'h8d5b;
8782: douta=16'h7497;
8783: douta=16'h7c97;
8784: douta=16'h7c97;
8785: douta=16'h84f8;
8786: douta=16'h7455;
8787: douta=16'h7434;
8788: douta=16'h6bd3;
8789: douta=16'h73f4;
8790: douta=16'h4acd;
8791: douta=16'h3aaf;
8792: douta=16'h4373;
8793: douta=16'h4bd6;
8794: douta=16'h4bd5;
8795: douta=16'h4395;
8796: douta=16'h5c58;
8797: douta=16'h6cb9;
8798: douta=16'h6478;
8799: douta=16'h5c58;
8800: douta=16'h751a;
8801: douta=16'h4395;
8802: douta=16'h5c16;
8803: douta=16'h74b9;
8804: douta=16'h7cfa;
8805: douta=16'h857b;
8806: douta=16'h857b;
8807: douta=16'h8d7c;
8808: douta=16'h7d3a;
8809: douta=16'h7d3a;
8810: douta=16'h857c;
8811: douta=16'h7d1a;
8812: douta=16'h855b;
8813: douta=16'h855b;
8814: douta=16'h7d3a;
8815: douta=16'h857b;
8816: douta=16'h7d3b;
8817: douta=16'h7cfa;
8818: douta=16'h855b;
8819: douta=16'h6457;
8820: douta=16'h7cfa;
8821: douta=16'h8d9c;
8822: douta=16'h7cf9;
8823: douta=16'h7d1a;
8824: douta=16'h7cd9;
8825: douta=16'h2126;
8826: douta=16'h42ef;
8827: douta=16'h4b30;
8828: douta=16'h6bb1;
8829: douta=16'h7c33;
8830: douta=16'h42ce;
8831: douta=16'h5b71;
8832: douta=16'h32d1;
8833: douta=16'h3b53;
8834: douta=16'h4374;
8835: douta=16'h222f;
8836: douta=16'h6436;
8837: douta=16'h63f4;
8838: douta=16'h7456;
8839: douta=16'h42d0;
8840: douta=16'h6bd3;
8841: douta=16'h52f0;
8842: douta=16'h6371;
8843: douta=16'h73f2;
8844: douta=16'h6391;
8845: douta=16'h632f;
8846: douta=16'ha515;
8847: douta=16'hd638;
8848: douta=16'h8411;
8849: douta=16'h9c91;
8850: douta=16'ha4b1;
8851: douta=16'hbd94;
8852: douta=16'hd657;
8853: douta=16'h942f;
8854: douta=16'ha4d3;
8855: douta=16'hb595;
8856: douta=16'h8bee;
8857: douta=16'h7b2a;
8858: douta=16'h7b4a;
8859: douta=16'h93cb;
8860: douta=16'h8b6a;
8861: douta=16'ha42c;
8862: douta=16'h9beb;
8863: douta=16'ha40c;
8864: douta=16'hbcad;
8865: douta=16'hcd6f;
8866: douta=16'hddf3;
8867: douta=16'hee75;
8868: douta=16'he655;
8869: douta=16'hddf2;
8870: douta=16'he613;
8871: douta=16'hd571;
8872: douta=16'hd591;
8873: douta=16'hcd6f;
8874: douta=16'ha42d;
8875: douta=16'h8308;
8876: douta=16'hb4ce;
8877: douta=16'ha40c;
8878: douta=16'hcd91;
8879: douta=16'hcdb2;
8880: douta=16'hc530;
8881: douta=16'hac8f;
8882: douta=16'h9c4e;
8883: douta=16'ha48f;
8884: douta=16'h8bef;
8885: douta=16'h52ac;
8886: douta=16'h5acc;
8887: douta=16'h424b;
8888: douta=16'h31ea;
8889: douta=16'h2188;
8890: douta=16'h10e6;
8891: douta=16'h422a;
8892: douta=16'h4a4a;
8893: douta=16'h10e4;
8894: douta=16'h10c4;
8895: douta=16'h10e5;
8896: douta=16'h10e5;
8897: douta=16'h2968;
8898: douta=16'h0000;
8899: douta=16'h1107;
8900: douta=16'h5b0e;
8901: douta=16'h5b2f;
8902: douta=16'h4a49;
8903: douta=16'h31a7;
8904: douta=16'h5269;
8905: douta=16'h4a89;
8906: douta=16'h3966;
8907: douta=16'h7bcc;
8908: douta=16'h29a9;
8909: douta=16'h29a9;
8910: douta=16'h10e6;
8911: douta=16'h08e6;
8912: douta=16'h3a2a;
8913: douta=16'h5b0d;
8914: douta=16'h21aa;
8915: douta=16'h4a8c;
8916: douta=16'h2a0c;
8917: douta=16'h1148;
8918: douta=16'h0044;
8919: douta=16'h838c;
8920: douta=16'h9d79;
8921: douta=16'h8d18;
8922: douta=16'h8d39;
8923: douta=16'h959a;
8924: douta=16'h7cb7;
8925: douta=16'h8d39;
8926: douta=16'h9559;
8927: douta=16'h9ddb;
8928: douta=16'h84f8;
8929: douta=16'h9579;
8930: douta=16'h9d9a;
8931: douta=16'h9559;
8932: douta=16'ha5fb;
8933: douta=16'ha5db;
8934: douta=16'h7c76;
8935: douta=16'h6416;
8936: douta=16'h7cd8;
8937: douta=16'h8519;
8938: douta=16'h957a;
8939: douta=16'h955a;
8940: douta=16'h9dbb;
8941: douta=16'h8d5a;
8942: douta=16'h7cf9;
8943: douta=16'h959b;
8944: douta=16'h8d5b;
8945: douta=16'hae1b;
8946: douta=16'hae1c;
8947: douta=16'h7cb8;
8948: douta=16'h8d39;
8949: douta=16'hb67d;
8950: douta=16'h8497;
8951: douta=16'h7cb7;
8952: douta=16'h84d8;
8953: douta=16'h834b;
8954: douta=16'h1105;
8955: douta=16'h18e5;
8956: douta=16'h5373;
8957: douta=16'h53d5;
8958: douta=16'h5bf5;
8959: douta=16'h5bf5;
8960: douta=16'h6457;
8961: douta=16'h63f5;
8962: douta=16'h5b93;
8963: douta=16'h5b93;
8964: douta=16'h6bf5;
8965: douta=16'h42cf;
8966: douta=16'h63b3;
8967: douta=16'h5352;
8968: douta=16'h7d1a;
8969: douta=16'h5c37;
8970: douta=16'h6457;
8971: douta=16'h5c16;
8972: douta=16'h6437;
8973: douta=16'h6436;
8974: douta=16'h63f5;
8975: douta=16'h7cb7;
8976: douta=16'h84d7;
8977: douta=16'h6c35;
8978: douta=16'h6c14;
8979: douta=16'h7413;
8980: douta=16'h73f1;
8981: douta=16'h4208;
8982: douta=16'h2126;
8983: douta=16'h10e5;
8984: douta=16'h3b34;
8985: douta=16'h4bb6;
8986: douta=16'h4bd6;
8987: douta=16'h53f7;
8988: douta=16'h4bf6;
8989: douta=16'h6479;
8990: douta=16'h5c78;
8991: douta=16'h3b33;
8992: douta=16'h6458;
8993: douta=16'h74fa;
8994: douta=16'h7d5b;
8995: douta=16'h751a;
8996: douta=16'h6cb9;
8997: douta=16'h857b;
8998: douta=16'h6c58;
8999: douta=16'h6c78;
9000: douta=16'h6c98;
9001: douta=16'h853a;
9002: douta=16'h8d9c;
9003: douta=16'h857b;
9004: douta=16'h857c;
9005: douta=16'h8d9c;
9006: douta=16'h8d9c;
9007: douta=16'h7d1a;
9008: douta=16'h7d3a;
9009: douta=16'h7d3a;
9010: douta=16'h7d1a;
9011: douta=16'h855b;
9012: douta=16'h855b;
9013: douta=16'h8d5b;
9014: douta=16'h7cf9;
9015: douta=16'h6478;
9016: douta=16'h7cfa;
9017: douta=16'h2146;
9018: douta=16'h5b72;
9019: douta=16'h9cd5;
9020: douta=16'h8cb4;
9021: douta=16'ha538;
9022: douta=16'h63b3;
9023: douta=16'h5372;
9024: douta=16'h3b34;
9025: douta=16'h222f;
9026: douta=16'h3333;
9027: douta=16'h2a90;
9028: douta=16'h6cb9;
9029: douta=16'h53d4;
9030: douta=16'h7476;
9031: douta=16'h6c56;
9032: douta=16'h5331;
9033: douta=16'h6bd3;
9034: douta=16'h7c34;
9035: douta=16'h8c54;
9036: douta=16'h7413;
9037: douta=16'h7c12;
9038: douta=16'had56;
9039: douta=16'h8c93;
9040: douta=16'h7bcf;
9041: douta=16'h8c50;
9042: douta=16'hc594;
9043: douta=16'hd657;
9044: douta=16'hd657;
9045: douta=16'hdeb7;
9046: douta=16'h6b2c;
9047: douta=16'h8c71;
9048: douta=16'h8c10;
9049: douta=16'h8b8b;
9050: douta=16'h8bab;
9051: douta=16'h8349;
9052: douta=16'h8b8b;
9053: douta=16'hac6b;
9054: douta=16'hb4ad;
9055: douta=16'hb48d;
9056: douta=16'hd56f;
9057: douta=16'hd5b1;
9058: douta=16'he675;
9059: douta=16'he675;
9060: douta=16'he675;
9061: douta=16'hddf3;
9062: douta=16'hddf3;
9063: douta=16'he613;
9064: douta=16'hc52f;
9065: douta=16'hbcae;
9066: douta=16'hbcce;
9067: douta=16'h9c0c;
9068: douta=16'hb4ae;
9069: douta=16'hacad;
9070: douta=16'hcd90;
9071: douta=16'hd5d2;
9072: douta=16'hcd70;
9073: douta=16'hbcf0;
9074: douta=16'hb4d0;
9075: douta=16'hac8f;
9076: douta=16'h942f;
9077: douta=16'h736e;
9078: douta=16'h7b6f;
9079: douta=16'h52ce;
9080: douta=16'h428c;
9081: douta=16'h3a2c;
9082: douta=16'h21a9;
9083: douta=16'h1906;
9084: douta=16'h08c5;
9085: douta=16'h0063;
9086: douta=16'h18a4;
9087: douta=16'h10e4;
9088: douta=16'h1084;
9089: douta=16'h08a4;
9090: douta=16'h2146;
9091: douta=16'h0000;
9092: douta=16'h2988;
9093: douta=16'h5b50;
9094: douta=16'h6baf;
9095: douta=16'h0001;
9096: douta=16'h52ca;
9097: douta=16'h08c3;
9098: douta=16'h62aa;
9099: douta=16'h2146;
9100: douta=16'h3186;
9101: douta=16'h6b4c;
9102: douta=16'h5269;
9103: douta=16'h7b8d;
9104: douta=16'hb532;
9105: douta=16'h4a4b;
9106: douta=16'h1948;
9107: douta=16'h636f;
9108: douta=16'h21a9;
9109: douta=16'h426c;
9110: douta=16'h7bef;
9111: douta=16'h8c0f;
9112: douta=16'h8d39;
9113: douta=16'h84b7;
9114: douta=16'h8d18;
9115: douta=16'h8d39;
9116: douta=16'h9579;
9117: douta=16'ha5ba;
9118: douta=16'h8518;
9119: douta=16'h8d39;
9120: douta=16'h8d38;
9121: douta=16'h9579;
9122: douta=16'ha5ba;
9123: douta=16'h9579;
9124: douta=16'h9d9a;
9125: douta=16'h9d9a;
9126: douta=16'h9dba;
9127: douta=16'hae3c;
9128: douta=16'h8d39;
9129: douta=16'h9d59;
9130: douta=16'h5bf6;
9131: douta=16'h9dbb;
9132: douta=16'ha5dc;
9133: douta=16'h957a;
9134: douta=16'h95bb;
9135: douta=16'ha5fc;
9136: douta=16'h853a;
9137: douta=16'h6c58;
9138: douta=16'h7cf9;
9139: douta=16'h8519;
9140: douta=16'ha5fc;
9141: douta=16'h74b8;
9142: douta=16'h7c76;
9143: douta=16'h8518;
9144: douta=16'ha5db;
9145: douta=16'h8bad;
9146: douta=16'h1925;
9147: douta=16'h1905;
9148: douta=16'h6c15;
9149: douta=16'h4b32;
9150: douta=16'h7497;
9151: douta=16'h7cd9;
9152: douta=16'h7497;
9153: douta=16'h7cd8;
9154: douta=16'h6c15;
9155: douta=16'h7cb7;
9156: douta=16'h6c35;
9157: douta=16'h7476;
9158: douta=16'h6415;
9159: douta=16'h4311;
9160: douta=16'h6415;
9161: douta=16'h5b73;
9162: douta=16'h5b94;
9163: douta=16'h6437;
9164: douta=16'h6c77;
9165: douta=16'h7cb8;
9166: douta=16'h63d4;
9167: douta=16'h5bb3;
9168: douta=16'h7c56;
9169: douta=16'h63d3;
9170: douta=16'h9d9a;
9171: douta=16'h84d7;
9172: douta=16'h6bd1;
9173: douta=16'h2967;
9174: douta=16'h1905;
9175: douta=16'h0884;
9176: douta=16'h7cd9;
9177: douta=16'h7477;
9178: douta=16'h6457;
9179: douta=16'h6cb9;
9180: douta=16'h5c37;
9181: douta=16'h5c58;
9182: douta=16'h6479;
9183: douta=16'h6499;
9184: douta=16'h74d9;
9185: douta=16'h5c37;
9186: douta=16'h53d5;
9187: douta=16'h6437;
9188: douta=16'h74f9;
9189: douta=16'h74d9;
9190: douta=16'h74d9;
9191: douta=16'h7d3a;
9192: douta=16'h7d1a;
9193: douta=16'h7477;
9194: douta=16'h6416;
9195: douta=16'h7d3a;
9196: douta=16'h853b;
9197: douta=16'h8d9c;
9198: douta=16'h7d3a;
9199: douta=16'h8d5b;
9200: douta=16'h7d1a;
9201: douta=16'h7d3a;
9202: douta=16'h74b9;
9203: douta=16'h7cd9;
9204: douta=16'h7d1a;
9205: douta=16'h8d9b;
9206: douta=16'h853a;
9207: douta=16'h7d1a;
9208: douta=16'h7498;
9209: douta=16'h39ea;
9210: douta=16'hb5b8;
9211: douta=16'hb5b8;
9212: douta=16'h7413;
9213: douta=16'h42af;
9214: douta=16'h8c94;
9215: douta=16'h9517;
9216: douta=16'h3b13;
9217: douta=16'h3b33;
9218: douta=16'h4b94;
9219: douta=16'h2a6f;
9220: douta=16'h53d5;
9221: douta=16'h4b73;
9222: douta=16'h63d4;
9223: douta=16'h7477;
9224: douta=16'h5b72;
9225: douta=16'h4b10;
9226: douta=16'h5b91;
9227: douta=16'h7c13;
9228: douta=16'h8473;
9229: douta=16'h8c73;
9230: douta=16'had34;
9231: douta=16'h5b2f;
9232: douta=16'h9c92;
9233: douta=16'hb574;
9234: douta=16'h9c90;
9235: douta=16'h9c91;
9236: douta=16'hbd94;
9237: douta=16'hbd94;
9238: douta=16'hb574;
9239: douta=16'hbe17;
9240: douta=16'h6b2b;
9241: douta=16'h8bab;
9242: douta=16'h838a;
9243: douta=16'h8b8b;
9244: douta=16'h9bca;
9245: douta=16'hac8c;
9246: douta=16'hb4ad;
9247: douta=16'hbcad;
9248: douta=16'hd5b0;
9249: douta=16'hde12;
9250: douta=16'hee96;
9251: douta=16'he675;
9252: douta=16'he634;
9253: douta=16'hddf2;
9254: douta=16'hd5d1;
9255: douta=16'hddb2;
9256: douta=16'h9c0d;
9257: douta=16'hc50f;
9258: douta=16'h8b8a;
9259: douta=16'h93aa;
9260: douta=16'ha44d;
9261: douta=16'hb4ad;
9262: douta=16'hcd91;
9263: douta=16'hd5d2;
9264: douta=16'hcd71;
9265: douta=16'hc530;
9266: douta=16'hbd10;
9267: douta=16'hac8f;
9268: douta=16'h9450;
9269: douta=16'h7b8f;
9270: douta=16'h7b8f;
9271: douta=16'h52ce;
9272: douta=16'h4acd;
9273: douta=16'h428d;
9274: douta=16'h29eb;
9275: douta=16'h29a9;
9276: douta=16'h1948;
9277: douta=16'h41e9;
9278: douta=16'h10a4;
9279: douta=16'h10c5;
9280: douta=16'h1084;
9281: douta=16'h1083;
9282: douta=16'h18e5;
9283: douta=16'h0000;
9284: douta=16'h0000;
9285: douta=16'h29ca;
9286: douta=16'h42ad;
9287: douta=16'h3166;
9288: douta=16'h0862;
9289: douta=16'h0000;
9290: douta=16'h18c3;
9291: douta=16'h2125;
9292: douta=16'h2105;
9293: douta=16'h3a09;
9294: douta=16'h4208;
9295: douta=16'h2988;
9296: douta=16'h9c70;
9297: douta=16'h31a8;
9298: douta=16'h5acd;
9299: douta=16'h4aad;
9300: douta=16'h424c;
9301: douta=16'h29a9;
9302: douta=16'h3a6b;
9303: douta=16'h628a;
9304: douta=16'h9d9a;
9305: douta=16'h9559;
9306: douta=16'h8d18;
9307: douta=16'h8d38;
9308: douta=16'h9559;
9309: douta=16'h8d18;
9310: douta=16'h8d18;
9311: douta=16'h8d18;
9312: douta=16'h9579;
9313: douta=16'h959a;
9314: douta=16'h959a;
9315: douta=16'h957a;
9316: douta=16'h84f8;
9317: douta=16'ha5ba;
9318: douta=16'h957a;
9319: douta=16'ha5fa;
9320: douta=16'hb63b;
9321: douta=16'hbe7c;
9322: douta=16'h8cf8;
9323: douta=16'h6457;
9324: douta=16'h7478;
9325: douta=16'h957b;
9326: douta=16'h7cf9;
9327: douta=16'h8539;
9328: douta=16'hbe9d;
9329: douta=16'h851a;
9330: douta=16'h8d7b;
9331: douta=16'h7498;
9332: douta=16'h955b;
9333: douta=16'h8d5a;
9334: douta=16'h63f5;
9335: douta=16'h5b93;
9336: douta=16'h8d19;
9337: douta=16'h93ef;
9338: douta=16'h2146;
9339: douta=16'h18e5;
9340: douta=16'ha5bb;
9341: douta=16'h8d18;
9342: douta=16'h6415;
9343: douta=16'h8539;
9344: douta=16'h8519;
9345: douta=16'h853a;
9346: douta=16'h7477;
9347: douta=16'h8d39;
9348: douta=16'h955a;
9349: douta=16'h7cd8;
9350: douta=16'h855b;
9351: douta=16'h7cd8;
9352: douta=16'h5373;
9353: douta=16'h6435;
9354: douta=16'h6c15;
9355: douta=16'h7cd9;
9356: douta=16'h74b7;
9357: douta=16'h6c36;
9358: douta=16'h84b7;
9359: douta=16'h63f4;
9360: douta=16'h63d3;
9361: douta=16'h63b3;
9362: douta=16'h6c35;
9363: douta=16'h957a;
9364: douta=16'h6bb1;
9365: douta=16'h2105;
9366: douta=16'h18e5;
9367: douta=16'h10e5;
9368: douta=16'h7cb8;
9369: douta=16'h6c77;
9370: douta=16'h7498;
9371: douta=16'h6458;
9372: douta=16'h6c99;
9373: douta=16'h4bd6;
9374: douta=16'h53d6;
9375: douta=16'h5c17;
9376: douta=16'h6478;
9377: douta=16'h6cb9;
9378: douta=16'h74d9;
9379: douta=16'h6457;
9380: douta=16'h6cb8;
9381: douta=16'h7d1a;
9382: douta=16'h6c98;
9383: douta=16'h7d1a;
9384: douta=16'h851a;
9385: douta=16'h851a;
9386: douta=16'h6c37;
9387: douta=16'h7cb9;
9388: douta=16'h74b9;
9389: douta=16'h7cf9;
9390: douta=16'h8dbc;
9391: douta=16'h7cda;
9392: douta=16'h8dbc;
9393: douta=16'h857b;
9394: douta=16'h8d7c;
9395: douta=16'h7d3b;
9396: douta=16'h855b;
9397: douta=16'h853a;
9398: douta=16'h7cd9;
9399: douta=16'h7d1a;
9400: douta=16'h7477;
9401: douta=16'h2968;
9402: douta=16'h7433;
9403: douta=16'hb5d8;
9404: douta=16'h73f3;
9405: douta=16'h7434;
9406: douta=16'h42d0;
9407: douta=16'h52ce;
9408: douta=16'h2a0d;
9409: douta=16'h4374;
9410: douta=16'h5c58;
9411: douta=16'h4bd6;
9412: douta=16'h3b33;
9413: douta=16'h53f6;
9414: douta=16'h63f5;
9415: douta=16'h7478;
9416: douta=16'h7436;
9417: douta=16'h63b2;
9418: douta=16'h5b93;
9419: douta=16'h4aef;
9420: douta=16'h73d2;
9421: douta=16'h8cb4;
9422: douta=16'hbdd8;
9423: douta=16'h8433;
9424: douta=16'h8411;
9425: douta=16'hcdf6;
9426: douta=16'hc5f5;
9427: douta=16'hd616;
9428: douta=16'hd657;
9429: douta=16'hb574;
9430: douta=16'h946f;
9431: douta=16'h938b;
9432: douta=16'h8b8b;
9433: douta=16'h9bcb;
9434: douta=16'hac4b;
9435: douta=16'hac6c;
9436: douta=16'hcd4e;
9437: douta=16'hbced;
9438: douta=16'hcd4e;
9439: douta=16'hd590;
9440: douta=16'he654;
9441: douta=16'hee96;
9442: douta=16'he654;
9443: douta=16'he654;
9444: douta=16'he654;
9445: douta=16'hde34;
9446: douta=16'hb4cf;
9447: douta=16'hbcd0;
9448: douta=16'h7b29;
9449: douta=16'h834a;
9450: douta=16'hd570;
9451: douta=16'hbd0e;
9452: douta=16'hbd2f;
9453: douta=16'hc52f;
9454: douta=16'hddf3;
9455: douta=16'hd5d2;
9456: douta=16'hd591;
9457: douta=16'hcd71;
9458: douta=16'hcd71;
9459: douta=16'hb4d0;
9460: douta=16'h9c50;
9461: douta=16'h8c10;
9462: douta=16'h7bcf;
9463: douta=16'h636f;
9464: douta=16'h5b2e;
9465: douta=16'h52cf;
9466: douta=16'h29eb;
9467: douta=16'h31eb;
9468: douta=16'h29ca;
9469: douta=16'h10e6;
9470: douta=16'h424a;
9471: douta=16'h10a4;
9472: douta=16'h10a4;
9473: douta=16'h10e4;
9474: douta=16'h1904;
9475: douta=16'h10c4;
9476: douta=16'h1906;
9477: douta=16'h2146;
9478: douta=16'h29eb;
9479: douta=16'h5b0e;
9480: douta=16'h3a6b;
9481: douta=16'h5a49;
9482: douta=16'h944d;
9483: douta=16'h3165;
9484: douta=16'h8bed;
9485: douta=16'h736c;
9486: douta=16'h5aa9;
9487: douta=16'h2146;
9488: douta=16'h0885;
9489: douta=16'h21a9;
9490: douta=16'h8c2f;
9491: douta=16'h5aab;
9492: douta=16'ha4d1;
9493: douta=16'h632d;
9494: douta=16'h426c;
9495: douta=16'h736e;
9496: douta=16'hb65c;
9497: douta=16'h9579;
9498: douta=16'h8d38;
9499: douta=16'h84f7;
9500: douta=16'h8d58;
9501: douta=16'h8d58;
9502: douta=16'h7cb7;
9503: douta=16'h84f8;
9504: douta=16'h8d38;
9505: douta=16'h8d39;
9506: douta=16'h9559;
9507: douta=16'h9579;
9508: douta=16'h8d39;
9509: douta=16'h8d39;
9510: douta=16'h9d9a;
9511: douta=16'h9559;
9512: douta=16'h9559;
9513: douta=16'h9dba;
9514: douta=16'h957a;
9515: douta=16'hadfa;
9516: douta=16'h9d9a;
9517: douta=16'ha5fb;
9518: douta=16'h9d9a;
9519: douta=16'h7cd9;
9520: douta=16'h7c97;
9521: douta=16'h957a;
9522: douta=16'hae3c;
9523: douta=16'h84f9;
9524: douta=16'ha5dc;
9525: douta=16'h957a;
9526: douta=16'h7435;
9527: douta=16'h84d7;
9528: douta=16'h7cb7;
9529: douta=16'h8474;
9530: douta=16'h5249;
9531: douta=16'h1905;
9532: douta=16'h5b91;
9533: douta=16'h9559;
9534: douta=16'h8d18;
9535: douta=16'h9579;
9536: douta=16'h9d9a;
9537: douta=16'h9dbb;
9538: douta=16'h8d3a;
9539: douta=16'h8d18;
9540: douta=16'h8d39;
9541: douta=16'h7cb8;
9542: douta=16'h7cf9;
9543: douta=16'h9ddc;
9544: douta=16'h84f9;
9545: douta=16'h7cb7;
9546: douta=16'h84d9;
9547: douta=16'h7cb7;
9548: douta=16'h6c35;
9549: douta=16'h6c14;
9550: douta=16'h84d7;
9551: douta=16'h9559;
9552: douta=16'h84d8;
9553: douta=16'h63d4;
9554: douta=16'h6bf4;
9555: douta=16'h6c35;
9556: douta=16'h39a8;
9557: douta=16'h2126;
9558: douta=16'h1905;
9559: douta=16'h4ad0;
9560: douta=16'h6436;
9561: douta=16'h5bf5;
9562: douta=16'h7498;
9563: douta=16'h6457;
9564: douta=16'h6cb9;
9565: douta=16'h6cda;
9566: douta=16'h751b;
9567: douta=16'h5c16;
9568: douta=16'h74f9;
9569: douta=16'h5c37;
9570: douta=16'h6c78;
9571: douta=16'h74b9;
9572: douta=16'h7cd9;
9573: douta=16'h7cf9;
9574: douta=16'h7498;
9575: douta=16'h74b8;
9576: douta=16'h7cd9;
9577: douta=16'h74b8;
9578: douta=16'h74b8;
9579: douta=16'h7cf9;
9580: douta=16'h8d5b;
9581: douta=16'h7cf9;
9582: douta=16'h851a;
9583: douta=16'h7d1a;
9584: douta=16'h6457;
9585: douta=16'h7cd9;
9586: douta=16'h7d1a;
9587: douta=16'h7d1a;
9588: douta=16'h7cd9;
9589: douta=16'h8d7b;
9590: douta=16'h7cf9;
9591: douta=16'h74b8;
9592: douta=16'h5b73;
9593: douta=16'h84d6;
9594: douta=16'ha598;
9595: douta=16'hbdf9;
9596: douta=16'h94d5;
9597: douta=16'h94b6;
9598: douta=16'h4aee;
9599: douta=16'h0800;
9600: douta=16'h222e;
9601: douta=16'h32f2;
9602: douta=16'h4b54;
9603: douta=16'h4375;
9604: douta=16'h4333;
9605: douta=16'h6458;
9606: douta=16'h5332;
9607: douta=16'h7cb9;
9608: douta=16'h63d4;
9609: douta=16'h4af0;
9610: douta=16'h7475;
9611: douta=16'h5b92;
9612: douta=16'h7c54;
9613: douta=16'h73f4;
9614: douta=16'hb576;
9615: douta=16'ha536;
9616: douta=16'h8c94;
9617: douta=16'hb534;
9618: douta=16'heef9;
9619: douta=16'hbd74;
9620: douta=16'hce36;
9621: douta=16'hc5f6;
9622: douta=16'h8369;
9623: douta=16'h93cb;
9624: douta=16'h938a;
9625: douta=16'hac4c;
9626: douta=16'hbc8b;
9627: douta=16'hbcad;
9628: douta=16'hc52e;
9629: douta=16'hd5b0;
9630: douta=16'hddf2;
9631: douta=16'he654;
9632: douta=16'hee75;
9633: douta=16'he674;
9634: douta=16'he654;
9635: douta=16'he674;
9636: douta=16'hde13;
9637: douta=16'hbcef;
9638: douta=16'hc551;
9639: douta=16'h9c2c;
9640: douta=16'hb4ae;
9641: douta=16'h93ec;
9642: douta=16'h838b;
9643: douta=16'hc550;
9644: douta=16'hde13;
9645: douta=16'hd5f3;
9646: douta=16'hde13;
9647: douta=16'hddf3;
9648: douta=16'hd5b2;
9649: douta=16'hcd71;
9650: douta=16'hcd50;
9651: douta=16'hc530;
9652: douta=16'h9c50;
9653: douta=16'h8c10;
9654: douta=16'h83d0;
9655: douta=16'h6b6f;
9656: douta=16'h6b70;
9657: douta=16'h634f;
9658: douta=16'h5330;
9659: douta=16'h42af;
9660: douta=16'h3a8e;
9661: douta=16'h29eb;
9662: douta=16'h2988;
9663: douta=16'h2126;
9664: douta=16'h10e4;
9665: douta=16'h10e4;
9666: douta=16'h10c3;
9667: douta=16'h10c3;
9668: douta=16'h10a4;
9669: douta=16'h10a4;
9670: douta=16'h10e5;
9671: douta=16'h3acf;
9672: douta=16'h10c6;
9673: douta=16'h08c5;
9674: douta=16'h2167;
9675: douta=16'h6b4b;
9676: douta=16'had11;
9677: douta=16'h39a6;
9678: douta=16'h39c6;
9679: douta=16'h5aca;
9680: douta=16'h4228;
9681: douta=16'h528a;
9682: douta=16'h8c50;
9683: douta=16'h942f;
9684: douta=16'h31c9;
9685: douta=16'h0085;
9686: douta=16'h1105;
9687: douta=16'h524a;
9688: douta=16'h7cd7;
9689: douta=16'h5bb4;
9690: douta=16'h9558;
9691: douta=16'h9559;
9692: douta=16'h9579;
9693: douta=16'hadfb;
9694: douta=16'h8d39;
9695: douta=16'h8d18;
9696: douta=16'h8d18;
9697: douta=16'h84d7;
9698: douta=16'h8d18;
9699: douta=16'h84f8;
9700: douta=16'h7cd7;
9701: douta=16'h957a;
9702: douta=16'h8d39;
9703: douta=16'h9579;
9704: douta=16'h9d9a;
9705: douta=16'h9559;
9706: douta=16'h9559;
9707: douta=16'h9559;
9708: douta=16'ha5db;
9709: douta=16'h9dbb;
9710: douta=16'ha5db;
9711: douta=16'h9dbb;
9712: douta=16'ha5db;
9713: douta=16'h9d9a;
9714: douta=16'h6c15;
9715: douta=16'h7cd9;
9716: douta=16'h9ddc;
9717: douta=16'h8d3a;
9718: douta=16'h8d18;
9719: douta=16'h84f8;
9720: douta=16'h8518;
9721: douta=16'h7435;
9722: douta=16'h838b;
9723: douta=16'h31a7;
9724: douta=16'h31c9;
9725: douta=16'h8cf8;
9726: douta=16'h84f8;
9727: douta=16'h8d39;
9728: douta=16'h9d7a;
9729: douta=16'ha5fb;
9730: douta=16'h957a;
9731: douta=16'h8d39;
9732: douta=16'h955a;
9733: douta=16'h8519;
9734: douta=16'h8d39;
9735: douta=16'h957b;
9736: douta=16'h7cb9;
9737: douta=16'h8539;
9738: douta=16'h8d5a;
9739: douta=16'h8d5a;
9740: douta=16'h957a;
9741: douta=16'h957a;
9742: douta=16'h6bf4;
9743: douta=16'h63d3;
9744: douta=16'h7435;
9745: douta=16'h9559;
9746: douta=16'h8518;
9747: douta=16'h7c55;
9748: douta=16'h2905;
9749: douta=16'h2146;
9750: douta=16'h10c5;
9751: douta=16'h5c15;
9752: douta=16'h5c16;
9753: douta=16'h7d5a;
9754: douta=16'h74d9;
9755: douta=16'h6cb9;
9756: douta=16'h6c79;
9757: douta=16'h6c98;
9758: douta=16'h74da;
9759: douta=16'h6cb9;
9760: douta=16'h6c98;
9761: douta=16'h74d9;
9762: douta=16'h74d9;
9763: douta=16'h74d9;
9764: douta=16'h74b9;
9765: douta=16'h6c56;
9766: douta=16'h74d9;
9767: douta=16'h7d1a;
9768: douta=16'h7498;
9769: douta=16'h63f6;
9770: douta=16'h8d5b;
9771: douta=16'h6c77;
9772: douta=16'h7cd9;
9773: douta=16'h851a;
9774: douta=16'h7478;
9775: douta=16'h7cf9;
9776: douta=16'h853b;
9777: douta=16'h7d1a;
9778: douta=16'h853a;
9779: douta=16'h8519;
9780: douta=16'h7cfa;
9781: douta=16'h853a;
9782: douta=16'h851a;
9783: douta=16'h853a;
9784: douta=16'h29cb;
9785: douta=16'hdefd;
9786: douta=16'h6c15;
9787: douta=16'h8cb6;
9788: douta=16'ha558;
9789: douta=16'h42ae;
9790: douta=16'h73b0;
9791: douta=16'h3a2a;
9792: douta=16'h3ad1;
9793: douta=16'h2a4f;
9794: douta=16'h4374;
9795: douta=16'h32b1;
9796: douta=16'h4374;
9797: douta=16'h53d5;
9798: douta=16'h3290;
9799: douta=16'h6415;
9800: douta=16'h5373;
9801: douta=16'h63b4;
9802: douta=16'h9559;
9803: douta=16'h7414;
9804: douta=16'h73f3;
9805: douta=16'h6bd2;
9806: douta=16'had36;
9807: douta=16'ha537;
9808: douta=16'h9d15;
9809: douta=16'had34;
9810: douta=16'hbd94;
9811: douta=16'hbd95;
9812: douta=16'he6f9;
9813: douta=16'h9cd3;
9814: douta=16'h93cb;
9815: douta=16'h93aa;
9816: douta=16'h93aa;
9817: douta=16'hb48c;
9818: douta=16'hc4cd;
9819: douta=16'hbccd;
9820: douta=16'hcd6f;
9821: douta=16'hddd1;
9822: douta=16'hde33;
9823: douta=16'hee75;
9824: douta=16'he675;
9825: douta=16'hee96;
9826: douta=16'he633;
9827: douta=16'hde34;
9828: douta=16'hddd2;
9829: douta=16'hbcef;
9830: douta=16'hc50f;
9831: douta=16'hb4ae;
9832: douta=16'hb4ce;
9833: douta=16'ha42d;
9834: douta=16'h838b;
9835: douta=16'ha48c;
9836: douta=16'hcd91;
9837: douta=16'hd5d2;
9838: douta=16'hde14;
9839: douta=16'hde13;
9840: douta=16'hd5b2;
9841: douta=16'hcd71;
9842: douta=16'hcd71;
9843: douta=16'hc551;
9844: douta=16'h9c50;
9845: douta=16'h9410;
9846: douta=16'h83cf;
9847: douta=16'h6b6f;
9848: douta=16'h634f;
9849: douta=16'h5b2f;
9850: douta=16'h52ef;
9851: douta=16'h42ef;
9852: douta=16'h42ae;
9853: douta=16'h3a6d;
9854: douta=16'h2189;
9855: douta=16'h6b4e;
9856: douta=16'h10e4;
9857: douta=16'h0883;
9858: douta=16'h10c4;
9859: douta=16'h10e4;
9860: douta=16'h10c4;
9861: douta=16'h10c5;
9862: douta=16'h2146;
9863: douta=16'h0000;
9864: douta=16'h2988;
9865: douta=16'h1947;
9866: douta=16'h10e5;
9867: douta=16'h10c5;
9868: douta=16'h738c;
9869: douta=16'h62ea;
9870: douta=16'h5289;
9871: douta=16'h528a;
9872: douta=16'h10c4;
9873: douta=16'h0043;
9874: douta=16'h6b8e;
9875: douta=16'hb551;
9876: douta=16'h944f;
9877: douta=16'h6b4d;
9878: douta=16'h29c9;
9879: douta=16'h0884;
9880: douta=16'h9539;
9881: douta=16'h7cf7;
9882: douta=16'h7455;
9883: douta=16'h7cb7;
9884: douta=16'h7c96;
9885: douta=16'h7cb7;
9886: douta=16'h9559;
9887: douta=16'h9579;
9888: douta=16'h9579;
9889: douta=16'h8d18;
9890: douta=16'h84d7;
9891: douta=16'h9d9a;
9892: douta=16'h8518;
9893: douta=16'h8d38;
9894: douta=16'h7cb7;
9895: douta=16'h8d18;
9896: douta=16'h9599;
9897: douta=16'h84d7;
9898: douta=16'h8d18;
9899: douta=16'h9d9a;
9900: douta=16'h9d9a;
9901: douta=16'ha5ba;
9902: douta=16'ha5ba;
9903: douta=16'ha5db;
9904: douta=16'h8d5a;
9905: douta=16'hae3c;
9906: douta=16'hb67d;
9907: douta=16'h8d39;
9908: douta=16'h7cd9;
9909: douta=16'h7cf9;
9910: douta=16'h8d39;
9911: douta=16'h84d8;
9912: douta=16'h84f8;
9913: douta=16'h84d7;
9914: douta=16'h93ed;
9915: douta=16'h4a08;
9916: douta=16'h10a5;
9917: douta=16'h6c15;
9918: douta=16'h8d19;
9919: douta=16'h8d39;
9920: douta=16'h8d39;
9921: douta=16'h84b7;
9922: douta=16'ha5ba;
9923: douta=16'h9d9a;
9924: douta=16'h9dbb;
9925: douta=16'h8d5a;
9926: douta=16'h8d59;
9927: douta=16'h8519;
9928: douta=16'h955a;
9929: douta=16'h7456;
9930: douta=16'h6c15;
9931: douta=16'h9559;
9932: douta=16'h9dbb;
9933: douta=16'h8d39;
9934: douta=16'h8cd8;
9935: douta=16'h7c55;
9936: douta=16'h7435;
9937: douta=16'h7c75;
9938: douta=16'h84f8;
9939: douta=16'h8d18;
9940: douta=16'h2105;
9941: douta=16'h2126;
9942: douta=16'h10e5;
9943: douta=16'h5c17;
9944: douta=16'h6437;
9945: douta=16'h6437;
9946: douta=16'h6458;
9947: douta=16'h6cba;
9948: douta=16'h74fa;
9949: douta=16'h74da;
9950: douta=16'h751a;
9951: douta=16'h74fa;
9952: douta=16'h855b;
9953: douta=16'h74b8;
9954: douta=16'h7498;
9955: douta=16'h74b8;
9956: douta=16'h7498;
9957: douta=16'h7cf9;
9958: douta=16'h74b8;
9959: douta=16'h7cd9;
9960: douta=16'h7498;
9961: douta=16'h7498;
9962: douta=16'h7cd8;
9963: douta=16'h8d9b;
9964: douta=16'h7478;
9965: douta=16'h7cd9;
9966: douta=16'h7cd9;
9967: douta=16'h7cd9;
9968: douta=16'h8d5b;
9969: douta=16'h7d1a;
9970: douta=16'h7d3a;
9971: douta=16'h7cda;
9972: douta=16'h8d3a;
9973: douta=16'h8d7b;
9974: douta=16'h855a;
9975: douta=16'h7d3a;
9976: douta=16'h31a9;
9977: douta=16'hb61a;
9978: douta=16'h5bb3;
9979: douta=16'hd69b;
9980: douta=16'h9d37;
9981: douta=16'h532f;
9982: douta=16'h39e8;
9983: douta=16'h4aad;
9984: douta=16'h328f;
9985: douta=16'h2a4f;
9986: douta=16'h3af3;
9987: douta=16'h3b33;
9988: douta=16'h4374;
9989: douta=16'h6457;
9990: douta=16'h4312;
9991: douta=16'h5373;
9992: douta=16'h5bf5;
9993: douta=16'h6415;
9994: douta=16'h84d7;
9995: douta=16'h7c96;
9996: douta=16'h8c94;
9997: douta=16'ha536;
9998: douta=16'h9cb4;
9999: douta=16'hbdd7;
10000: douta=16'hb5b6;
10001: douta=16'had34;
10002: douta=16'h8c31;
10003: douta=16'had76;
10004: douta=16'had13;
10005: douta=16'h832a;
10006: douta=16'hac4b;
10007: douta=16'ha40b;
10008: douta=16'hac4c;
10009: douta=16'hcd4e;
10010: douta=16'hcd0d;
10011: douta=16'hd58f;
10012: douta=16'hde13;
10013: douta=16'hcd90;
10014: douta=16'he654;
10015: douta=16'heeb6;
10016: douta=16'he675;
10017: douta=16'he654;
10018: douta=16'hac6c;
10019: douta=16'hb4ae;
10020: douta=16'hddd1;
10021: douta=16'ha42d;
10022: douta=16'h72a6;
10023: douta=16'h9c2b;
10024: douta=16'hac6d;
10025: douta=16'hac8d;
10026: douta=16'hc50f;
10027: douta=16'hcd71;
10028: douta=16'hd5b2;
10029: douta=16'hddf3;
10030: douta=16'hde34;
10031: douta=16'hde13;
10032: douta=16'hd5b2;
10033: douta=16'hd591;
10034: douta=16'hd591;
10035: douta=16'hc530;
10036: douta=16'hacb1;
10037: douta=16'h9c51;
10038: douta=16'h9430;
10039: douta=16'h7bd1;
10040: douta=16'h73b1;
10041: douta=16'h6b70;
10042: douta=16'h6371;
10043: douta=16'h5b50;
10044: douta=16'h530f;
10045: douta=16'h428d;
10046: douta=16'h3a2c;
10047: douta=16'h320c;
10048: douta=16'h6b2c;
10049: douta=16'h1906;
10050: douta=16'h18e4;
10051: douta=16'h10c4;
10052: douta=16'h10c3;
10053: douta=16'h10e4;
10054: douta=16'h10c4;
10055: douta=16'h10e5;
10056: douta=16'h1906;
10057: douta=16'h2167;
10058: douta=16'h2189;
10059: douta=16'h1946;
10060: douta=16'h0884;
10061: douta=16'h3a07;
10062: douta=16'h08a4;
10063: douta=16'h2947;
10064: douta=16'h944f;
10065: douta=16'h2124;
10066: douta=16'h18a3;
10067: douta=16'h630c;
10068: douta=16'h2146;
10069: douta=16'h8c30;
10070: douta=16'h52cc;
10071: douta=16'h83ed;
10072: douta=16'h6bd2;
10073: douta=16'hae3c;
10074: douta=16'ha5db;
10075: douta=16'h7415;
10076: douta=16'h7cb6;
10077: douta=16'h8cf8;
10078: douta=16'ha5db;
10079: douta=16'h7cb7;
10080: douta=16'h9559;
10081: douta=16'h84f8;
10082: douta=16'hb65b;
10083: douta=16'hb63b;
10084: douta=16'ha5ba;
10085: douta=16'h8d59;
10086: douta=16'h9559;
10087: douta=16'h8d39;
10088: douta=16'h8d18;
10089: douta=16'h9559;
10090: douta=16'ha5ba;
10091: douta=16'h957a;
10092: douta=16'h9559;
10093: douta=16'h9d9a;
10094: douta=16'h957a;
10095: douta=16'h9559;
10096: douta=16'h9dba;
10097: douta=16'ha5ba;
10098: douta=16'h9dba;
10099: douta=16'h9dba;
10100: douta=16'ha5db;
10101: douta=16'h8d5a;
10102: douta=16'hadfb;
10103: douta=16'h8d39;
10104: douta=16'h7c77;
10105: douta=16'h84d8;
10106: douta=16'ha4f2;
10107: douta=16'h8b8b;
10108: douta=16'h10c4;
10109: douta=16'h2167;
10110: douta=16'h7cb8;
10111: douta=16'h9559;
10112: douta=16'ha5db;
10113: douta=16'h84f8;
10114: douta=16'ha5ba;
10115: douta=16'h9d58;
10116: douta=16'h9d79;
10117: douta=16'h84b6;
10118: douta=16'h8d39;
10119: douta=16'h9dbb;
10120: douta=16'ha61c;
10121: douta=16'h9d9a;
10122: douta=16'h9518;
10123: douta=16'h8495;
10124: douta=16'h8cb4;
10125: douta=16'h7c12;
10126: douta=16'h8cd7;
10127: douta=16'h84b7;
10128: douta=16'h8cf8;
10129: douta=16'h84d8;
10130: douta=16'h84d7;
10131: douta=16'h7476;
10132: douta=16'h2146;
10133: douta=16'h1905;
10134: douta=16'h18e5;
10135: douta=16'h8ddf;
10136: douta=16'h4333;
10137: douta=16'h3b12;
10138: douta=16'h6499;
10139: douta=16'h5c58;
10140: douta=16'h6cda;
10141: douta=16'h4b94;
10142: douta=16'h5394;
10143: douta=16'h5c16;
10144: douta=16'h7519;
10145: douta=16'h74d9;
10146: douta=16'h7cd9;
10147: douta=16'h7d19;
10148: douta=16'h7498;
10149: douta=16'h851a;
10150: douta=16'h851a;
10151: douta=16'h853a;
10152: douta=16'h7cd9;
10153: douta=16'h7cd9;
10154: douta=16'h7cd9;
10155: douta=16'h8d5a;
10156: douta=16'h7498;
10157: douta=16'h7498;
10158: douta=16'h8d5a;
10159: douta=16'h6c57;
10160: douta=16'h853a;
10161: douta=16'h853a;
10162: douta=16'h959b;
10163: douta=16'h853a;
10164: douta=16'h8519;
10165: douta=16'h8d7b;
10166: douta=16'h7cf9;
10167: douta=16'h7cf9;
10168: douta=16'h52ac;
10169: douta=16'h8434;
10170: douta=16'hadb9;
10171: douta=16'h7c33;
10172: douta=16'h8495;
10173: douta=16'h3a8f;
10174: douta=16'h0041;
10175: douta=16'ha577;
10176: douta=16'h2106;
10177: douta=16'h2a90;
10178: douta=16'h3af2;
10179: douta=16'h751c;
10180: douta=16'h2a4f;
10181: douta=16'h3b12;
10182: douta=16'h53b4;
10183: douta=16'h63f5;
10184: douta=16'h5bb4;
10185: douta=16'h6c35;
10186: douta=16'h7cb7;
10187: douta=16'h6392;
10188: douta=16'h4ace;
10189: douta=16'h8433;
10190: douta=16'ha536;
10191: douta=16'hbdb7;
10192: douta=16'hc618;
10193: douta=16'h8411;
10194: douta=16'h9493;
10195: douta=16'h834b;
10196: douta=16'h834a;
10197: douta=16'h8b8b;
10198: douta=16'hac2a;
10199: douta=16'hb4ac;
10200: douta=16'hc4ed;
10201: douta=16'hd58f;
10202: douta=16'hd5b0;
10203: douta=16'hddd1;
10204: douta=16'hde13;
10205: douta=16'hee75;
10206: douta=16'hde13;
10207: douta=16'hee95;
10208: douta=16'he634;
10209: douta=16'hde12;
10210: douta=16'hcd71;
10211: douta=16'hbcf0;
10212: douta=16'h9beb;
10213: douta=16'h7285;
10214: douta=16'hb4ce;
10215: douta=16'hbd30;
10216: douta=16'hbd2f;
10217: douta=16'hc54f;
10218: douta=16'hc550;
10219: douta=16'hd5b1;
10220: douta=16'he634;
10221: douta=16'he634;
10222: douta=16'he655;
10223: douta=16'hde13;
10224: douta=16'hddf3;
10225: douta=16'hcd71;
10226: douta=16'hcd50;
10227: douta=16'hc531;
10228: douta=16'hacb1;
10229: douta=16'ha471;
10230: douta=16'h9c51;
10231: douta=16'h8411;
10232: douta=16'h8411;
10233: douta=16'h73d1;
10234: douta=16'h6370;
10235: douta=16'h5b50;
10236: douta=16'h6350;
10237: douta=16'h5330;
10238: douta=16'h6372;
10239: douta=16'h29a9;
10240: douta=16'h10e6;
10241: douta=16'h2146;
10242: douta=16'h39ea;
10243: douta=16'h10a4;
10244: douta=16'h10e4;
10245: douta=16'h10c4;
10246: douta=16'h10c4;
10247: douta=16'h10a3;
10248: douta=16'h10c5;
10249: douta=16'h1084;
10250: douta=16'h0042;
10251: douta=16'h2188;
10252: douta=16'h18c5;
10253: douta=16'h840d;
10254: douta=16'h39a6;
10255: douta=16'h5ac9;
10256: douta=16'h39a7;
10257: douta=16'h3186;
10258: douta=16'hb510;
10259: douta=16'h630c;
10260: douta=16'h2967;
10261: douta=16'h29a9;
10262: douta=16'h2187;
10263: douta=16'h5acb;
10264: douta=16'h6b4d;
10265: douta=16'h7c95;
10266: douta=16'h84d7;
10267: douta=16'h8d38;
10268: douta=16'h84f8;
10269: douta=16'h957a;
10270: douta=16'h7476;
10271: douta=16'h7c97;
10272: douta=16'h84b8;
10273: douta=16'h9dba;
10274: douta=16'h7456;
10275: douta=16'h5352;
10276: douta=16'h84f7;
10277: douta=16'ha5ba;
10278: douta=16'h8d18;
10279: douta=16'ha5ba;
10280: douta=16'h9579;
10281: douta=16'h9579;
10282: douta=16'h9d9a;
10283: douta=16'ha5da;
10284: douta=16'ha5da;
10285: douta=16'h8d59;
10286: douta=16'h9d9a;
10287: douta=16'h9d9a;
10288: douta=16'hadfa;
10289: douta=16'ha5db;
10290: douta=16'h9559;
10291: douta=16'h9d9a;
10292: douta=16'ha5fb;
10293: douta=16'h8d59;
10294: douta=16'h8539;
10295: douta=16'h959a;
10296: douta=16'h957a;
10297: douta=16'h9dbb;
10298: douta=16'h94f6;
10299: douta=16'hbccf;
10300: douta=16'h18e5;
10301: douta=16'h0042;
10302: douta=16'h9ddc;
10303: douta=16'h8d39;
10304: douta=16'h8d39;
10305: douta=16'h84b8;
10306: douta=16'h84d8;
10307: douta=16'h957a;
10308: douta=16'h7c76;
10309: douta=16'h9539;
10310: douta=16'h9d9a;
10311: douta=16'h9559;
10312: douta=16'h8cf8;
10313: douta=16'h9d99;
10314: douta=16'h9d58;
10315: douta=16'h94f6;
10316: douta=16'h8c75;
10317: douta=16'h8d18;
10318: douta=16'h7455;
10319: douta=16'h7455;
10320: douta=16'h84b7;
10321: douta=16'h84f8;
10322: douta=16'h7cd8;
10323: douta=16'h8d7b;
10324: douta=16'h2126;
10325: douta=16'h10e5;
10326: douta=16'h2104;
10327: douta=16'h5c16;
10328: douta=16'h6478;
10329: douta=16'h751a;
10330: douta=16'h5c36;
10331: douta=16'h3b34;
10332: douta=16'h5417;
10333: douta=16'h6cb9;
10334: douta=16'h53f6;
10335: douta=16'h5c16;
10336: douta=16'h6c77;
10337: douta=16'h857b;
10338: douta=16'h8d9c;
10339: douta=16'h6c77;
10340: douta=16'h7498;
10341: douta=16'h7cd9;
10342: douta=16'h7cd9;
10343: douta=16'h7cf9;
10344: douta=16'h853a;
10345: douta=16'h853a;
10346: douta=16'h7cd9;
10347: douta=16'h7cd9;
10348: douta=16'h7cd9;
10349: douta=16'h8d5a;
10350: douta=16'h959b;
10351: douta=16'h74b8;
10352: douta=16'h853a;
10353: douta=16'h8d5a;
10354: douta=16'h7cf9;
10355: douta=16'h853a;
10356: douta=16'h8dbc;
10357: douta=16'h6477;
10358: douta=16'h8d7b;
10359: douta=16'h8d5b;
10360: douta=16'h7c95;
10361: douta=16'hbe3a;
10362: douta=16'h63f4;
10363: douta=16'h7c33;
10364: douta=16'h9d16;
10365: douta=16'h94f6;
10366: douta=16'h7c33;
10367: douta=16'h5310;
10368: douta=16'h2106;
10369: douta=16'h53f7;
10370: douta=16'h32b0;
10371: douta=16'h4bb5;
10372: douta=16'h3ad1;
10373: douta=16'h5394;
10374: douta=16'h6457;
10375: douta=16'h7c98;
10376: douta=16'h7478;
10377: douta=16'h63f5;
10378: douta=16'h63b3;
10379: douta=16'h5b92;
10380: douta=16'h9493;
10381: douta=16'h94f6;
10382: douta=16'h7bd2;
10383: douta=16'h9493;
10384: douta=16'h73f1;
10385: douta=16'hbd96;
10386: douta=16'hb596;
10387: douta=16'h8329;
10388: douta=16'h93ab;
10389: douta=16'h93cb;
10390: douta=16'hbcab;
10391: douta=16'hc50d;
10392: douta=16'hcd2e;
10393: douta=16'hd5b0;
10394: douta=16'hd5b0;
10395: douta=16'hddf3;
10396: douta=16'hde13;
10397: douta=16'heeb6;
10398: douta=16'heeb6;
10399: douta=16'hddf3;
10400: douta=16'he655;
10401: douta=16'hd5d2;
10402: douta=16'hbd10;
10403: douta=16'hc510;
10404: douta=16'ha44c;
10405: douta=16'h8b69;
10406: douta=16'ha44d;
10407: douta=16'hb4ee;
10408: douta=16'hc550;
10409: douta=16'hc570;
10410: douta=16'hddd1;
10411: douta=16'hddf3;
10412: douta=16'hde13;
10413: douta=16'hde13;
10414: douta=16'he634;
10415: douta=16'hde34;
10416: douta=16'hde14;
10417: douta=16'hd591;
10418: douta=16'hcd50;
10419: douta=16'hc511;
10420: douta=16'hb4d1;
10421: douta=16'ha491;
10422: douta=16'h9c72;
10423: douta=16'h8c32;
10424: douta=16'h8412;
10425: douta=16'h7bf2;
10426: douta=16'h6bb1;
10427: douta=16'h6391;
10428: douta=16'h6bb1;
10429: douta=16'h5b72;
10430: douta=16'h4acf;
10431: douta=16'h31a8;
10432: douta=16'h39ca;
10433: douta=16'h10e5;
10434: douta=16'h3a2b;
10435: douta=16'h1083;
10436: douta=16'h10a4;
10437: douta=16'h10e4;
10438: douta=16'h10c3;
10439: douta=16'h18c4;
10440: douta=16'h18e5;
10441: douta=16'h1905;
10442: douta=16'h10c4;
10443: douta=16'h08c5;
10444: douta=16'h4a8b;
10445: douta=16'h4aaa;
10446: douta=16'h5228;
10447: douta=16'h840e;
10448: douta=16'h840f;
10449: douta=16'hb4f1;
10450: douta=16'h83ac;
10451: douta=16'h5aca;
10452: douta=16'h18e4;
10453: douta=16'h736d;
10454: douta=16'h2967;
10455: douta=16'h630c;
10456: douta=16'h5a6a;
10457: douta=16'h63d2;
10458: douta=16'h9559;
10459: douta=16'h9539;
10460: douta=16'h84d7;
10461: douta=16'h7c96;
10462: douta=16'h8d18;
10463: douta=16'h84d8;
10464: douta=16'h6415;
10465: douta=16'h7476;
10466: douta=16'hae1c;
10467: douta=16'h9d9a;
10468: douta=16'h5372;
10469: douta=16'h7c75;
10470: douta=16'h8d18;
10471: douta=16'hbe5c;
10472: douta=16'hadfb;
10473: douta=16'ha5fa;
10474: douta=16'h957a;
10475: douta=16'h9dba;
10476: douta=16'h9d7a;
10477: douta=16'h9d9a;
10478: douta=16'h9dba;
10479: douta=16'ha5da;
10480: douta=16'h9d99;
10481: douta=16'hb63b;
10482: douta=16'hae1b;
10483: douta=16'h9579;
10484: douta=16'h9559;
10485: douta=16'h9d9a;
10486: douta=16'h8d18;
10487: douta=16'h8539;
10488: douta=16'h9579;
10489: douta=16'h8d18;
10490: douta=16'h94f7;
10491: douta=16'hb4d0;
10492: douta=16'h1105;
10493: douta=16'h1083;
10494: douta=16'h8519;
10495: douta=16'h84f8;
10496: douta=16'h957a;
10497: douta=16'h957a;
10498: douta=16'h84b8;
10499: douta=16'h84d7;
10500: douta=16'h9559;
10501: douta=16'h7c76;
10502: douta=16'h84d7;
10503: douta=16'ha5ba;
10504: douta=16'h9539;
10505: douta=16'h9558;
10506: douta=16'h8495;
10507: douta=16'h9517;
10508: douta=16'h9516;
10509: douta=16'h9518;
10510: douta=16'h9559;
10511: douta=16'h84d8;
10512: douta=16'h6c55;
10513: douta=16'h84f8;
10514: douta=16'h7cd8;
10515: douta=16'h8d9b;
10516: douta=16'h1906;
10517: douta=16'h08c4;
10518: douta=16'h2125;
10519: douta=16'h6478;
10520: douta=16'h5c37;
10521: douta=16'h74b9;
10522: douta=16'h6cb9;
10523: douta=16'h53f7;
10524: douta=16'h4353;
10525: douta=16'h74fa;
10526: douta=16'h855b;
10527: douta=16'h32f2;
10528: douta=16'h6cb9;
10529: douta=16'h5bd5;
10530: douta=16'h6c57;
10531: douta=16'h74d9;
10532: douta=16'h7cf9;
10533: douta=16'h74d9;
10534: douta=16'h8d5b;
10535: douta=16'h6c77;
10536: douta=16'h7cf9;
10537: douta=16'h7497;
10538: douta=16'h8d3a;
10539: douta=16'h7cf9;
10540: douta=16'h84f9;
10541: douta=16'h7498;
10542: douta=16'h8519;
10543: douta=16'h7cd9;
10544: douta=16'h7498;
10545: douta=16'h7cb8;
10546: douta=16'h7497;
10547: douta=16'h6c36;
10548: douta=16'h74b8;
10549: douta=16'h7cd9;
10550: douta=16'h6c77;
10551: douta=16'h63f3;
10552: douta=16'h6bf3;
10553: douta=16'ha5b9;
10554: douta=16'h6c34;
10555: douta=16'h7c33;
10556: douta=16'h63b1;
10557: douta=16'h8432;
10558: douta=16'h9d58;
10559: douta=16'h8c95;
10560: douta=16'h10c2;
10561: douta=16'h4354;
10562: douta=16'h2a6f;
10563: douta=16'h3b12;
10564: douta=16'h116b;
10565: douta=16'h226f;
10566: douta=16'h6436;
10567: douta=16'h7456;
10568: douta=16'h7d1a;
10569: douta=16'h74b9;
10570: douta=16'h63f4;
10571: douta=16'h5331;
10572: douta=16'h7413;
10573: douta=16'h9d16;
10574: douta=16'h7c13;
10575: douta=16'h9cd4;
10576: douta=16'h8411;
10577: douta=16'hb556;
10578: douta=16'h7b2b;
10579: douta=16'h93cb;
10580: douta=16'hac4b;
10581: douta=16'hac4b;
10582: douta=16'hcd6f;
10583: douta=16'hcd6f;
10584: douta=16'hd5b0;
10585: douta=16'hde34;
10586: douta=16'he655;
10587: douta=16'he674;
10588: douta=16'heeb6;
10589: douta=16'he634;
10590: douta=16'he675;
10591: douta=16'he634;
10592: douta=16'hcd92;
10593: douta=16'hd5d2;
10594: douta=16'ha42c;
10595: douta=16'ha42c;
10596: douta=16'h8b8a;
10597: douta=16'ha42c;
10598: douta=16'ha44d;
10599: douta=16'hac8d;
10600: douta=16'hd591;
10601: douta=16'hd5b1;
10602: douta=16'hddf2;
10603: douta=16'he654;
10604: douta=16'he654;
10605: douta=16'he654;
10606: douta=16'he654;
10607: douta=16'hddf3;
10608: douta=16'hddf3;
10609: douta=16'hc531;
10610: douta=16'hc531;
10611: douta=16'hbd11;
10612: douta=16'hacb0;
10613: douta=16'h8c31;
10614: douta=16'h9431;
10615: douta=16'h8c72;
10616: douta=16'h8c53;
10617: douta=16'h8c53;
10618: douta=16'h8c74;
10619: douta=16'h7c33;
10620: douta=16'ha556;
10621: douta=16'h69e3;
10622: douta=16'hb50f;
10623: douta=16'h3a0b;
10624: douta=16'h4209;
10625: douta=16'h2987;
10626: douta=16'h1906;
10627: douta=16'h2147;
10628: douta=16'h2147;
10629: douta=16'h0863;
10630: douta=16'h10a4;
10631: douta=16'h10c4;
10632: douta=16'h10a4;
10633: douta=16'h18e5;
10634: douta=16'h18c4;
10635: douta=16'h1906;
10636: douta=16'h08e5;
10637: douta=16'h84f7;
10638: douta=16'h4aac;
10639: douta=16'h6bce;
10640: douta=16'h08a3;
10641: douta=16'h8c0f;
10642: douta=16'h5aca;
10643: douta=16'h736c;
10644: douta=16'h5a8a;
10645: douta=16'h5269;
10646: douta=16'h39a6;
10647: douta=16'hbd92;
10648: douta=16'h9c70;
10649: douta=16'h6aca;
10650: douta=16'ha61c;
10651: douta=16'h9d7a;
10652: douta=16'h8d39;
10653: douta=16'h8d59;
10654: douta=16'h8d39;
10655: douta=16'h8d39;
10656: douta=16'h8d18;
10657: douta=16'h7c96;
10658: douta=16'h84f8;
10659: douta=16'h84d7;
10660: douta=16'h84f8;
10661: douta=16'h84d7;
10662: douta=16'h9579;
10663: douta=16'h8d39;
10664: douta=16'h9559;
10665: douta=16'h8518;
10666: douta=16'h6c15;
10667: douta=16'haddb;
10668: douta=16'hadfb;
10669: douta=16'hadda;
10670: douta=16'hb63b;
10671: douta=16'h9d9a;
10672: douta=16'h8d18;
10673: douta=16'h9579;
10674: douta=16'h9599;
10675: douta=16'h9599;
10676: douta=16'hadfa;
10677: douta=16'ha5ba;
10678: douta=16'ha5da;
10679: douta=16'h9d9a;
10680: douta=16'ha5ba;
10681: douta=16'h8518;
10682: douta=16'h9dba;
10683: douta=16'h9538;
10684: douta=16'h1083;
10685: douta=16'h0063;
10686: douta=16'h29e9;
10687: douta=16'h9538;
10688: douta=16'h8d39;
10689: douta=16'h6c35;
10690: douta=16'h8539;
10691: douta=16'h8d39;
10692: douta=16'h84f8;
10693: douta=16'h9d79;
10694: douta=16'h8496;
10695: douta=16'h84b6;
10696: douta=16'h7c55;
10697: douta=16'h8cb6;
10698: douta=16'h8496;
10699: douta=16'h8cd6;
10700: douta=16'h8cb6;
10701: douta=16'h9538;
10702: douta=16'h9dbb;
10703: douta=16'h9dbb;
10704: douta=16'h8d39;
10705: douta=16'h959b;
10706: douta=16'h8d9b;
10707: douta=16'h63d3;
10708: douta=16'h1083;
10709: douta=16'h2146;
10710: douta=16'h426c;
10711: douta=16'h7d1a;
10712: douta=16'h7d3b;
10713: douta=16'h7d1a;
10714: douta=16'h6c98;
10715: douta=16'h857b;
10716: douta=16'h857b;
10717: douta=16'h857b;
10718: douta=16'h9ddd;
10719: douta=16'h5c17;
10720: douta=16'h5c16;
10721: douta=16'h7d3b;
10722: douta=16'h74b9;
10723: douta=16'h6437;
10724: douta=16'h6437;
10725: douta=16'h74b8;
10726: douta=16'h7d1a;
10727: douta=16'h6c36;
10728: douta=16'h7477;
10729: douta=16'h7477;
10730: douta=16'h855a;
10731: douta=16'h959b;
10732: douta=16'h853a;
10733: douta=16'h7cfa;
10734: douta=16'h84f9;
10735: douta=16'h8d9b;
10736: douta=16'h851a;
10737: douta=16'h74b8;
10738: douta=16'h95dc;
10739: douta=16'h7cd8;
10740: douta=16'h6416;
10741: douta=16'h853a;
10742: douta=16'h41ea;
10743: douta=16'h52cd;
10744: douta=16'h6c13;
10745: douta=16'h6392;
10746: douta=16'h9d58;
10747: douta=16'h9d79;
10748: douta=16'h9559;
10749: douta=16'h0800;
10750: douta=16'h8474;
10751: douta=16'h8474;
10752: douta=16'h1082;
10753: douta=16'h53f7;
10754: douta=16'h21ed;
10755: douta=16'h2a4e;
10756: douta=16'h4354;
10757: douta=16'h32f2;
10758: douta=16'h74d9;
10759: douta=16'h7477;
10760: douta=16'h74b8;
10761: douta=16'h6c36;
10762: douta=16'h7435;
10763: douta=16'h8497;
10764: douta=16'h8cb6;
10765: douta=16'h9d16;
10766: douta=16'h5b30;
10767: douta=16'h6b90;
10768: douta=16'h8c72;
10769: douta=16'h8bcb;
10770: douta=16'h93ac;
10771: douta=16'ha42b;
10772: douta=16'hbcad;
10773: douta=16'hbccd;
10774: douta=16'hd5b1;
10775: douta=16'hcd6f;
10776: douta=16'hd5b0;
10777: douta=16'hee95;
10778: douta=16'hee96;
10779: douta=16'hee96;
10780: douta=16'hddf3;
10781: douta=16'heeb6;
10782: douta=16'he654;
10783: douta=16'hd5d1;
10784: douta=16'hc50e;
10785: douta=16'hbd0f;
10786: douta=16'h8349;
10787: douta=16'h8b8a;
10788: douta=16'h93eb;
10789: douta=16'hac4c;
10790: douta=16'hc54f;
10791: douta=16'hc54f;
10792: douta=16'hd5d2;
10793: douta=16'hde13;
10794: douta=16'he675;
10795: douta=16'he654;
10796: douta=16'hde14;
10797: douta=16'he634;
10798: douta=16'hde13;
10799: douta=16'he613;
10800: douta=16'hcd91;
10801: douta=16'hbd12;
10802: douta=16'hbcf1;
10803: douta=16'hb4d1;
10804: douta=16'hacb1;
10805: douta=16'h8c12;
10806: douta=16'h9452;
10807: douta=16'h8c53;
10808: douta=16'h8c33;
10809: douta=16'h6b70;
10810: douta=16'h8c73;
10811: douta=16'h5b2f;
10812: douta=16'h2947;
10813: douta=16'hd590;
10814: douta=16'h9c2e;
10815: douta=16'h422b;
10816: douta=16'h422a;
10817: douta=16'h31ea;
10818: douta=16'h2147;
10819: douta=16'h1927;
10820: douta=16'h1906;
10821: douta=16'h4a8c;
10822: douta=16'h1084;
10823: douta=16'h10e4;
10824: douta=16'h10c4;
10825: douta=16'h10e4;
10826: douta=16'h10e4;
10827: douta=16'h10c5;
10828: douta=16'h2187;
10829: douta=16'h0000;
10830: douta=16'h5371;
10831: douta=16'h3a4c;
10832: douta=16'h940d;
10833: douta=16'h630c;
10834: douta=16'h0883;
10835: douta=16'h0861;
10836: douta=16'h10c3;
10837: douta=16'h1905;
10838: douta=16'h8c0d;
10839: douta=16'h8c4e;
10840: douta=16'h39e8;
10841: douta=16'h8bef;
10842: douta=16'h6c13;
10843: douta=16'h8518;
10844: douta=16'h8d39;
10845: douta=16'h8d39;
10846: douta=16'h8d38;
10847: douta=16'h8d38;
10848: douta=16'h9579;
10849: douta=16'h8d18;
10850: douta=16'h7c96;
10851: douta=16'h7cb6;
10852: douta=16'h9558;
10853: douta=16'h9538;
10854: douta=16'h84d7;
10855: douta=16'h8d39;
10856: douta=16'h8d58;
10857: douta=16'h7476;
10858: douta=16'ha5db;
10859: douta=16'h9579;
10860: douta=16'h8518;
10861: douta=16'hadda;
10862: douta=16'ha5ba;
10863: douta=16'h8d59;
10864: douta=16'h959a;
10865: douta=16'h7cb7;
10866: douta=16'h8d38;
10867: douta=16'h9d99;
10868: douta=16'h959a;
10869: douta=16'h9579;
10870: douta=16'h9d9a;
10871: douta=16'ha5ba;
10872: douta=16'h9d99;
10873: douta=16'h9db9;
10874: douta=16'h9579;
10875: douta=16'h957a;
10876: douta=16'hc530;
10877: douta=16'h2926;
10878: douta=16'h1082;
10879: douta=16'h955a;
10880: douta=16'h9559;
10881: douta=16'h8d18;
10882: douta=16'h8d39;
10883: douta=16'h6c35;
10884: douta=16'h84b7;
10885: douta=16'h8cf7;
10886: douta=16'h84d7;
10887: douta=16'h7c75;
10888: douta=16'h9538;
10889: douta=16'h7c13;
10890: douta=16'h73f2;
10891: douta=16'h7c54;
10892: douta=16'h8cb6;
10893: douta=16'h84f8;
10894: douta=16'h7477;
10895: douta=16'h7497;
10896: douta=16'h84f9;
10897: douta=16'h851a;
10898: douta=16'h7476;
10899: douta=16'h2905;
10900: douta=16'h2167;
10901: douta=16'h31c8;
10902: douta=16'h5bf4;
10903: douta=16'h74b8;
10904: douta=16'h7d3a;
10905: douta=16'h74f9;
10906: douta=16'h6c78;
10907: douta=16'h6457;
10908: douta=16'h7d1a;
10909: douta=16'h8d7b;
10910: douta=16'h7cd9;
10911: douta=16'h9dfd;
10912: douta=16'h9dfd;
10913: douta=16'h7cd9;
10914: douta=16'h6417;
10915: douta=16'h6c98;
10916: douta=16'h74fa;
10917: douta=16'h5c37;
10918: douta=16'h7498;
10919: douta=16'h853a;
10920: douta=16'h7498;
10921: douta=16'h7cd9;
10922: douta=16'h6c36;
10923: douta=16'h74b8;
10924: douta=16'h7cf9;
10925: douta=16'h8d7a;
10926: douta=16'h8539;
10927: douta=16'h84d9;
10928: douta=16'h6c77;
10929: douta=16'h8d5b;
10930: douta=16'h84f9;
10931: douta=16'h7cb8;
10932: douta=16'h855a;
10933: douta=16'h6416;
10934: douta=16'h6391;
10935: douta=16'h8d3a;
10936: douta=16'h7c95;
10937: douta=16'h9d58;
10938: douta=16'h7454;
10939: douta=16'h7497;
10940: douta=16'h73f3;
10941: douta=16'h2167;
10942: douta=16'h9517;
10943: douta=16'h5351;
10944: douta=16'h1083;
10945: douta=16'h3ad0;
10946: douta=16'h2a90;
10947: douta=16'h3af2;
10948: douta=16'h32d1;
10949: douta=16'h2a70;
10950: douta=16'h6478;
10951: douta=16'h63d4;
10952: douta=16'h6416;
10953: douta=16'h7477;
10954: douta=16'h63b3;
10955: douta=16'h63f3;
10956: douta=16'h6bd2;
10957: douta=16'h94d6;
10958: douta=16'ha536;
10959: douta=16'had35;
10960: douta=16'h8c72;
10961: douta=16'h8b8a;
10962: douta=16'h8bab;
10963: douta=16'hac6b;
10964: douta=16'hb4ab;
10965: douta=16'hc50e;
10966: douta=16'hddd1;
10967: douta=16'hd5b0;
10968: douta=16'hd5b1;
10969: douta=16'hee96;
10970: douta=16'hee96;
10971: douta=16'hee96;
10972: douta=16'hcd4f;
10973: douta=16'hf6b6;
10974: douta=16'hee96;
10975: douta=16'hcd6f;
10976: douta=16'hcd30;
10977: douta=16'hb4cd;
10978: douta=16'h834a;
10979: douta=16'h9c2d;
10980: douta=16'ha42c;
10981: douta=16'hb48d;
10982: douta=16'hc54f;
10983: douta=16'hcd90;
10984: douta=16'hde13;
10985: douta=16'hde33;
10986: douta=16'he674;
10987: douta=16'he655;
10988: douta=16'he654;
10989: douta=16'he654;
10990: douta=16'hddf3;
10991: douta=16'hddf3;
10992: douta=16'hcd91;
10993: douta=16'hbcf1;
10994: douta=16'hb4d1;
10995: douta=16'hb4b2;
10996: douta=16'ha4b1;
10997: douta=16'h7bf2;
10998: douta=16'h9432;
10999: douta=16'h7bf2;
11000: douta=16'h7c12;
11001: douta=16'h6b70;
11002: douta=16'h6b70;
11003: douta=16'h5249;
11004: douta=16'h59e5;
11005: douta=16'hddd0;
11006: douta=16'h9c2e;
11007: douta=16'h524b;
11008: douta=16'h528b;
11009: douta=16'h3a2b;
11010: douta=16'h21a8;
11011: douta=16'h1105;
11012: douta=16'h10a4;
11013: douta=16'h1904;
11014: douta=16'h2987;
11015: douta=16'h10c4;
11016: douta=16'h10a4;
11017: douta=16'h10c4;
11018: douta=16'h10c4;
11019: douta=16'h10c5;
11020: douta=16'h1905;
11021: douta=16'h18e4;
11022: douta=16'h0000;
11023: douta=16'h5330;
11024: douta=16'h9cb4;
11025: douta=16'h528a;
11026: douta=16'h630b;
11027: douta=16'h9470;
11028: douta=16'h8c2e;
11029: douta=16'h2145;
11030: douta=16'h62aa;
11031: douta=16'h2124;
11032: douta=16'h7bad;
11033: douta=16'h738d;
11034: douta=16'h52ed;
11035: douta=16'h8d39;
11036: douta=16'h957a;
11037: douta=16'h8d39;
11038: douta=16'ha5db;
11039: douta=16'h8d59;
11040: douta=16'h9559;
11041: douta=16'h8d38;
11042: douta=16'h9579;
11043: douta=16'h8d38;
11044: douta=16'h8d18;
11045: douta=16'h8cf7;
11046: douta=16'h84d7;
11047: douta=16'h9559;
11048: douta=16'h9579;
11049: douta=16'h9559;
11050: douta=16'h84f8;
11051: douta=16'h8d59;
11052: douta=16'h957a;
11053: douta=16'h84f8;
11054: douta=16'h9d9a;
11055: douta=16'h9579;
11056: douta=16'h9d9a;
11057: douta=16'ha5da;
11058: douta=16'h9d99;
11059: douta=16'h9d99;
11060: douta=16'ha5da;
11061: douta=16'h9d79;
11062: douta=16'h9d9a;
11063: douta=16'h9d99;
11064: douta=16'h8d18;
11065: douta=16'ha5fa;
11066: douta=16'ha5da;
11067: douta=16'h9d9a;
11068: douta=16'hee73;
11069: douta=16'h9c0c;
11070: douta=16'h0882;
11071: douta=16'ha5db;
11072: douta=16'h8d17;
11073: douta=16'h84d8;
11074: douta=16'h8d39;
11075: douta=16'ha5ba;
11076: douta=16'h9d79;
11077: douta=16'h7c75;
11078: douta=16'h84d7;
11079: douta=16'h8495;
11080: douta=16'h8495;
11081: douta=16'h9d57;
11082: douta=16'h8cb5;
11083: douta=16'h94f6;
11084: douta=16'h7413;
11085: douta=16'h84f8;
11086: douta=16'h8519;
11087: douta=16'h7cd8;
11088: douta=16'h7498;
11089: douta=16'h8d7c;
11090: douta=16'h3a2b;
11091: douta=16'h2125;
11092: douta=16'h2188;
11093: douta=16'h2125;
11094: douta=16'h63f5;
11095: douta=16'h6c77;
11096: douta=16'h7cd8;
11097: douta=16'h853b;
11098: douta=16'h7d19;
11099: douta=16'h7d1a;
11100: douta=16'h74d9;
11101: douta=16'h8d9c;
11102: douta=16'h95bc;
11103: douta=16'h74b8;
11104: douta=16'ha63d;
11105: douta=16'h9dfd;
11106: douta=16'h95bc;
11107: douta=16'h853a;
11108: douta=16'h7d3a;
11109: douta=16'h6cb8;
11110: douta=16'h6c77;
11111: douta=16'h6436;
11112: douta=16'h851a;
11113: douta=16'h851a;
11114: douta=16'h7cb8;
11115: douta=16'h7498;
11116: douta=16'h6437;
11117: douta=16'h6c57;
11118: douta=16'h853a;
11119: douta=16'h8d5a;
11120: douta=16'h7cf9;
11121: douta=16'h7cd8;
11122: douta=16'h95bc;
11123: douta=16'h8d5a;
11124: douta=16'h7477;
11125: douta=16'h6350;
11126: douta=16'h9d9a;
11127: douta=16'h8d3a;
11128: douta=16'h63b2;
11129: douta=16'h5b93;
11130: douta=16'h7c55;
11131: douta=16'hbe5d;
11132: douta=16'h738f;
11133: douta=16'h5b50;
11134: douta=16'h8475;
11135: douta=16'h7413;
11136: douta=16'h2105;
11137: douta=16'h4334;
11138: douta=16'h32b1;
11139: douta=16'h3290;
11140: douta=16'h4354;
11141: douta=16'h2a90;
11142: douta=16'h4b53;
11143: douta=16'h63d4;
11144: douta=16'h7497;
11145: douta=16'h6c56;
11146: douta=16'h6372;
11147: douta=16'h7414;
11148: douta=16'h7414;
11149: douta=16'h7c33;
11150: douta=16'h73d2;
11151: douta=16'had77;
11152: douta=16'h9c0b;
11153: douta=16'h93eb;
11154: douta=16'h93ab;
11155: douta=16'hbcec;
11156: douta=16'hcd2e;
11157: douta=16'hd5b1;
11158: douta=16'hde12;
11159: douta=16'he654;
11160: douta=16'hddf2;
11161: douta=16'hee95;
11162: douta=16'heed7;
11163: douta=16'he675;
11164: douta=16'hddf3;
11165: douta=16'hddf3;
11166: douta=16'hcd70;
11167: douta=16'hc52f;
11168: douta=16'hac6c;
11169: douta=16'h93ca;
11170: douta=16'ha42c;
11171: douta=16'ha42c;
11172: douta=16'hb48d;
11173: douta=16'hd5d1;
11174: douta=16'hd5f2;
11175: douta=16'hddf3;
11176: douta=16'he674;
11177: douta=16'he634;
11178: douta=16'he675;
11179: douta=16'hee75;
11180: douta=16'he654;
11181: douta=16'he613;
11182: douta=16'hddd2;
11183: douta=16'hd591;
11184: douta=16'hc531;
11185: douta=16'hb4d1;
11186: douta=16'ha491;
11187: douta=16'h9452;
11188: douta=16'h9c92;
11189: douta=16'h6b91;
11190: douta=16'h4aad;
11191: douta=16'h8c32;
11192: douta=16'h7b8f;
11193: douta=16'h630e;
11194: douta=16'h8328;
11195: douta=16'hac6c;
11196: douta=16'ha42a;
11197: douta=16'hddd2;
11198: douta=16'ha44d;
11199: douta=16'h8bae;
11200: douta=16'h630d;
11201: douta=16'h630d;
11202: douta=16'h5aee;
11203: douta=16'h2167;
11204: douta=16'h2126;
11205: douta=16'h2126;
11206: douta=16'h10a4;
11207: douta=16'h2947;
11208: douta=16'h29a8;
11209: douta=16'h10a3;
11210: douta=16'h10c3;
11211: douta=16'h10a4;
11212: douta=16'h10c5;
11213: douta=16'h10c4;
11214: douta=16'h10a4;
11215: douta=16'h0042;
11216: douta=16'h1905;
11217: douta=16'h10e5;
11218: douta=16'h2146;
11219: douta=16'h83cd;
11220: douta=16'hd655;
11221: douta=16'ha490;
11222: douta=16'h6b0b;
11223: douta=16'h4a49;
11224: douta=16'h5acb;
11225: douta=16'h9c2e;
11226: douta=16'h62cb;
11227: douta=16'ha5fc;
11228: douta=16'h9559;
11229: douta=16'h9559;
11230: douta=16'h8518;
11231: douta=16'h957a;
11232: douta=16'h84f8;
11233: douta=16'h8d18;
11234: douta=16'h8d17;
11235: douta=16'h8d17;
11236: douta=16'h8d38;
11237: douta=16'h9538;
11238: douta=16'h84d7;
11239: douta=16'h8d18;
11240: douta=16'h84d7;
11241: douta=16'h8cf8;
11242: douta=16'h84d7;
11243: douta=16'h84d7;
11244: douta=16'h8d7a;
11245: douta=16'h84d8;
11246: douta=16'h74b7;
11247: douta=16'h8d5a;
11248: douta=16'h8d39;
11249: douta=16'h8d59;
11250: douta=16'h9dbb;
11251: douta=16'ha5da;
11252: douta=16'hadfb;
11253: douta=16'ha5ba;
11254: douta=16'h9d9a;
11255: douta=16'h959a;
11256: douta=16'h9d79;
11257: douta=16'h9579;
11258: douta=16'ha5da;
11259: douta=16'ha5ba;
11260: douta=16'hde13;
11261: douta=16'hff37;
11262: douta=16'hac0d;
11263: douta=16'h0001;
11264: douta=16'h2168;
11265: douta=16'hae1b;
11266: douta=16'h9d9a;
11267: douta=16'h9d9a;
11268: douta=16'h9d79;
11269: douta=16'h8cf6;
11270: douta=16'ha598;
11271: douta=16'h9537;
11272: douta=16'h8475;
11273: douta=16'h634f;
11274: douta=16'h73d2;
11275: douta=16'h7c95;
11276: douta=16'h7cb7;
11277: douta=16'h7cd8;
11278: douta=16'h7cf9;
11279: douta=16'h74d9;
11280: douta=16'h74b9;
11281: douta=16'h2146;
11282: douta=16'h18c3;
11283: douta=16'h21a8;
11284: douta=16'h0884;
11285: douta=16'h7cb8;
11286: douta=16'h6415;
11287: douta=16'h84b8;
11288: douta=16'h6c98;
11289: douta=16'h6c36;
11290: douta=16'h8d3a;
11291: douta=16'h8539;
11292: douta=16'h8d5a;
11293: douta=16'h8519;
11294: douta=16'h8519;
11295: douta=16'h7cd9;
11296: douta=16'h851a;
11297: douta=16'h8d5b;
11298: douta=16'h8d5a;
11299: douta=16'h8d5b;
11300: douta=16'h7d3a;
11301: douta=16'h7cf9;
11302: douta=16'h8d7b;
11303: douta=16'h853a;
11304: douta=16'h95bd;
11305: douta=16'h5bf6;
11306: douta=16'h7d19;
11307: douta=16'h7498;
11308: douta=16'h851a;
11309: douta=16'h74d9;
11310: douta=16'h8d5a;
11311: douta=16'h7cd9;
11312: douta=16'h6c57;
11313: douta=16'h7cd9;
11314: douta=16'h7cd8;
11315: douta=16'h6c37;
11316: douta=16'h74d9;
11317: douta=16'h5353;
11318: douta=16'ha5fc;
11319: douta=16'h9d79;
11320: douta=16'h4b31;
11321: douta=16'h63d2;
11322: douta=16'h84d7;
11323: douta=16'h49e9;
11324: douta=16'h1881;
11325: douta=16'h9517;
11326: douta=16'h6391;
11327: douta=16'h7c75;
11328: douta=16'h2905;
11329: douta=16'h29ea;
11330: douta=16'h2250;
11331: douta=16'h3ad1;
11332: douta=16'h32d2;
11333: douta=16'h32d1;
11334: douta=16'h53b5;
11335: douta=16'h5b93;
11336: douta=16'h5bb4;
11337: douta=16'h6c56;
11338: douta=16'h7c14;
11339: douta=16'h7435;
11340: douta=16'h7c76;
11341: douta=16'h9d17;
11342: douta=16'h94b5;
11343: douta=16'h734e;
11344: douta=16'h93aa;
11345: douta=16'ha42c;
11346: douta=16'hac4b;
11347: douta=16'hcd2e;
11348: douta=16'hd570;
11349: douta=16'hddd2;
11350: douta=16'he674;
11351: douta=16'heed7;
11352: douta=16'hf6f7;
11353: douta=16'he613;
11354: douta=16'hddd2;
11355: douta=16'he695;
11356: douta=16'hd5b1;
11357: douta=16'hc52f;
11358: douta=16'hcd90;
11359: douta=16'hbcce;
11360: douta=16'h8b69;
11361: douta=16'hac6d;
11362: douta=16'hac8d;
11363: douta=16'hb4ed;
11364: douta=16'hc50e;
11365: douta=16'hde13;
11366: douta=16'he655;
11367: douta=16'he654;
11368: douta=16'hee96;
11369: douta=16'heeb6;
11370: douta=16'hee75;
11371: douta=16'he634;
11372: douta=16'he654;
11373: douta=16'he654;
11374: douta=16'hd591;
11375: douta=16'hbd10;
11376: douta=16'hac91;
11377: douta=16'h9c52;
11378: douta=16'h9c72;
11379: douta=16'h9c92;
11380: douta=16'h8431;
11381: douta=16'h73d1;
11382: douta=16'h5aee;
11383: douta=16'h39ea;
11384: douta=16'h4a6b;
11385: douta=16'h5a26;
11386: douta=16'h93cb;
11387: douta=16'hcd2e;
11388: douta=16'he5f2;
11389: douta=16'hd58f;
11390: douta=16'hb48d;
11391: douta=16'h93ac;
11392: douta=16'h630d;
11393: douta=16'h630e;
11394: douta=16'h630e;
11395: douta=16'h3a4c;
11396: douta=16'h322c;
11397: douta=16'h322b;
11398: douta=16'h2988;
11399: douta=16'h1906;
11400: douta=16'h1084;
11401: douta=16'h0883;
11402: douta=16'h10a3;
11403: douta=16'h10c4;
11404: douta=16'h1905;
11405: douta=16'h10a4;
11406: douta=16'h10c5;
11407: douta=16'h2146;
11408: douta=16'h29a8;
11409: douta=16'h10c5;
11410: douta=16'h2126;
11411: douta=16'h1926;
11412: douta=16'h2167;
11413: douta=16'h8c6f;
11414: douta=16'h8c2e;
11415: douta=16'h1063;
11416: douta=16'h3986;
11417: douta=16'h31a6;
11418: douta=16'h6b0b;
11419: douta=16'h6391;
11420: douta=16'h7cb7;
11421: douta=16'h7496;
11422: douta=16'h9d7a;
11423: douta=16'h9559;
11424: douta=16'h9579;
11425: douta=16'h8d38;
11426: douta=16'h8d38;
11427: douta=16'h9579;
11428: douta=16'h8d38;
11429: douta=16'h8d18;
11430: douta=16'h84f8;
11431: douta=16'h9d99;
11432: douta=16'h8d58;
11433: douta=16'h8d18;
11434: douta=16'h8d18;
11435: douta=16'h9559;
11436: douta=16'h84d8;
11437: douta=16'h8d18;
11438: douta=16'h9559;
11439: douta=16'h9d9a;
11440: douta=16'h8d39;
11441: douta=16'h8518;
11442: douta=16'h8d18;
11443: douta=16'h957a;
11444: douta=16'h9d9a;
11445: douta=16'h9559;
11446: douta=16'h8d39;
11447: douta=16'h8d39;
11448: douta=16'h9d9a;
11449: douta=16'h9d9a;
11450: douta=16'h9d9a;
11451: douta=16'h9d79;
11452: douta=16'h8d5a;
11453: douta=16'had34;
11454: douta=16'hff98;
11455: douta=16'h29eb;
11456: douta=16'h1106;
11457: douta=16'h0043;
11458: douta=16'ha5fb;
11459: douta=16'h9d79;
11460: douta=16'h9538;
11461: douta=16'h9d58;
11462: douta=16'h9d58;
11463: douta=16'h8c94;
11464: douta=16'h8473;
11465: douta=16'h9d16;
11466: douta=16'h9537;
11467: douta=16'h73f4;
11468: douta=16'h6cb8;
11469: douta=16'h53f5;
11470: douta=16'h753c;
11471: douta=16'h7d5c;
11472: douta=16'h39ea;
11473: douta=16'h20e5;
11474: douta=16'h322c;
11475: douta=16'h1927;
11476: douta=16'h7d1a;
11477: douta=16'h7d3a;
11478: douta=16'h853a;
11479: douta=16'h853a;
11480: douta=16'h8d5a;
11481: douta=16'h84f9;
11482: douta=16'h6c36;
11483: douta=16'h7498;
11484: douta=16'h853a;
11485: douta=16'h853a;
11486: douta=16'h853a;
11487: douta=16'h8519;
11488: douta=16'h8519;
11489: douta=16'h8d5a;
11490: douta=16'h8d7b;
11491: douta=16'h851a;
11492: douta=16'h855a;
11493: douta=16'h8d7b;
11494: douta=16'h853a;
11495: douta=16'h853b;
11496: douta=16'h853a;
11497: douta=16'h7cfa;
11498: douta=16'h855a;
11499: douta=16'h5394;
11500: douta=16'h8d7b;
11501: douta=16'h7cd9;
11502: douta=16'h959b;
11503: douta=16'h8d5a;
11504: douta=16'h7498;
11505: douta=16'h74d8;
11506: douta=16'h74d8;
11507: douta=16'h6cda;
11508: douta=16'h72cb;
11509: douta=16'ha5fb;
11510: douta=16'h7414;
11511: douta=16'h5351;
11512: douta=16'h7c76;
11513: douta=16'h7cb7;
11514: douta=16'h84f8;
11515: douta=16'h0800;
11516: douta=16'h5330;
11517: douta=16'h6c14;
11518: douta=16'h7454;
11519: douta=16'h7c95;
11520: douta=16'h2925;
11521: douta=16'h29a9;
11522: douta=16'h4bd6;
11523: douta=16'h222e;
11524: douta=16'h3312;
11525: douta=16'h220d;
11526: douta=16'h3ad1;
11527: douta=16'h5b94;
11528: douta=16'h7cb8;
11529: douta=16'h7498;
11530: douta=16'h324c;
11531: douta=16'h5b92;
11532: douta=16'h6c14;
11533: douta=16'h8c94;
11534: douta=16'h94d4;
11535: douta=16'h62a9;
11536: douta=16'h93cb;
11537: douta=16'hac4b;
11538: douta=16'hb48b;
11539: douta=16'hcd4f;
11540: douta=16'hd590;
11541: douta=16'hddf2;
11542: douta=16'hee96;
11543: douta=16'heeb6;
11544: douta=16'heeb6;
11545: douta=16'he695;
11546: douta=16'hde13;
11547: douta=16'he634;
11548: douta=16'hd570;
11549: douta=16'hcd4f;
11550: douta=16'hc52e;
11551: douta=16'h938a;
11552: douta=16'hb48d;
11553: douta=16'ha44c;
11554: douta=16'hbcee;
11555: douta=16'hbced;
11556: douta=16'hd591;
11557: douta=16'he634;
11558: douta=16'he675;
11559: douta=16'he675;
11560: douta=16'hee96;
11561: douta=16'hee96;
11562: douta=16'he654;
11563: douta=16'he613;
11564: douta=16'hde13;
11565: douta=16'he613;
11566: douta=16'hd592;
11567: douta=16'hbcef;
11568: douta=16'h9c51;
11569: douta=16'h9c71;
11570: douta=16'h9c72;
11571: douta=16'h9452;
11572: douta=16'h8432;
11573: douta=16'h7bf2;
11574: douta=16'h6b6f;
11575: douta=16'h2988;
11576: douta=16'h20e6;
11577: douta=16'h82e7;
11578: douta=16'hac6c;
11579: douta=16'hddb1;
11580: douta=16'he654;
11581: douta=16'hddd1;
11582: douta=16'hbcac;
11583: douta=16'h9bed;
11584: douta=16'h632d;
11585: douta=16'h5b0d;
11586: douta=16'h6b6f;
11587: douta=16'h5310;
11588: douta=16'h42af;
11589: douta=16'h42ae;
11590: douta=16'h29cb;
11591: douta=16'h2168;
11592: douta=16'h10c4;
11593: douta=16'h428d;
11594: douta=16'h10a4;
11595: douta=16'h18e5;
11596: douta=16'h10e5;
11597: douta=16'h10a4;
11598: douta=16'h10a4;
11599: douta=16'h10a3;
11600: douta=16'h1905;
11601: douta=16'h10e5;
11602: douta=16'h1926;
11603: douta=16'h1926;
11604: douta=16'h08c5;
11605: douta=16'h52aa;
11606: douta=16'hc5d4;
11607: douta=16'ha4d2;
11608: douta=16'h9c2f;
11609: douta=16'h630b;
11610: douta=16'h20c3;
11611: douta=16'h3988;
11612: douta=16'h9dbb;
11613: douta=16'h84d7;
11614: douta=16'h9559;
11615: douta=16'h9d9a;
11616: douta=16'h9dba;
11617: douta=16'h9dba;
11618: douta=16'h84f7;
11619: douta=16'h8d39;
11620: douta=16'h84f8;
11621: douta=16'h84f8;
11622: douta=16'h84f8;
11623: douta=16'h8d38;
11624: douta=16'h8d39;
11625: douta=16'h9d7a;
11626: douta=16'h8d39;
11627: douta=16'h84f8;
11628: douta=16'h8539;
11629: douta=16'h8d18;
11630: douta=16'h7cb7;
11631: douta=16'h8d39;
11632: douta=16'h8d39;
11633: douta=16'h957a;
11634: douta=16'h9559;
11635: douta=16'h84d7;
11636: douta=16'h8d38;
11637: douta=16'h9dba;
11638: douta=16'h84f8;
11639: douta=16'h8517;
11640: douta=16'h8d39;
11641: douta=16'ha5da;
11642: douta=16'h957a;
11643: douta=16'h8d39;
11644: douta=16'h9dbb;
11645: douta=16'h8519;
11646: douta=16'hf6b4;
11647: douta=16'h426d;
11648: douta=16'h4b0f;
11649: douta=16'h0001;
11650: douta=16'h3aae;
11651: douta=16'h9dbb;
11652: douta=16'ha5fb;
11653: douta=16'h9d79;
11654: douta=16'h9517;
11655: douta=16'ha557;
11656: douta=16'h8c93;
11657: douta=16'h8493;
11658: douta=16'h7c74;
11659: douta=16'h7d3a;
11660: douta=16'h5c37;
11661: douta=16'h5c58;
11662: douta=16'h4b94;
11663: douta=16'h322c;
11664: douta=16'h2904;
11665: douta=16'h3a8d;
11666: douta=16'h2189;
11667: douta=16'h4311;
11668: douta=16'h7cfa;
11669: douta=16'h5c15;
11670: douta=16'h7d19;
11671: douta=16'h95bb;
11672: douta=16'h8d7a;
11673: douta=16'h959b;
11674: douta=16'h8d1a;
11675: douta=16'h53b4;
11676: douta=16'h7497;
11677: douta=16'h8d5a;
11678: douta=16'h959c;
11679: douta=16'h853a;
11680: douta=16'h7498;
11681: douta=16'h7498;
11682: douta=16'h84f9;
11683: douta=16'h8d7b;
11684: douta=16'h959c;
11685: douta=16'h8d7c;
11686: douta=16'h8d7b;
11687: douta=16'h7cf9;
11688: douta=16'h853a;
11689: douta=16'h853a;
11690: douta=16'h95bc;
11691: douta=16'h6457;
11692: douta=16'h7498;
11693: douta=16'h8d5b;
11694: douta=16'h74b8;
11695: douta=16'h6c78;
11696: douta=16'h7d3a;
11697: douta=16'h7cf9;
11698: douta=16'h53d6;
11699: douta=16'h3af1;
11700: douta=16'h736f;
11701: douta=16'h5330;
11702: douta=16'h9d9a;
11703: douta=16'h8cf8;
11704: douta=16'h8d18;
11705: douta=16'h63f4;
11706: douta=16'h63d4;
11707: douta=16'h2946;
11708: douta=16'h7cd8;
11709: douta=16'hadfa;
11710: douta=16'h5b72;
11711: douta=16'h6c13;
11712: douta=16'h3146;
11713: douta=16'h2126;
11714: douta=16'h3ad1;
11715: douta=16'h2a90;
11716: douta=16'h53f7;
11717: douta=16'h4374;
11718: douta=16'h32f1;
11719: douta=16'h326f;
11720: douta=16'h7c98;
11721: douta=16'h6c57;
11722: douta=16'h4acf;
11723: douta=16'h5b72;
11724: douta=16'h6bd3;
11725: douta=16'h9d37;
11726: douta=16'h8b8b;
11727: douta=16'h93aa;
11728: douta=16'hac6b;
11729: douta=16'hbc8b;
11730: douta=16'hd56f;
11731: douta=16'hd5b0;
11732: douta=16'hddd1;
11733: douta=16'hee95;
11734: douta=16'hee95;
11735: douta=16'hee96;
11736: douta=16'heeb6;
11737: douta=16'he674;
11738: douta=16'he654;
11739: douta=16'hcd70;
11740: douta=16'hc4cf;
11741: douta=16'hb48d;
11742: douta=16'h8b69;
11743: douta=16'h9bea;
11744: douta=16'hac6c;
11745: douta=16'hb4ad;
11746: douta=16'hcd6f;
11747: douta=16'hd5b0;
11748: douta=16'hddf3;
11749: douta=16'he655;
11750: douta=16'he675;
11751: douta=16'he675;
11752: douta=16'he674;
11753: douta=16'he654;
11754: douta=16'he654;
11755: douta=16'hddf2;
11756: douta=16'hdd92;
11757: douta=16'hcd70;
11758: douta=16'hbcef;
11759: douta=16'h9c30;
11760: douta=16'h9451;
11761: douta=16'h7bd1;
11762: douta=16'h7bf2;
11763: douta=16'h734e;
11764: douta=16'h7b8f;
11765: douta=16'h6b4f;
11766: douta=16'h630e;
11767: douta=16'h7b08;
11768: douta=16'h938a;
11769: douta=16'ha42c;
11770: douta=16'hd590;
11771: douta=16'he634;
11772: douta=16'he613;
11773: douta=16'hdd8f;
11774: douta=16'hcd0e;
11775: douta=16'ha42d;
11776: douta=16'h838e;
11777: douta=16'h732e;
11778: douta=16'h634e;
11779: douta=16'h6350;
11780: douta=16'h4aef;
11781: douta=16'h5b51;
11782: douta=16'h42cf;
11783: douta=16'h324d;
11784: douta=16'h29ec;
11785: douta=16'h2168;
11786: douta=16'h0884;
11787: douta=16'h5b0e;
11788: douta=16'h10c4;
11789: douta=16'h18e4;
11790: douta=16'h10e5;
11791: douta=16'h10c4;
11792: douta=16'h10c5;
11793: douta=16'h10a3;
11794: douta=16'h2146;
11795: douta=16'h10e4;
11796: douta=16'h18e5;
11797: douta=16'h6bb1;
11798: douta=16'h2966;
11799: douta=16'hd678;
11800: douta=16'h840e;
11801: douta=16'h2946;
11802: douta=16'h528a;
11803: douta=16'h0002;
11804: douta=16'h41c7;
11805: douta=16'h5b70;
11806: douta=16'h84f8;
11807: douta=16'h84f7;
11808: douta=16'h8d39;
11809: douta=16'h7c96;
11810: douta=16'h8d39;
11811: douta=16'h957a;
11812: douta=16'ha5fb;
11813: douta=16'h9d7a;
11814: douta=16'h84d7;
11815: douta=16'h84f8;
11816: douta=16'h84f8;
11817: douta=16'h9559;
11818: douta=16'h84d7;
11819: douta=16'h84d7;
11820: douta=16'h7496;
11821: douta=16'h84f8;
11822: douta=16'h7c96;
11823: douta=16'h7cb6;
11824: douta=16'h84f8;
11825: douta=16'h7c96;
11826: douta=16'h84d7;
11827: douta=16'h84d7;
11828: douta=16'h9d9a;
11829: douta=16'h8d38;
11830: douta=16'h9559;
11831: douta=16'h9559;
11832: douta=16'h8d39;
11833: douta=16'h9579;
11834: douta=16'h9d9a;
11835: douta=16'h9d9a;
11836: douta=16'h84f8;
11837: douta=16'h9559;
11838: douta=16'ha5db;
11839: douta=16'h7b4c;
11840: douta=16'h7b6e;
11841: douta=16'h7476;
11842: douta=16'h322d;
11843: douta=16'h1906;
11844: douta=16'h18c4;
11845: douta=16'h21eb;
11846: douta=16'h63d3;
11847: douta=16'h7bce;
11848: douta=16'h0882;
11849: douta=16'h1968;
11850: douta=16'h4c39;
11851: douta=16'h2a2c;
11852: douta=16'h1082;
11853: douta=16'h3145;
11854: douta=16'h5a6a;
11855: douta=16'h49a7;
11856: douta=16'h6c98;
11857: douta=16'h29a9;
11858: douta=16'h324c;
11859: douta=16'h7cf9;
11860: douta=16'h7cd8;
11861: douta=16'h84f9;
11862: douta=16'h7c98;
11863: douta=16'h7cd9;
11864: douta=16'h8d5a;
11865: douta=16'h957b;
11866: douta=16'h959b;
11867: douta=16'h9dbc;
11868: douta=16'h9dbc;
11869: douta=16'h8d7a;
11870: douta=16'h9ddc;
11871: douta=16'h8d3a;
11872: douta=16'h6436;
11873: douta=16'h7497;
11874: douta=16'h7cd8;
11875: douta=16'h8d3a;
11876: douta=16'h957b;
11877: douta=16'h8d7b;
11878: douta=16'h74b8;
11879: douta=16'h6415;
11880: douta=16'h6c56;
11881: douta=16'h9ddc;
11882: douta=16'h8d5a;
11883: douta=16'h8d5b;
11884: douta=16'h851a;
11885: douta=16'h74d9;
11886: douta=16'h853a;
11887: douta=16'h6437;
11888: douta=16'h5bd5;
11889: douta=16'h4b53;
11890: douta=16'h7b8e;
11891: douta=16'h6b90;
11892: douta=16'h3880;
11893: douta=16'h4b72;
11894: douta=16'h9559;
11895: douta=16'hadb9;
11896: douta=16'h53b4;
11897: douta=16'h7456;
11898: douta=16'h5350;
11899: douta=16'h9559;
11900: douta=16'ha599;
11901: douta=16'h9d98;
11902: douta=16'h1084;
11903: douta=16'h0000;
11904: douta=16'h2945;
11905: douta=16'h18e4;
11906: douta=16'h328f;
11907: douta=16'h3290;
11908: douta=16'h4bb5;
11909: douta=16'h4374;
11910: douta=16'h2a2e;
11911: douta=16'h5bf5;
11912: douta=16'h84d8;
11913: douta=16'h7456;
11914: douta=16'h5b72;
11915: douta=16'h5b51;
11916: douta=16'h7434;
11917: douta=16'ha599;
11918: douta=16'h9bca;
11919: douta=16'hac4c;
11920: douta=16'hb4ad;
11921: douta=16'hc4ed;
11922: douta=16'hd5af;
11923: douta=16'he613;
11924: douta=16'he633;
11925: douta=16'heeb6;
11926: douta=16'hee75;
11927: douta=16'heeb6;
11928: douta=16'he674;
11929: douta=16'hd5b2;
11930: douta=16'hd5b1;
11931: douta=16'hcd70;
11932: douta=16'hac6c;
11933: douta=16'h8308;
11934: douta=16'ha40b;
11935: douta=16'h9beb;
11936: douta=16'hbccd;
11937: douta=16'hc50e;
11938: douta=16'hcd90;
11939: douta=16'hde12;
11940: douta=16'he675;
11941: douta=16'hee96;
11942: douta=16'hee95;
11943: douta=16'he675;
11944: douta=16'he674;
11945: douta=16'he613;
11946: douta=16'hddd2;
11947: douta=16'hd591;
11948: douta=16'hc530;
11949: douta=16'hc510;
11950: douta=16'h9c50;
11951: douta=16'h9431;
11952: douta=16'h9431;
11953: douta=16'h6aed;
11954: douta=16'h630e;
11955: douta=16'h736f;
11956: douta=16'h6b0e;
11957: douta=16'h49e8;
11958: douta=16'h4185;
11959: douta=16'h9c0c;
11960: douta=16'h9bcb;
11961: douta=16'hc52f;
11962: douta=16'he5f2;
11963: douta=16'he654;
11964: douta=16'he654;
11965: douta=16'hd58f;
11966: douta=16'hc4ee;
11967: douta=16'ha42d;
11968: douta=16'h838d;
11969: douta=16'h7b4d;
11970: douta=16'h632e;
11971: douta=16'h634f;
11972: douta=16'h6b71;
11973: douta=16'h5b50;
11974: douta=16'h52f0;
11975: douta=16'h3a8e;
11976: douta=16'h320c;
11977: douta=16'h2189;
11978: douta=16'h2168;
11979: douta=16'h0884;
11980: douta=16'h10a4;
11981: douta=16'h10e4;
11982: douta=16'h18c4;
11983: douta=16'h10c4;
11984: douta=16'h10a4;
11985: douta=16'h10c4;
11986: douta=16'h18e4;
11987: douta=16'h1905;
11988: douta=16'h1906;
11989: douta=16'h6b90;
11990: douta=16'h6b90;
11991: douta=16'h52ed;
11992: douta=16'h4228;
11993: douta=16'h5269;
11994: douta=16'h62cb;
11995: douta=16'h8c0f;
11996: douta=16'h6b2b;
11997: douta=16'h5269;
11998: douta=16'h84f8;
11999: douta=16'h8d38;
12000: douta=16'h7cb6;
12001: douta=16'h8d18;
12002: douta=16'h84b7;
12003: douta=16'h8d59;
12004: douta=16'h84f8;
12005: douta=16'h8d39;
12006: douta=16'h9579;
12007: douta=16'ha5ba;
12008: douta=16'h9558;
12009: douta=16'h7476;
12010: douta=16'h8d18;
12011: douta=16'h7496;
12012: douta=16'h7cb7;
12013: douta=16'h7c96;
12014: douta=16'h84d7;
12015: douta=16'h8d38;
12016: douta=16'h9579;
12017: douta=16'h8d39;
12018: douta=16'h84f8;
12019: douta=16'h84f7;
12020: douta=16'h8d18;
12021: douta=16'h9559;
12022: douta=16'h84f8;
12023: douta=16'h8d18;
12024: douta=16'h9559;
12025: douta=16'h9559;
12026: douta=16'h84f8;
12027: douta=16'h8d18;
12028: douta=16'ha5db;
12029: douta=16'h9559;
12030: douta=16'h7496;
12031: douta=16'ha5fc;
12032: douta=16'h9db9;
12033: douta=16'h6330;
12034: douta=16'h4a8d;
12035: douta=16'h1989;
12036: douta=16'h1968;
12037: douta=16'h1948;
12038: douta=16'h10e5;
12039: douta=16'h0064;
12040: douta=16'h2146;
12041: douta=16'h1905;
12042: douta=16'h1061;
12043: douta=16'h4a08;
12044: douta=16'h834c;
12045: douta=16'h8b4b;
12046: douta=16'h6c14;
12047: douta=16'h63f4;
12048: douta=16'h5350;
12049: douta=16'h7c97;
12050: douta=16'h853b;
12051: douta=16'h8519;
12052: douta=16'h6c78;
12053: douta=16'h6c37;
12054: douta=16'h959c;
12055: douta=16'h74b8;
12056: douta=16'h7cb8;
12057: douta=16'h7c98;
12058: douta=16'h8d3a;
12059: douta=16'h8d5a;
12060: douta=16'ha61c;
12061: douta=16'h851a;
12062: douta=16'h8d5b;
12063: douta=16'h95bb;
12064: douta=16'h95dc;
12065: douta=16'h95bc;
12066: douta=16'h95bc;
12067: douta=16'h7d19;
12068: douta=16'h74b8;
12069: douta=16'h7477;
12070: douta=16'h959c;
12071: douta=16'h8d7b;
12072: douta=16'h95bb;
12073: douta=16'h6c16;
12074: douta=16'h5bf5;
12075: douta=16'h74b8;
12076: douta=16'h7cf9;
12077: douta=16'h851a;
12078: douta=16'h7cd9;
12079: douta=16'h7d1a;
12080: douta=16'h857b;
12081: douta=16'h857c;
12082: douta=16'h7c98;
12083: douta=16'h63d4;
12084: douta=16'h4374;
12085: douta=16'h72a6;
12086: douta=16'h3965;
12087: douta=16'h2a4d;
12088: douta=16'h7499;
12089: douta=16'h6c56;
12090: douta=16'h4165;
12091: douta=16'ha5db;
12092: douta=16'h84b6;
12093: douta=16'h63d5;
12094: douta=16'h2125;
12095: douta=16'h1083;
12096: douta=16'h3166;
12097: douta=16'h1083;
12098: douta=16'h328e;
12099: douta=16'h4b94;
12100: douta=16'h4353;
12101: douta=16'h3af2;
12102: douta=16'h4353;
12103: douta=16'h5bf5;
12104: douta=16'h84d8;
12105: douta=16'h7457;
12106: douta=16'h5b52;
12107: douta=16'h6bb3;
12108: douta=16'h84b6;
12109: douta=16'h73f3;
12110: douta=16'hac4b;
12111: douta=16'hb4ac;
12112: douta=16'hbcad;
12113: douta=16'hc50e;
12114: douta=16'hd5d0;
12115: douta=16'he634;
12116: douta=16'he654;
12117: douta=16'hee96;
12118: douta=16'he675;
12119: douta=16'he633;
12120: douta=16'hee95;
12121: douta=16'hd591;
12122: douta=16'hd590;
12123: douta=16'hcd4f;
12124: douta=16'h93aa;
12125: douta=16'h9bcb;
12126: douta=16'hac6c;
12127: douta=16'ha44c;
12128: douta=16'hbcee;
12129: douta=16'hc50e;
12130: douta=16'hd5b1;
12131: douta=16'hde13;
12132: douta=16'he675;
12133: douta=16'hee96;
12134: douta=16'hee75;
12135: douta=16'hee75;
12136: douta=16'hee75;
12137: douta=16'he632;
12138: douta=16'hddb2;
12139: douta=16'hcd71;
12140: douta=16'hc4f0;
12141: douta=16'hbcd0;
12142: douta=16'h9c50;
12143: douta=16'h8c11;
12144: douta=16'h83f1;
12145: douta=16'h62cd;
12146: douta=16'h62cd;
12147: douta=16'h5acc;
12148: douta=16'h5aab;
12149: douta=16'h4164;
12150: douta=16'h7ac7;
12151: douta=16'hb48e;
12152: douta=16'hbcae;
12153: douta=16'hd5b1;
12154: douta=16'he634;
12155: douta=16'hee55;
12156: douta=16'he633;
12157: douta=16'hd58f;
12158: douta=16'hbcad;
12159: douta=16'ha42d;
12160: douta=16'ha42e;
12161: douta=16'h838d;
12162: douta=16'h734f;
12163: douta=16'h634f;
12164: douta=16'h6b71;
12165: douta=16'h6371;
12166: douta=16'h4af0;
12167: douta=16'h42ae;
12168: douta=16'h322c;
12169: douta=16'h29ea;
12170: douta=16'h21a9;
12171: douta=16'h2128;
12172: douta=16'h4a8d;
12173: douta=16'h10a3;
12174: douta=16'h10e5;
12175: douta=16'h10a3;
12176: douta=16'h18e4;
12177: douta=16'h10a4;
12178: douta=16'h10a3;
12179: douta=16'h10c5;
12180: douta=16'h18e5;
12181: douta=16'h18e5;
12182: douta=16'h7433;
12183: douta=16'h5b50;
12184: douta=16'h6b2c;
12185: douta=16'h8bce;
12186: douta=16'h8bcd;
12187: douta=16'h8c30;
12188: douta=16'h734d;
12189: douta=16'ha4f1;
12190: douta=16'h8d7a;
12191: douta=16'h7cb6;
12192: douta=16'h7c96;
12193: douta=16'h7475;
12194: douta=16'h84d7;
12195: douta=16'h6c14;
12196: douta=16'h8d38;
12197: douta=16'h8cf8;
12198: douta=16'h7c96;
12199: douta=16'h9d9a;
12200: douta=16'ha5db;
12201: douta=16'ha599;
12202: douta=16'h84f8;
12203: douta=16'h84f8;
12204: douta=16'h7c97;
12205: douta=16'h8d38;
12206: douta=16'h84f8;
12207: douta=16'h84b7;
12208: douta=16'h8d17;
12209: douta=16'h8d18;
12210: douta=16'h8d18;
12211: douta=16'h8cd8;
12212: douta=16'h84d7;
12213: douta=16'h8d39;
12214: douta=16'h9559;
12215: douta=16'h8d18;
12216: douta=16'h8d18;
12217: douta=16'h9dba;
12218: douta=16'h9559;
12219: douta=16'h8d59;
12220: douta=16'h8d18;
12221: douta=16'h959a;
12222: douta=16'h957a;
12223: douta=16'h7c97;
12224: douta=16'h957b;
12225: douta=16'h8495;
12226: douta=16'h424b;
12227: douta=16'h4aae;
12228: douta=16'h3a6d;
12229: douta=16'h21a9;
12230: douta=16'h21a9;
12231: douta=16'h1947;
12232: douta=16'h0882;
12233: douta=16'h2125;
12234: douta=16'h49e8;
12235: douta=16'ha40e;
12236: douta=16'h936c;
12237: douta=16'h7bf2;
12238: douta=16'h5350;
12239: douta=16'h3a0a;
12240: douta=16'h4a8d;
12241: douta=16'ha61d;
12242: douta=16'h8d19;
12243: douta=16'h8d3a;
12244: douta=16'h9539;
12245: douta=16'h7c77;
12246: douta=16'h5394;
12247: douta=16'h957b;
12248: douta=16'h7cb8;
12249: douta=16'h74b8;
12250: douta=16'h7c98;
12251: douta=16'h851a;
12252: douta=16'h8d5b;
12253: douta=16'ha63d;
12254: douta=16'h8d7a;
12255: douta=16'h8d5a;
12256: douta=16'h8d5b;
12257: douta=16'h851a;
12258: douta=16'h8d9b;
12259: douta=16'h853a;
12260: douta=16'h7c98;
12261: douta=16'h7cd8;
12262: douta=16'h6415;
12263: douta=16'h95bc;
12264: douta=16'h853a;
12265: douta=16'h95bc;
12266: douta=16'h6c57;
12267: douta=16'h6c77;
12268: douta=16'h7cd9;
12269: douta=16'h74b8;
12270: douta=16'h6c77;
12271: douta=16'h74b8;
12272: douta=16'h751b;
12273: douta=16'h7d3a;
12274: douta=16'h63f5;
12275: douta=16'h9d9a;
12276: douta=16'h63f4;
12277: douta=16'h959a;
12278: douta=16'h6249;
12279: douta=16'h40e1;
12280: douta=16'h53b5;
12281: douta=16'h7d5c;
12282: douta=16'h1000;
12283: douta=16'h9559;
12284: douta=16'hbe7b;
12285: douta=16'h7455;
12286: douta=16'h2967;
12287: douta=16'h1083;
12288: douta=16'h39a7;
12289: douta=16'h18a4;
12290: douta=16'h322b;
12291: douta=16'h3b12;
12292: douta=16'h3b13;
12293: douta=16'h53f6;
12294: douta=16'h2a4f;
12295: douta=16'h6c36;
12296: douta=16'h7cb7;
12297: douta=16'h7476;
12298: douta=16'h5b52;
12299: douta=16'h6b92;
12300: douta=16'h84b6;
12301: douta=16'h7bf2;
12302: douta=16'hbcad;
12303: douta=16'hbced;
12304: douta=16'hcd4f;
12305: douta=16'hd590;
12306: douta=16'hde13;
12307: douta=16'hee75;
12308: douta=16'he654;
12309: douta=16'hee95;
12310: douta=16'he653;
12311: douta=16'hddf2;
12312: douta=16'hc50d;
12313: douta=16'hd590;
12314: douta=16'hc4ee;
12315: douta=16'h9bea;
12316: douta=16'hac4c;
12317: douta=16'hac6d;
12318: douta=16'hb4ad;
12319: douta=16'hac6c;
12320: douta=16'hcd8f;
12321: douta=16'hcd90;
12322: douta=16'hde33;
12323: douta=16'hee75;
12324: douta=16'he695;
12325: douta=16'hee96;
12326: douta=16'hee95;
12327: douta=16'he675;
12328: douta=16'he613;
12329: douta=16'hde33;
12330: douta=16'hd5d2;
12331: douta=16'ha46f;
12332: douta=16'ha450;
12333: douta=16'h9c50;
12334: douta=16'h83d0;
12335: douta=16'h83f0;
12336: douta=16'h6b0d;
12337: douta=16'h630c;
12338: douta=16'h630c;
12339: douta=16'h41e8;
12340: douta=16'h8b48;
12341: douta=16'h9c0b;
12342: douta=16'h9c0c;
12343: douta=16'hd5b1;
12344: douta=16'hde13;
12345: douta=16'hee95;
12346: douta=16'hee75;
12347: douta=16'hde13;
12348: douta=16'hddd1;
12349: douta=16'hcd0e;
12350: douta=16'hc4cd;
12351: douta=16'ha42d;
12352: douta=16'h9c0e;
12353: douta=16'h93ce;
12354: douta=16'h8bcf;
12355: douta=16'h7bb0;
12356: douta=16'h6b91;
12357: douta=16'h6bb1;
12358: douta=16'h6392;
12359: douta=16'h4b10;
12360: douta=16'h42ae;
12361: douta=16'h322c;
12362: douta=16'h324d;
12363: douta=16'h2a0b;
12364: douta=16'h2189;
12365: douta=16'h3a4b;
12366: douta=16'h5b0f;
12367: douta=16'h18e4;
12368: douta=16'h10c4;
12369: douta=16'h10a3;
12370: douta=16'h10c4;
12371: douta=16'h10c5;
12372: douta=16'h18e5;
12373: douta=16'h1926;
12374: douta=16'h18e5;
12375: douta=16'h2988;
12376: douta=16'h5b50;
12377: douta=16'h4b2f;
12378: douta=16'h0842;
12379: douta=16'h9cb0;
12380: douta=16'h83ee;
12381: douta=16'h5aaa;
12382: douta=16'h7b8c;
12383: douta=16'h31ea;
12384: douta=16'h9559;
12385: douta=16'h6c34;
12386: douta=16'h7c96;
12387: douta=16'h7cb7;
12388: douta=16'h9559;
12389: douta=16'h84f8;
12390: douta=16'h84f8;
12391: douta=16'h84f8;
12392: douta=16'h84d7;
12393: douta=16'h84d7;
12394: douta=16'h9559;
12395: douta=16'h6c14;
12396: douta=16'h6c14;
12397: douta=16'ha5db;
12398: douta=16'h9dba;
12399: douta=16'h9559;
12400: douta=16'h9579;
12401: douta=16'h9559;
12402: douta=16'h9d9a;
12403: douta=16'h9558;
12404: douta=16'h9d7a;
12405: douta=16'h84f7;
12406: douta=16'h9559;
12407: douta=16'h8518;
12408: douta=16'h8d18;
12409: douta=16'h9559;
12410: douta=16'h9dbb;
12411: douta=16'h9559;
12412: douta=16'h84f8;
12413: douta=16'h957a;
12414: douta=16'h9559;
12415: douta=16'h957a;
12416: douta=16'h8d59;
12417: douta=16'h9559;
12418: douta=16'h9579;
12419: douta=16'h8d18;
12420: douta=16'h7cb6;
12421: douta=16'h528c;
12422: douta=16'h4aad;
12423: douta=16'h5c56;
12424: douta=16'h32ae;
12425: douta=16'h6414;
12426: douta=16'h6c76;
12427: douta=16'h3a09;
12428: douta=16'h5aef;
12429: douta=16'h9d9a;
12430: douta=16'h8d7a;
12431: douta=16'h8539;
12432: douta=16'h8d59;
12433: douta=16'h957a;
12434: douta=16'h957a;
12435: douta=16'h8d39;
12436: douta=16'h9dbb;
12437: douta=16'h8d7a;
12438: douta=16'h8d5a;
12439: douta=16'ha61c;
12440: douta=16'h8539;
12441: douta=16'h8518;
12442: douta=16'h7cb8;
12443: douta=16'h7cd9;
12444: douta=16'h8519;
12445: douta=16'h8d7b;
12446: douta=16'h84d9;
12447: douta=16'h853a;
12448: douta=16'h74b8;
12449: douta=16'h7cf9;
12450: douta=16'h959b;
12451: douta=16'h95bb;
12452: douta=16'h957b;
12453: douta=16'h851a;
12454: douta=16'h8d5a;
12455: douta=16'h95bb;
12456: douta=16'h959c;
12457: douta=16'h7cb8;
12458: douta=16'h7498;
12459: douta=16'h7cd9;
12460: douta=16'h7d1a;
12461: douta=16'h7cd9;
12462: douta=16'h7cd9;
12463: douta=16'h7414;
12464: douta=16'h6c55;
12465: douta=16'h7d3b;
12466: douta=16'h4b11;
12467: douta=16'h63f5;
12468: douta=16'h95bc;
12469: douta=16'h63f5;
12470: douta=16'h5bf5;
12471: douta=16'h7477;
12472: douta=16'h851a;
12473: douta=16'h838d;
12474: douta=16'h0000;
12475: douta=16'h2290;
12476: douta=16'h43b5;
12477: douta=16'h74b7;
12478: douta=16'h8433;
12479: douta=16'h10a3;
12480: douta=16'h3986;
12481: douta=16'h18e3;
12482: douta=16'h31ca;
12483: douta=16'h4bb5;
12484: douta=16'h4374;
12485: douta=16'h4bb5;
12486: douta=16'h3ad1;
12487: douta=16'h6415;
12488: douta=16'h63d4;
12489: douta=16'h7477;
12490: douta=16'h5b72;
12491: douta=16'h6392;
12492: douta=16'h84b6;
12493: douta=16'h7bf2;
12494: douta=16'hc4ed;
12495: douta=16'hbced;
12496: douta=16'hcd8f;
12497: douta=16'hde13;
12498: douta=16'hee75;
12499: douta=16'heeb6;
12500: douta=16'hee95;
12501: douta=16'he654;
12502: douta=16'he633;
12503: douta=16'hd5b0;
12504: douta=16'hd570;
12505: douta=16'hac4c;
12506: douta=16'hbcee;
12507: douta=16'h8348;
12508: douta=16'hb48d;
12509: douta=16'hb4cd;
12510: douta=16'hbccd;
12511: douta=16'hc4ee;
12512: douta=16'hde33;
12513: douta=16'hd5b0;
12514: douta=16'he654;
12515: douta=16'he675;
12516: douta=16'hee95;
12517: douta=16'heeb6;
12518: douta=16'hee75;
12519: douta=16'he654;
12520: douta=16'hddd1;
12521: douta=16'hd590;
12522: douta=16'hd570;
12523: douta=16'h9c30;
12524: douta=16'h83d0;
12525: douta=16'h8c10;
12526: douta=16'h6b2e;
12527: douta=16'h734f;
12528: douta=16'h732e;
12529: douta=16'h4a29;
12530: douta=16'h2925;
12531: douta=16'h9308;
12532: douta=16'hac2b;
12533: douta=16'hcd2f;
12534: douta=16'hd56f;
12535: douta=16'hee75;
12536: douta=16'hee95;
12537: douta=16'heeb6;
12538: douta=16'hee75;
12539: douta=16'hee54;
12540: douta=16'hddf2;
12541: douta=16'hcd0f;
12542: douta=16'hc4cf;
12543: douta=16'hb46e;
12544: douta=16'h9bee;
12545: douta=16'h93ce;
12546: douta=16'h93ef;
12547: douta=16'h8410;
12548: douta=16'h7bf2;
12549: douta=16'h7bf2;
12550: douta=16'h63b2;
12551: douta=16'h5b91;
12552: douta=16'h4b10;
12553: douta=16'h320c;
12554: douta=16'h29cb;
12555: douta=16'h29aa;
12556: douta=16'h2a0c;
12557: douta=16'h31eb;
12558: douta=16'h2146;
12559: douta=16'h3a0b;
12560: douta=16'h1905;
12561: douta=16'h1926;
12562: douta=16'h18e5;
12563: douta=16'h2147;
12564: douta=16'h1926;
12565: douta=16'h18e5;
12566: douta=16'h18e5;
12567: douta=16'h18e5;
12568: douta=16'h31ea;
12569: douta=16'h10e4;
12570: douta=16'h18e5;
12571: douta=16'h630c;
12572: douta=16'h6b6d;
12573: douta=16'h526a;
12574: douta=16'h8c2f;
12575: douta=16'h8bed;
12576: douta=16'h29a9;
12577: douta=16'h84f7;
12578: douta=16'h7cb7;
12579: douta=16'h84b7;
12580: douta=16'h8d38;
12581: douta=16'h84f8;
12582: douta=16'h84d7;
12583: douta=16'h7c96;
12584: douta=16'h63f4;
12585: douta=16'h8d18;
12586: douta=16'h84f8;
12587: douta=16'h8d38;
12588: douta=16'h84d7;
12589: douta=16'h84f7;
12590: douta=16'h8d18;
12591: douta=16'h9559;
12592: douta=16'ha5fb;
12593: douta=16'hbe7c;
12594: douta=16'hae1b;
12595: douta=16'ha5ba;
12596: douta=16'h8d39;
12597: douta=16'h8d59;
12598: douta=16'h9559;
12599: douta=16'h9559;
12600: douta=16'ha5fb;
12601: douta=16'h8d18;
12602: douta=16'h8d39;
12603: douta=16'h84f8;
12604: douta=16'h957a;
12605: douta=16'h8d18;
12606: douta=16'h7456;
12607: douta=16'h8d18;
12608: douta=16'h957a;
12609: douta=16'h957a;
12610: douta=16'h8d18;
12611: douta=16'h9d9a;
12612: douta=16'h9ddb;
12613: douta=16'h8539;
12614: douta=16'h853a;
12615: douta=16'h734f;
12616: douta=16'h4a4b;
12617: douta=16'h2188;
12618: douta=16'h2906;
12619: douta=16'h9ddc;
12620: douta=16'h8d59;
12621: douta=16'h8518;
12622: douta=16'h959a;
12623: douta=16'h959a;
12624: douta=16'ha5db;
12625: douta=16'h9d9a;
12626: douta=16'h8539;
12627: douta=16'h74b8;
12628: douta=16'h8519;
12629: douta=16'h7cf8;
12630: douta=16'h8d59;
12631: douta=16'h8519;
12632: douta=16'h9dbb;
12633: douta=16'h959a;
12634: douta=16'h9ddb;
12635: douta=16'h959a;
12636: douta=16'h8519;
12637: douta=16'h853a;
12638: douta=16'h8d3a;
12639: douta=16'h7d19;
12640: douta=16'h8d5b;
12641: douta=16'h855a;
12642: douta=16'h8d3a;
12643: douta=16'h8d1a;
12644: douta=16'h7498;
12645: douta=16'h95bb;
12646: douta=16'h957b;
12647: douta=16'h853a;
12648: douta=16'h8d9b;
12649: douta=16'h853a;
12650: douta=16'h95bc;
12651: douta=16'h8d7b;
12652: douta=16'h6c56;
12653: douta=16'h74b8;
12654: douta=16'h6c98;
12655: douta=16'h84d8;
12656: douta=16'h32ae;
12657: douta=16'h5372;
12658: douta=16'h8d18;
12659: douta=16'hae1c;
12660: douta=16'h6416;
12661: douta=16'h5bd4;
12662: douta=16'h4b33;
12663: douta=16'h5372;
12664: douta=16'h9ddc;
12665: douta=16'h0000;
12666: douta=16'hb71f;
12667: douta=16'h6b0a;
12668: douta=16'h61e4;
12669: douta=16'h2947;
12670: douta=16'h7c96;
12671: douta=16'h0882;
12672: douta=16'h3166;
12673: douta=16'h18e4;
12674: douta=16'h31c9;
12675: douta=16'h4374;
12676: douta=16'h3290;
12677: douta=16'h5c16;
12678: douta=16'h2a50;
12679: douta=16'h5bf5;
12680: douta=16'h6c36;
12681: douta=16'h6c36;
12682: douta=16'h5b92;
12683: douta=16'h6392;
12684: douta=16'h7414;
12685: douta=16'h73d1;
12686: douta=16'hc4ed;
12687: douta=16'hc50e;
12688: douta=16'hcd8f;
12689: douta=16'he613;
12690: douta=16'hee95;
12691: douta=16'hf6b6;
12692: douta=16'hf6d7;
12693: douta=16'he654;
12694: douta=16'hddf2;
12695: douta=16'hd56f;
12696: douta=16'hcd2f;
12697: douta=16'h9baa;
12698: douta=16'h7ae7;
12699: douta=16'hb48d;
12700: douta=16'hbd2e;
12701: douta=16'hbd0d;
12702: douta=16'hbcee;
12703: douta=16'hcd6f;
12704: douta=16'he655;
12705: douta=16'hd5b0;
12706: douta=16'heeb6;
12707: douta=16'hee75;
12708: douta=16'heeb6;
12709: douta=16'hee96;
12710: douta=16'hee95;
12711: douta=16'he654;
12712: douta=16'hddb2;
12713: douta=16'hcd50;
12714: douta=16'hcd30;
12715: douta=16'h8bd0;
12716: douta=16'h7bb0;
12717: douta=16'h7bd0;
12718: douta=16'h6b2f;
12719: douta=16'h6b2d;
12720: douta=16'h7b8f;
12721: douta=16'h28e3;
12722: douta=16'h51a5;
12723: douta=16'h9be9;
12724: douta=16'hc4ee;
12725: douta=16'hd5b1;
12726: douta=16'hddf2;
12727: douta=16'hee96;
12728: douta=16'heeb6;
12729: douta=16'hee95;
12730: douta=16'he634;
12731: douta=16'he634;
12732: douta=16'hddf2;
12733: douta=16'hcd0f;
12734: douta=16'hbcae;
12735: douta=16'hac4e;
12736: douta=16'ha42e;
12737: douta=16'ha42f;
12738: douta=16'h8c10;
12739: douta=16'h8c11;
12740: douta=16'h8412;
12741: douta=16'h8433;
12742: douta=16'h7414;
12743: douta=16'h63b2;
12744: douta=16'h5b51;
12745: douta=16'h428e;
12746: douta=16'h3a8d;
12747: douta=16'h3a6d;
12748: douta=16'h3af0;
12749: douta=16'h31c9;
12750: douta=16'h31c9;
12751: douta=16'h42ae;
12752: douta=16'h5310;
12753: douta=16'h1927;
12754: douta=16'h18e5;
12755: douta=16'h1906;
12756: douta=16'h1926;
12757: douta=16'h1925;
12758: douta=16'h18e5;
12759: douta=16'h1905;
12760: douta=16'h10c5;
12761: douta=16'h18e5;
12762: douta=16'h10e5;
12763: douta=16'h0001;
12764: douta=16'h2987;
12765: douta=16'h7b6e;
12766: douta=16'h5acb;
12767: douta=16'h9c70;
12768: douta=16'h4a28;
12769: douta=16'hae3d;
12770: douta=16'h7c96;
12771: douta=16'h7455;
12772: douta=16'h9579;
12773: douta=16'h9d9a;
12774: douta=16'h84f8;
12775: douta=16'h7c96;
12776: douta=16'h7455;
12777: douta=16'h7c76;
12778: douta=16'h8d18;
12779: douta=16'h9559;
12780: douta=16'h9579;
12781: douta=16'h84d7;
12782: douta=16'h84d7;
12783: douta=16'h84b6;
12784: douta=16'h9539;
12785: douta=16'hadda;
12786: douta=16'hb63b;
12787: douta=16'h8d18;
12788: douta=16'h8d39;
12789: douta=16'h9559;
12790: douta=16'h957a;
12791: douta=16'h8d39;
12792: douta=16'h7cb7;
12793: douta=16'h8d59;
12794: douta=16'h9559;
12795: douta=16'h955a;
12796: douta=16'h8518;
12797: douta=16'h8d59;
12798: douta=16'h84f8;
12799: douta=16'h6c55;
12800: douta=16'h6c15;
12801: douta=16'h84f9;
12802: douta=16'h8d39;
12803: douta=16'h8d59;
12804: douta=16'h84f8;
12805: douta=16'h957a;
12806: douta=16'h8d5a;
12807: douta=16'h8432;
12808: douta=16'h4a6b;
12809: douta=16'h1041;
12810: douta=16'h39e9;
12811: douta=16'h8519;
12812: douta=16'h959a;
12813: douta=16'h9d9a;
12814: douta=16'h957a;
12815: douta=16'h957a;
12816: douta=16'h957a;
12817: douta=16'h959a;
12818: douta=16'h9dbb;
12819: douta=16'h8d59;
12820: douta=16'h9dbb;
12821: douta=16'h957a;
12822: douta=16'h957a;
12823: douta=16'h9ddb;
12824: douta=16'h8d7a;
12825: douta=16'h9dbb;
12826: douta=16'h959b;
12827: douta=16'h959a;
12828: douta=16'ha61c;
12829: douta=16'h7cf9;
12830: douta=16'h8519;
12831: douta=16'h7cf9;
12832: douta=16'h957a;
12833: douta=16'h853a;
12834: douta=16'h7cd9;
12835: douta=16'h8d5a;
12836: douta=16'h7cd8;
12837: douta=16'h7cd9;
12838: douta=16'h8d3a;
12839: douta=16'h9e1d;
12840: douta=16'h9e1e;
12841: douta=16'h853a;
12842: douta=16'h8d5b;
12843: douta=16'h8d7b;
12844: douta=16'h8d7b;
12845: douta=16'h7d7c;
12846: douta=16'h6b2c;
12847: douta=16'h9dfd;
12848: douta=16'h74b9;
12849: douta=16'h74b9;
12850: douta=16'h7cb7;
12851: douta=16'h6c57;
12852: douta=16'h5bd4;
12853: douta=16'h9dbb;
12854: douta=16'h6c35;
12855: douta=16'h9d7a;
12856: douta=16'h5394;
12857: douta=16'h1860;
12858: douta=16'h8d5a;
12859: douta=16'h95bb;
12860: douta=16'h84b6;
12861: douta=16'h7225;
12862: douta=16'h3a4c;
12863: douta=16'h1883;
12864: douta=16'h3986;
12865: douta=16'h2925;
12866: douta=16'h31a8;
12867: douta=16'h2a6f;
12868: douta=16'h2a4e;
12869: douta=16'h3b12;
12870: douta=16'h32b0;
12871: douta=16'h6436;
12872: douta=16'h5352;
12873: douta=16'h7455;
12874: douta=16'h6393;
12875: douta=16'h5b72;
12876: douta=16'h7434;
12877: douta=16'h7c13;
12878: douta=16'hcd2e;
12879: douta=16'hcd6f;
12880: douta=16'hddf2;
12881: douta=16'hee75;
12882: douta=16'heeb6;
12883: douta=16'hee75;
12884: douta=16'he654;
12885: douta=16'hee95;
12886: douta=16'hac6d;
12887: douta=16'hb46e;
12888: douta=16'hb48d;
12889: douta=16'ha42c;
12890: douta=16'hb4ad;
12891: douta=16'haccd;
12892: douta=16'hc52e;
12893: douta=16'hde13;
12894: douta=16'hc54f;
12895: douta=16'he676;
12896: douta=16'hee96;
12897: douta=16'he654;
12898: douta=16'hee96;
12899: douta=16'hee96;
12900: douta=16'he633;
12901: douta=16'he675;
12902: douta=16'he613;
12903: douta=16'he633;
12904: douta=16'hb4af;
12905: douta=16'hb48f;
12906: douta=16'hac8f;
12907: douta=16'h83cf;
12908: douta=16'h734f;
12909: douta=16'h732e;
12910: douta=16'h62ec;
12911: douta=16'h5aab;
12912: douta=16'h20c4;
12913: douta=16'hb46c;
12914: douta=16'hac4c;
12915: douta=16'hbccc;
12916: douta=16'he612;
12917: douta=16'he654;
12918: douta=16'hee75;
12919: douta=16'heeb6;
12920: douta=16'heeb6;
12921: douta=16'he655;
12922: douta=16'he613;
12923: douta=16'hddd2;
12924: douta=16'hddb2;
12925: douta=16'hbccf;
12926: douta=16'hbcaf;
12927: douta=16'hac6e;
12928: douta=16'h8bef;
12929: douta=16'h9410;
12930: douta=16'h9451;
12931: douta=16'h9452;
12932: douta=16'h9473;
12933: douta=16'h8c53;
12934: douta=16'h8454;
12935: douta=16'h7c54;
12936: douta=16'h7414;
12937: douta=16'h6bd2;
12938: douta=16'h6bf2;
12939: douta=16'h4b32;
12940: douta=16'hb46f;
12941: douta=16'h42ae;
12942: douta=16'h322b;
12943: douta=16'h31ea;
12944: douta=16'h1906;
12945: douta=16'h2988;
12946: douta=16'h0863;
12947: douta=16'h0883;
12948: douta=16'h10a3;
12949: douta=16'h10c3;
12950: douta=16'h10a4;
12951: douta=16'h10c4;
12952: douta=16'h18e5;
12953: douta=16'h1905;
12954: douta=16'h10c4;
12955: douta=16'h10a3;
12956: douta=16'h18e5;
12957: douta=16'h1905;
12958: douta=16'hbd72;
12959: douta=16'h8430;
12960: douta=16'h9491;
12961: douta=16'hd635;
12962: douta=16'h31eb;
12963: douta=16'h7cb7;
12964: douta=16'h8d38;
12965: douta=16'h8d18;
12966: douta=16'h9d9a;
12967: douta=16'h84f8;
12968: douta=16'h7cb7;
12969: douta=16'h9d7a;
12970: douta=16'h8d38;
12971: douta=16'h9579;
12972: douta=16'h9559;
12973: douta=16'h7434;
12974: douta=16'h63d3;
12975: douta=16'h84d7;
12976: douta=16'h8d18;
12977: douta=16'h7c96;
12978: douta=16'h7c97;
12979: douta=16'h6c15;
12980: douta=16'h6c35;
12981: douta=16'h8518;
12982: douta=16'h9559;
12983: douta=16'h959a;
12984: douta=16'h959a;
12985: douta=16'h7cb7;
12986: douta=16'h8518;
12987: douta=16'h8518;
12988: douta=16'h7cb7;
12989: douta=16'h7cd8;
12990: douta=16'h8518;
12991: douta=16'h955a;
12992: douta=16'h8d39;
12993: douta=16'h8539;
12994: douta=16'h957a;
12995: douta=16'h7cd7;
12996: douta=16'h7cd8;
12997: douta=16'h959a;
12998: douta=16'h8d59;
12999: douta=16'h9473;
13000: douta=16'h4a6c;
13001: douta=16'h1062;
13002: douta=16'h39e9;
13003: douta=16'h8519;
13004: douta=16'h8d59;
13005: douta=16'h7cf8;
13006: douta=16'h9ddb;
13007: douta=16'h959a;
13008: douta=16'h9dbb;
13009: douta=16'hae3c;
13010: douta=16'h8539;
13011: douta=16'h8539;
13012: douta=16'h8539;
13013: douta=16'h959a;
13014: douta=16'h8d39;
13015: douta=16'h959b;
13016: douta=16'h9ddb;
13017: douta=16'h7cf9;
13018: douta=16'ha5fb;
13019: douta=16'h959b;
13020: douta=16'h8d5a;
13021: douta=16'ha61c;
13022: douta=16'ha5fb;
13023: douta=16'h8539;
13024: douta=16'ha5fc;
13025: douta=16'h7497;
13026: douta=16'h7497;
13027: douta=16'h9dbb;
13028: douta=16'h957b;
13029: douta=16'h95bb;
13030: douta=16'h8d3a;
13031: douta=16'h8519;
13032: douta=16'h7cd9;
13033: douta=16'h7cd8;
13034: douta=16'h853a;
13035: douta=16'h7d3a;
13036: douta=16'h524a;
13037: douta=16'h0000;
13038: douta=16'h2127;
13039: douta=16'h4921;
13040: douta=16'h74fa;
13041: douta=16'h95dc;
13042: douta=16'h53b4;
13043: douta=16'h53b4;
13044: douta=16'h9dbc;
13045: douta=16'h9dbb;
13046: douta=16'h8d39;
13047: douta=16'h8518;
13048: douta=16'h5184;
13049: douta=16'h53f5;
13050: douta=16'h7477;
13051: douta=16'hcefe;
13052: douta=16'h8d19;
13053: douta=16'h8d39;
13054: douta=16'h6cba;
13055: douta=16'h3964;
13056: douta=16'h3966;
13057: douta=16'h3145;
13058: douta=16'h1083;
13059: douta=16'h32d1;
13060: douta=16'h32b1;
13061: douta=16'h32b1;
13062: douta=16'h4353;
13063: douta=16'h5394;
13064: douta=16'h7456;
13065: douta=16'h7cb7;
13066: douta=16'h63f5;
13067: douta=16'h6372;
13068: douta=16'h7c55;
13069: douta=16'h6bd2;
13070: douta=16'hbcef;
13071: douta=16'hd58e;
13072: douta=16'he654;
13073: douta=16'hee76;
13074: douta=16'heeb6;
13075: douta=16'he634;
13076: douta=16'he613;
13077: douta=16'hd570;
13078: douta=16'hcd70;
13079: douta=16'h7b07;
13080: douta=16'h51c4;
13081: douta=16'hb4ad;
13082: douta=16'hbcee;
13083: douta=16'hd5b1;
13084: douta=16'hd5b1;
13085: douta=16'hd5d3;
13086: douta=16'hc570;
13087: douta=16'heeb6;
13088: douta=16'hddf3;
13089: douta=16'hf6f8;
13090: douta=16'he675;
13091: douta=16'hee95;
13092: douta=16'he654;
13093: douta=16'he613;
13094: douta=16'hde12;
13095: douta=16'hd5b1;
13096: douta=16'hb4ae;
13097: douta=16'ha46f;
13098: douta=16'h83af;
13099: douta=16'h7b8f;
13100: douta=16'h6b2c;
13101: douta=16'h62ec;
13102: douta=16'h5a6a;
13103: douta=16'h3145;
13104: douta=16'ha388;
13105: douta=16'hb46b;
13106: douta=16'hc4cc;
13107: douta=16'hddd1;
13108: douta=16'he634;
13109: douta=16'hde33;
13110: douta=16'he654;
13111: douta=16'heeb6;
13112: douta=16'heeb6;
13113: douta=16'he654;
13114: douta=16'he613;
13115: douta=16'hd572;
13116: douta=16'hcd71;
13117: douta=16'hbcb0;
13118: douta=16'hac50;
13119: douta=16'h9c30;
13120: douta=16'h9451;
13121: douta=16'h8c31;
13122: douta=16'h8c11;
13123: douta=16'h8c32;
13124: douta=16'h8412;
13125: douta=16'h8412;
13126: douta=16'h73b1;
13127: douta=16'h736f;
13128: douta=16'h632e;
13129: douta=16'h62ac;
13130: douta=16'h6a8a;
13131: douta=16'hd52b;
13132: douta=16'ha48f;
13133: douta=16'h4ace;
13134: douta=16'h29eb;
13135: douta=16'h3a8c;
13136: douta=16'h2147;
13137: douta=16'h1905;
13138: douta=16'h2947;
13139: douta=16'h5b0e;
13140: douta=16'h39ea;
13141: douta=16'h10c5;
13142: douta=16'h10e5;
13143: douta=16'h18e5;
13144: douta=16'h18e5;
13145: douta=16'h18c4;
13146: douta=16'h2106;
13147: douta=16'h18e5;
13148: douta=16'h0883;
13149: douta=16'h0863;
13150: douta=16'h8453;
13151: douta=16'h9492;
13152: douta=16'ha4b2;
13153: douta=16'h7c0f;
13154: douta=16'h634d;
13155: douta=16'h39e8;
13156: douta=16'h8d18;
13157: douta=16'h8d18;
13158: douta=16'h84d7;
13159: douta=16'h8d38;
13160: douta=16'h9579;
13161: douta=16'h8d18;
13162: douta=16'h8d38;
13163: douta=16'h9579;
13164: douta=16'h9579;
13165: douta=16'h84b6;
13166: douta=16'h8d18;
13167: douta=16'h8d39;
13168: douta=16'h6c35;
13169: douta=16'h84d7;
13170: douta=16'h8d18;
13171: douta=16'h8518;
13172: douta=16'h7c96;
13173: douta=16'h84f8;
13174: douta=16'h7435;
13175: douta=16'h5352;
13176: douta=16'h7496;
13177: douta=16'h84f8;
13178: douta=16'h9dbb;
13179: douta=16'h8d59;
13180: douta=16'h84f8;
13181: douta=16'h8518;
13182: douta=16'h959a;
13183: douta=16'h84f8;
13184: douta=16'h8539;
13185: douta=16'h8d5a;
13186: douta=16'h8d59;
13187: douta=16'h7cf8;
13188: douta=16'h8518;
13189: douta=16'h7cb7;
13190: douta=16'h8518;
13191: douta=16'h8c52;
13192: douta=16'h528c;
13193: douta=16'h18a2;
13194: douta=16'h31c9;
13195: douta=16'h8d59;
13196: douta=16'h8538;
13197: douta=16'h9ddb;
13198: douta=16'h8539;
13199: douta=16'h8518;
13200: douta=16'h7cd8;
13201: douta=16'h959b;
13202: douta=16'h9ddb;
13203: douta=16'h959a;
13204: douta=16'h9ddb;
13205: douta=16'h95ba;
13206: douta=16'ha5db;
13207: douta=16'h8519;
13208: douta=16'h8d9a;
13209: douta=16'h8d7a;
13210: douta=16'h8d59;
13211: douta=16'ha5db;
13212: douta=16'ha5fb;
13213: douta=16'h8d5a;
13214: douta=16'h957a;
13215: douta=16'h9d9b;
13216: douta=16'h8519;
13217: douta=16'h7cd9;
13218: douta=16'h8d3a;
13219: douta=16'h84f9;
13220: douta=16'h7497;
13221: douta=16'h7cb8;
13222: douta=16'h853a;
13223: douta=16'h957b;
13224: douta=16'h95bb;
13225: douta=16'h851a;
13226: douta=16'h84f9;
13227: douta=16'h62cb;
13228: douta=16'h2903;
13229: douta=16'h10a2;
13230: douta=16'h0020;
13231: douta=16'h8d39;
13232: douta=16'h4060;
13233: douta=16'h29ec;
13234: douta=16'h5bf5;
13235: douta=16'h84f9;
13236: douta=16'h7cd7;
13237: douta=16'h6c56;
13238: douta=16'h42f1;
13239: douta=16'h3af1;
13240: douta=16'h0800;
13241: douta=16'h8d7a;
13242: douta=16'h9dba;
13243: douta=16'h7c76;
13244: douta=16'h8497;
13245: douta=16'h6436;
13246: douta=16'h6c15;
13247: douta=16'h0020;
13248: douta=16'h3966;
13249: douta=16'h3165;
13250: douta=16'h1063;
13251: douta=16'h4333;
13252: douta=16'h2a2e;
13253: douta=16'h3270;
13254: douta=16'h2a8f;
13255: douta=16'h4332;
13256: douta=16'h6c36;
13257: douta=16'h7456;
13258: douta=16'h7456;
13259: douta=16'h6bb3;
13260: douta=16'h7c55;
13261: douta=16'h7413;
13262: douta=16'h9c52;
13263: douta=16'hddb0;
13264: douta=16'he654;
13265: douta=16'hee96;
13266: douta=16'hee95;
13267: douta=16'hde33;
13268: douta=16'hddf2;
13269: douta=16'hcd6f;
13270: douta=16'hbcee;
13271: douta=16'h7b28;
13272: douta=16'h72c7;
13273: douta=16'hbcee;
13274: douta=16'hbcef;
13275: douta=16'hd612;
13276: douta=16'hddf3;
13277: douta=16'hde34;
13278: douta=16'hcd91;
13279: douta=16'heed7;
13280: douta=16'hddf3;
13281: douta=16'hee95;
13282: douta=16'he675;
13283: douta=16'heeb5;
13284: douta=16'he654;
13285: douta=16'he613;
13286: douta=16'hd5d1;
13287: douta=16'hd591;
13288: douta=16'ha40f;
13289: douta=16'h940e;
13290: douta=16'h7b90;
13291: douta=16'h6b0c;
13292: douta=16'h6b2c;
13293: douta=16'h6b0c;
13294: douta=16'h49e9;
13295: douta=16'h8306;
13296: douta=16'hb44b;
13297: douta=16'hc4ed;
13298: douta=16'hd54f;
13299: douta=16'hddf2;
13300: douta=16'he654;
13301: douta=16'he654;
13302: douta=16'hee95;
13303: douta=16'he654;
13304: douta=16'hee75;
13305: douta=16'hee54;
13306: douta=16'hddf3;
13307: douta=16'hd571;
13308: douta=16'hd591;
13309: douta=16'hac91;
13310: douta=16'h9431;
13311: douta=16'ha471;
13312: douta=16'h8c31;
13313: douta=16'h9432;
13314: douta=16'h83f1;
13315: douta=16'h7c12;
13316: douta=16'h73d1;
13317: douta=16'h73b0;
13318: douta=16'h736f;
13319: douta=16'h6b2e;
13320: douta=16'h5aee;
13321: douta=16'h7a87;
13322: douta=16'h9368;
13323: douta=16'hd56e;
13324: douta=16'h9c4f;
13325: douta=16'h4ace;
13326: douta=16'h322b;
13327: douta=16'h4aee;
13328: douta=16'h2168;
13329: douta=16'h10e5;
13330: douta=16'h10c5;
13331: douta=16'h2988;
13332: douta=16'h5ace;
13333: douta=16'h0062;
13334: douta=16'h18e5;
13335: douta=16'h18e5;
13336: douta=16'h18e5;
13337: douta=16'h18e5;
13338: douta=16'h10e4;
13339: douta=16'h10c4;
13340: douta=16'h1905;
13341: douta=16'h0022;
13342: douta=16'h4b31;
13343: douta=16'h5b70;
13344: douta=16'h4a6c;
13345: douta=16'h4a6a;
13346: douta=16'h8c70;
13347: douta=16'h7b8e;
13348: douta=16'h2189;
13349: douta=16'ha61c;
13350: douta=16'h8d18;
13351: douta=16'h8518;
13352: douta=16'h84d7;
13353: douta=16'h8d39;
13354: douta=16'h8d38;
13355: douta=16'h9579;
13356: douta=16'h8d38;
13357: douta=16'h8cd7;
13358: douta=16'h8496;
13359: douta=16'h84f7;
13360: douta=16'h8d18;
13361: douta=16'h7476;
13362: douta=16'h7c96;
13363: douta=16'h84d7;
13364: douta=16'h84f8;
13365: douta=16'h84d7;
13366: douta=16'h84b7;
13367: douta=16'h7c76;
13368: douta=16'h6c35;
13369: douta=16'h6c35;
13370: douta=16'h84f8;
13371: douta=16'h8518;
13372: douta=16'h7cd7;
13373: douta=16'h7476;
13374: douta=16'h8518;
13375: douta=16'h84f9;
13376: douta=16'h8d39;
13377: douta=16'h8539;
13378: douta=16'h8539;
13379: douta=16'h8d7a;
13380: douta=16'h8539;
13381: douta=16'h7cf8;
13382: douta=16'h8518;
13383: douta=16'h8c73;
13384: douta=16'h52ad;
13385: douta=16'h1861;
13386: douta=16'h39e9;
13387: douta=16'h8539;
13388: douta=16'h8d5a;
13389: douta=16'h8519;
13390: douta=16'h9dbb;
13391: douta=16'h959a;
13392: douta=16'h84f9;
13393: douta=16'h8d59;
13394: douta=16'h959a;
13395: douta=16'h8d7a;
13396: douta=16'h8d59;
13397: douta=16'h8d7a;
13398: douta=16'h9d9a;
13399: douta=16'h7cd9;
13400: douta=16'h9ddb;
13401: douta=16'h959a;
13402: douta=16'h959a;
13403: douta=16'h9ddb;
13404: douta=16'h957a;
13405: douta=16'h95bb;
13406: douta=16'h957a;
13407: douta=16'h9d9a;
13408: douta=16'h959a;
13409: douta=16'h8d59;
13410: douta=16'h8519;
13411: douta=16'h959a;
13412: douta=16'h95bb;
13413: douta=16'h8519;
13414: douta=16'h6c37;
13415: douta=16'h957b;
13416: douta=16'h8d7b;
13417: douta=16'h74b8;
13418: douta=16'h6b2e;
13419: douta=16'h6244;
13420: douta=16'h3124;
13421: douta=16'h18c3;
13422: douta=16'h0882;
13423: douta=16'h6c57;
13424: douta=16'h942e;
13425: douta=16'h3880;
13426: douta=16'h6416;
13427: douta=16'h4311;
13428: douta=16'h5bb4;
13429: douta=16'hae3d;
13430: douta=16'h6c15;
13431: douta=16'h95dd;
13432: douta=16'h29a9;
13433: douta=16'h4b32;
13434: douta=16'hb65c;
13435: douta=16'h9dbb;
13436: douta=16'h9dbb;
13437: douta=16'h6436;
13438: douta=16'h6415;
13439: douta=16'h0000;
13440: douta=16'h3966;
13441: douta=16'h3146;
13442: douta=16'h18c4;
13443: douta=16'h29eb;
13444: douta=16'h220d;
13445: douta=16'h4312;
13446: douta=16'h3290;
13447: douta=16'h4332;
13448: douta=16'h6416;
13449: douta=16'h6c36;
13450: douta=16'h7cd9;
13451: douta=16'h63b3;
13452: douta=16'h4acf;
13453: douta=16'h7413;
13454: douta=16'h73d1;
13455: douta=16'h8c75;
13456: douta=16'hee96;
13457: douta=16'hee75;
13458: douta=16'hde13;
13459: douta=16'hd5d1;
13460: douta=16'hcd71;
13461: douta=16'hb4ad;
13462: douta=16'h7b07;
13463: douta=16'hbcee;
13464: douta=16'hbcee;
13465: douta=16'hc52f;
13466: douta=16'hcd71;
13467: douta=16'he655;
13468: douta=16'hde13;
13469: douta=16'he696;
13470: douta=16'he696;
13471: douta=16'he675;
13472: douta=16'hee96;
13473: douta=16'hddd2;
13474: douta=16'hee95;
13475: douta=16'heed6;
13476: douta=16'hddf2;
13477: douta=16'hcd70;
13478: douta=16'hbcf0;
13479: douta=16'hac8f;
13480: douta=16'h8bf0;
13481: douta=16'h7b8f;
13482: douta=16'h6b2e;
13483: douta=16'h6b0c;
13484: douta=16'h5a6a;
13485: douta=16'h3125;
13486: douta=16'habea;
13487: douta=16'hbc8c;
13488: douta=16'hcd2d;
13489: douta=16'he654;
13490: douta=16'hee95;
13491: douta=16'he675;
13492: douta=16'he674;
13493: douta=16'hee75;
13494: douta=16'hee95;
13495: douta=16'he633;
13496: douta=16'hee75;
13497: douta=16'hd5b3;
13498: douta=16'hc552;
13499: douta=16'hbd12;
13500: douta=16'hbd11;
13501: douta=16'ha492;
13502: douta=16'h9c93;
13503: douta=16'h9472;
13504: douta=16'h8432;
13505: douta=16'h8432;
13506: douta=16'h7391;
13507: douta=16'h6b2e;
13508: douta=16'h630e;
13509: douta=16'h62ec;
13510: douta=16'h5a6a;
13511: douta=16'h6226;
13512: douta=16'hb46b;
13513: douta=16'hddd0;
13514: douta=16'he633;
13515: douta=16'he634;
13516: douta=16'hbcf0;
13517: douta=16'h7391;
13518: douta=16'h6330;
13519: douta=16'h8412;
13520: douta=16'h3a2c;
13521: douta=16'h31ca;
13522: douta=16'h3a2c;
13523: douta=16'h2989;
13524: douta=16'h2127;
13525: douta=16'h0863;
13526: douta=16'h5b51;
13527: douta=16'h0842;
13528: douta=16'h10c5;
13529: douta=16'h10c4;
13530: douta=16'h18e5;
13531: douta=16'h18e4;
13532: douta=16'h10a4;
13533: douta=16'h18e5;
13534: douta=16'h0001;
13535: douta=16'h0862;
13536: douta=16'h7c74;
13537: douta=16'h42cf;
13538: douta=16'h424a;
13539: douta=16'h52ac;
13540: douta=16'h2988;
13541: douta=16'h7bae;
13542: douta=16'h29ca;
13543: douta=16'hae3d;
13544: douta=16'hae3d;
13545: douta=16'h7cf8;
13546: douta=16'h9579;
13547: douta=16'h8d59;
13548: douta=16'h8d38;
13549: douta=16'h8d18;
13550: douta=16'h9538;
13551: douta=16'h84f7;
13552: douta=16'ha5fb;
13553: douta=16'h7476;
13554: douta=16'h7cb7;
13555: douta=16'h84f8;
13556: douta=16'h959a;
13557: douta=16'h7cb7;
13558: douta=16'h9579;
13559: douta=16'ha59a;
13560: douta=16'h7c96;
13561: douta=16'h84d7;
13562: douta=16'h84d7;
13563: douta=16'h7435;
13564: douta=16'h7c96;
13565: douta=16'h7476;
13566: douta=16'h6c15;
13567: douta=16'h84d8;
13568: douta=16'h8519;
13569: douta=16'h8d7b;
13570: douta=16'h7cb7;
13571: douta=16'h8d5a;
13572: douta=16'h8d5a;
13573: douta=16'h84f9;
13574: douta=16'h8d39;
13575: douta=16'h8d18;
13576: douta=16'h5208;
13577: douta=16'h3146;
13578: douta=16'h7455;
13579: douta=16'h84f8;
13580: douta=16'h8539;
13581: douta=16'h8d59;
13582: douta=16'h957a;
13583: douta=16'h9559;
13584: douta=16'h8d39;
13585: douta=16'h959a;
13586: douta=16'h8519;
13587: douta=16'h74b8;
13588: douta=16'h8d59;
13589: douta=16'h8d5a;
13590: douta=16'h8d19;
13591: douta=16'ha61c;
13592: douta=16'h9dba;
13593: douta=16'h9ddb;
13594: douta=16'h8539;
13595: douta=16'h959a;
13596: douta=16'h957a;
13597: douta=16'h959a;
13598: douta=16'h957a;
13599: douta=16'h9dbb;
13600: douta=16'h8d3a;
13601: douta=16'h9ddb;
13602: douta=16'h9ddb;
13603: douta=16'h959a;
13604: douta=16'h8d5a;
13605: douta=16'h8559;
13606: douta=16'h8dbc;
13607: douta=16'had57;
13608: douta=16'h7b6e;
13609: douta=16'h5417;
13610: douta=16'h6498;
13611: douta=16'h6b2c;
13612: douta=16'h51e4;
13613: douta=16'h4144;
13614: douta=16'h1083;
13615: douta=16'h0000;
13616: douta=16'h7cda;
13617: douta=16'h74fa;
13618: douta=16'h4b53;
13619: douta=16'h84f8;
13620: douta=16'h6c35;
13621: douta=16'h8d18;
13622: douta=16'h74ba;
13623: douta=16'h7390;
13624: douta=16'h855a;
13625: douta=16'h6415;
13626: douta=16'h7497;
13627: douta=16'h7cb8;
13628: douta=16'h7c98;
13629: douta=16'hb65d;
13630: douta=16'h4aef;
13631: douta=16'h0821;
13632: douta=16'h3985;
13633: douta=16'h3145;
13634: douta=16'h3146;
13635: douta=16'h29a9;
13636: douta=16'h21ed;
13637: douta=16'h32b0;
13638: douta=16'h32d1;
13639: douta=16'h63f6;
13640: douta=16'h3aaf;
13641: douta=16'h4af0;
13642: douta=16'h7477;
13643: douta=16'h42af;
13644: douta=16'h5330;
13645: douta=16'h6bd3;
13646: douta=16'ha557;
13647: douta=16'had98;
13648: douta=16'hee73;
13649: douta=16'hee75;
13650: douta=16'he654;
13651: douta=16'hc550;
13652: douta=16'hc50e;
13653: douta=16'h8b6a;
13654: douta=16'hbcee;
13655: douta=16'hbd0f;
13656: douta=16'hbd0e;
13657: douta=16'hcd90;
13658: douta=16'he634;
13659: douta=16'hde54;
13660: douta=16'hde14;
13661: douta=16'heeb7;
13662: douta=16'he655;
13663: douta=16'heeb6;
13664: douta=16'hee75;
13665: douta=16'he635;
13666: douta=16'hac2d;
13667: douta=16'hac2d;
13668: douta=16'hee94;
13669: douta=16'hbcf0;
13670: douta=16'hac70;
13671: douta=16'h9c50;
13672: douta=16'h7b8f;
13673: douta=16'h6b4d;
13674: douta=16'h62cc;
13675: douta=16'h4a09;
13676: douta=16'h6206;
13677: douta=16'hc4ab;
13678: douta=16'hbc8b;
13679: douta=16'hcd2e;
13680: douta=16'he633;
13681: douta=16'hee75;
13682: douta=16'he654;
13683: douta=16'heeb6;
13684: douta=16'hee74;
13685: douta=16'hde13;
13686: douta=16'hddf3;
13687: douta=16'hbcf1;
13688: douta=16'hcd52;
13689: douta=16'hcd72;
13690: douta=16'hacd2;
13691: douta=16'hb4f2;
13692: douta=16'ha4b3;
13693: douta=16'h9c94;
13694: douta=16'h9473;
13695: douta=16'h8433;
13696: douta=16'h73b1;
13697: douta=16'h736f;
13698: douta=16'h6b2f;
13699: douta=16'h6b0d;
13700: douta=16'h6b0e;
13701: douta=16'h62ad;
13702: douta=16'h8b28;
13703: douta=16'hc46c;
13704: douta=16'hcd6e;
13705: douta=16'hde11;
13706: douta=16'hde12;
13707: douta=16'he612;
13708: douta=16'hcd71;
13709: douta=16'h8c10;
13710: douta=16'h7bd0;
13711: douta=16'h9474;
13712: douta=16'h5b91;
13713: douta=16'h3a6c;
13714: douta=16'h324c;
13715: douta=16'h324d;
13716: douta=16'h322b;
13717: douta=16'h1947;
13718: douta=16'h08a4;
13719: douta=16'h5b51;
13720: douta=16'h10a4;
13721: douta=16'h18e5;
13722: douta=16'h10c5;
13723: douta=16'h18c5;
13724: douta=16'h10e4;
13725: douta=16'h10c5;
13726: douta=16'h10e5;
13727: douta=16'h1906;
13728: douta=16'h0042;
13729: douta=16'h7c54;
13730: douta=16'h31ea;
13731: douta=16'h0000;
13732: douta=16'h52ed;
13733: douta=16'h4a6a;
13734: douta=16'h73f3;
13735: douta=16'h41c8;
13736: douta=16'h2169;
13737: douta=16'h9d9a;
13738: douta=16'h9d79;
13739: douta=16'h8d18;
13740: douta=16'h9559;
13741: douta=16'h84d6;
13742: douta=16'h7c96;
13743: douta=16'h8d18;
13744: douta=16'h84b7;
13745: douta=16'h84d7;
13746: douta=16'h7476;
13747: douta=16'h9579;
13748: douta=16'h7c76;
13749: douta=16'h8d38;
13750: douta=16'h8d38;
13751: douta=16'h8d18;
13752: douta=16'h9579;
13753: douta=16'h9559;
13754: douta=16'h8d39;
13755: douta=16'h9559;
13756: douta=16'h84d7;
13757: douta=16'h7cb7;
13758: douta=16'h9d9a;
13759: douta=16'h6391;
13760: douta=16'h63b2;
13761: douta=16'h6bd2;
13762: douta=16'h7cb7;
13763: douta=16'h8d7a;
13764: douta=16'h7cb8;
13765: douta=16'h7cd8;
13766: douta=16'h8519;
13767: douta=16'h8539;
13768: douta=16'h857b;
13769: douta=16'h95bc;
13770: douta=16'h7cd8;
13771: douta=16'h95bb;
13772: douta=16'h74b8;
13773: douta=16'h84f9;
13774: douta=16'h84d8;
13775: douta=16'h957a;
13776: douta=16'h8d59;
13777: douta=16'h8d19;
13778: douta=16'h8d19;
13779: douta=16'h8519;
13780: douta=16'h959a;
13781: douta=16'h957a;
13782: douta=16'h959a;
13783: douta=16'h8d5a;
13784: douta=16'ha5db;
13785: douta=16'h957a;
13786: douta=16'ha5fc;
13787: douta=16'ha5db;
13788: douta=16'h9dbb;
13789: douta=16'h9dda;
13790: douta=16'h959a;
13791: douta=16'h959a;
13792: douta=16'hb65c;
13793: douta=16'h959a;
13794: douta=16'h8d7a;
13795: douta=16'h957a;
13796: douta=16'ha5dc;
13797: douta=16'h9dfc;
13798: douta=16'h5b0e;
13799: douta=16'h5c38;
13800: douta=16'h5c79;
13801: douta=16'h5c16;
13802: douta=16'h5373;
13803: douta=16'h6cba;
13804: douta=16'h7b08;
13805: douta=16'h6245;
13806: douta=16'h20e3;
13807: douta=16'h0862;
13808: douta=16'h5331;
13809: douta=16'h857c;
13810: douta=16'h61c3;
13811: douta=16'h10a5;
13812: douta=16'h8518;
13813: douta=16'h7456;
13814: douta=16'h7c32;
13815: douta=16'h3040;
13816: douta=16'h21ec;
13817: douta=16'h5352;
13818: douta=16'h63d3;
13819: douta=16'hbe5c;
13820: douta=16'h84d8;
13821: douta=16'h6c78;
13822: douta=16'h29a8;
13823: douta=16'h4acd;
13824: douta=16'h3965;
13825: douta=16'h3165;
13826: douta=16'h2926;
13827: douta=16'h3a4d;
13828: douta=16'h324f;
13829: douta=16'h3af1;
13830: douta=16'h53d6;
13831: douta=16'h4b73;
13832: douta=16'h4b32;
13833: douta=16'h63f4;
13834: douta=16'h7cb8;
13835: douta=16'h5331;
13836: douta=16'h5351;
13837: douta=16'h5b72;
13838: douta=16'h8c73;
13839: douta=16'h9d16;
13840: douta=16'hddd1;
13841: douta=16'he675;
13842: douta=16'hddf3;
13843: douta=16'ha42c;
13844: douta=16'ha44c;
13845: douta=16'h8348;
13846: douta=16'hbcee;
13847: douta=16'hbd0f;
13848: douta=16'hc50e;
13849: douta=16'hd5d2;
13850: douta=16'he675;
13851: douta=16'hde54;
13852: douta=16'he655;
13853: douta=16'heeb7;
13854: douta=16'he655;
13855: douta=16'hee96;
13856: douta=16'hee75;
13857: douta=16'hddf3;
13858: douta=16'hcd50;
13859: douta=16'h9c0d;
13860: douta=16'hd591;
13861: douta=16'hac50;
13862: douta=16'h9c70;
13863: douta=16'h9c50;
13864: douta=16'h736d;
13865: douta=16'h6b2c;
13866: douta=16'h62cc;
13867: douta=16'h2905;
13868: douta=16'hb42a;
13869: douta=16'hcd2d;
13870: douta=16'hc4ed;
13871: douta=16'hcd4f;
13872: douta=16'he654;
13873: douta=16'hf6b6;
13874: douta=16'hee96;
13875: douta=16'he654;
13876: douta=16'he654;
13877: douta=16'hddb1;
13878: douta=16'hddb1;
13879: douta=16'hbd12;
13880: douta=16'hac91;
13881: douta=16'hd5b2;
13882: douta=16'h9c92;
13883: douta=16'hacd3;
13884: douta=16'ha4d3;
13885: douta=16'h9473;
13886: douta=16'h8c53;
13887: douta=16'h8412;
13888: douta=16'h7390;
13889: douta=16'h736f;
13890: douta=16'h732e;
13891: douta=16'h632e;
13892: douta=16'h5229;
13893: douta=16'h6228;
13894: douta=16'hb3eb;
13895: douta=16'hcd0e;
13896: douta=16'hddd1;
13897: douta=16'he654;
13898: douta=16'he634;
13899: douta=16'he613;
13900: douta=16'hcd71;
13901: douta=16'h8c10;
13902: douta=16'h83f1;
13903: douta=16'h8c32;
13904: douta=16'h7433;
13905: douta=16'h3a6d;
13906: douta=16'h426d;
13907: douta=16'h322c;
13908: douta=16'h2a0b;
13909: douta=16'h21a9;
13910: douta=16'h2127;
13911: douta=16'h2107;
13912: douta=16'h10c4;
13913: douta=16'h1063;
13914: douta=16'h10c4;
13915: douta=16'h10c5;
13916: douta=16'h10c5;
13917: douta=16'h10e4;
13918: douta=16'h18e4;
13919: douta=16'h10a4;
13920: douta=16'h2147;
13921: douta=16'h10e5;
13922: douta=16'h2167;
13923: douta=16'h0842;
13924: douta=16'h10c4;
13925: douta=16'h0883;
13926: douta=16'h9cf5;
13927: douta=16'hb573;
13928: douta=16'h9c90;
13929: douta=16'h29aa;
13930: douta=16'ha5db;
13931: douta=16'ha5da;
13932: douta=16'ha5ba;
13933: douta=16'h9559;
13934: douta=16'h8d18;
13935: douta=16'h9559;
13936: douta=16'h84d7;
13937: douta=16'h84d7;
13938: douta=16'h7c96;
13939: douta=16'h8d59;
13940: douta=16'h8d18;
13941: douta=16'h7cb7;
13942: douta=16'h9dba;
13943: douta=16'h9dba;
13944: douta=16'h7cb6;
13945: douta=16'h9559;
13946: douta=16'h8d39;
13947: douta=16'h84f8;
13948: douta=16'h8d18;
13949: douta=16'h84b7;
13950: douta=16'h7476;
13951: douta=16'h7c55;
13952: douta=16'h6bb3;
13953: douta=16'h7434;
13954: douta=16'h6bd4;
13955: douta=16'h5b93;
13956: douta=16'h7cb7;
13957: douta=16'h7d18;
13958: douta=16'h8519;
13959: douta=16'h7cf8;
13960: douta=16'h8539;
13961: douta=16'h8d5b;
13962: douta=16'h851a;
13963: douta=16'h8539;
13964: douta=16'h84f8;
13965: douta=16'h95bb;
13966: douta=16'h8539;
13967: douta=16'h84f8;
13968: douta=16'h84f8;
13969: douta=16'h8d59;
13970: douta=16'h9d9a;
13971: douta=16'h8518;
13972: douta=16'h959a;
13973: douta=16'h9dbb;
13974: douta=16'h8d59;
13975: douta=16'h8d5a;
13976: douta=16'h959a;
13977: douta=16'h9dbb;
13978: douta=16'h959a;
13979: douta=16'hadfc;
13980: douta=16'h9d9a;
13981: douta=16'h959a;
13982: douta=16'h9dbb;
13983: douta=16'h8d5a;
13984: douta=16'h8d5a;
13985: douta=16'hae3c;
13986: douta=16'hb67d;
13987: douta=16'ha61d;
13988: douta=16'ha61c;
13989: douta=16'h632e;
13990: douta=16'h4bf7;
13991: douta=16'h6478;
13992: douta=16'h5c57;
13993: douta=16'h53f5;
13994: douta=16'h6498;
13995: douta=16'h5c78;
13996: douta=16'h8308;
13997: douta=16'h72a6;
13998: douta=16'h2923;
13999: douta=16'h0862;
14000: douta=16'h1926;
14001: douta=16'h4bd4;
14002: douta=16'ha535;
14003: douta=16'h4060;
14004: douta=16'h7d3c;
14005: douta=16'h63d4;
14006: douta=16'h734b;
14007: douta=16'h1800;
14008: douta=16'h5bb3;
14009: douta=16'h5bb4;
14010: douta=16'h4b32;
14011: douta=16'h6bd3;
14012: douta=16'h7455;
14013: douta=16'h5310;
14014: douta=16'h7433;
14015: douta=16'h5b8f;
14016: douta=16'h3945;
14017: douta=16'h3966;
14018: douta=16'h2945;
14019: douta=16'h1083;
14020: douta=16'h5bf7;
14021: douta=16'h32b0;
14022: douta=16'h4333;
14023: douta=16'h5373;
14024: douta=16'h5c15;
14025: douta=16'h5bd4;
14026: douta=16'h7498;
14027: douta=16'h5351;
14028: douta=16'h5b92;
14029: douta=16'h5b72;
14030: douta=16'h9d36;
14031: douta=16'h8cb4;
14032: douta=16'had57;
14033: douta=16'hee95;
14034: douta=16'h836c;
14035: douta=16'hac6c;
14036: douta=16'hbcee;
14037: douta=16'hc530;
14038: douta=16'hcd91;
14039: douta=16'hd5b1;
14040: douta=16'hcdb1;
14041: douta=16'hee96;
14042: douta=16'heeb7;
14043: douta=16'hee96;
14044: douta=16'he675;
14045: douta=16'heeb7;
14046: douta=16'hee97;
14047: douta=16'hee96;
14048: douta=16'hd613;
14049: douta=16'hd5d2;
14050: douta=16'hbd30;
14051: douta=16'hbd30;
14052: douta=16'hb4f1;
14053: douta=16'ha430;
14054: douta=16'ha4b1;
14055: douta=16'h7baf;
14056: douta=16'h62eb;
14057: douta=16'h6b0d;
14058: douta=16'h3125;
14059: douta=16'hbcab;
14060: douta=16'hc4cc;
14061: douta=16'hc4ec;
14062: douta=16'hddd2;
14063: douta=16'hde14;
14064: douta=16'hee95;
14065: douta=16'heeb7;
14066: douta=16'he654;
14067: douta=16'he614;
14068: douta=16'hddf2;
14069: douta=16'hcd30;
14070: douta=16'hcd50;
14071: douta=16'hbd11;
14072: douta=16'hbcf1;
14073: douta=16'h8bf1;
14074: douta=16'hbd53;
14075: douta=16'h8c52;
14076: douta=16'h9473;
14077: douta=16'h8c53;
14078: douta=16'h7bf1;
14079: douta=16'h7bd0;
14080: douta=16'h732e;
14081: douta=16'h630e;
14082: douta=16'h6b0d;
14083: douta=16'h7aa7;
14084: douta=16'hac09;
14085: douta=16'hb46b;
14086: douta=16'hddaf;
14087: douta=16'he612;
14088: douta=16'he654;
14089: douta=16'he613;
14090: douta=16'hde13;
14091: douta=16'hddd1;
14092: douta=16'hc511;
14093: douta=16'ha470;
14094: douta=16'ha491;
14095: douta=16'h8453;
14096: douta=16'h8454;
14097: douta=16'h7c34;
14098: douta=16'h5b71;
14099: douta=16'h42cf;
14100: douta=16'h42ae;
14101: douta=16'h3a2c;
14102: douta=16'h322c;
14103: douta=16'h2167;
14104: douta=16'h08a3;
14105: douta=16'h29a9;
14106: douta=16'h2167;
14107: douta=16'h18e5;
14108: douta=16'h18e5;
14109: douta=16'h10e4;
14110: douta=16'h10c5;
14111: douta=16'h18e4;
14112: douta=16'h10c5;
14113: douta=16'h10c4;
14114: douta=16'h2126;
14115: douta=16'h0883;
14116: douta=16'h1926;
14117: douta=16'h1905;
14118: douta=16'h10a4;
14119: douta=16'hd655;
14120: douta=16'h944e;
14121: douta=16'hc5f4;
14122: douta=16'h39e8;
14123: douta=16'h630d;
14124: douta=16'h428d;
14125: douta=16'h8d39;
14126: douta=16'h84d7;
14127: douta=16'h9579;
14128: douta=16'h9dba;
14129: douta=16'h9d9a;
14130: douta=16'h84f8;
14131: douta=16'h7455;
14132: douta=16'h9d9a;
14133: douta=16'h8d38;
14134: douta=16'h84d7;
14135: douta=16'h84f7;
14136: douta=16'h8d38;
14137: douta=16'h84f8;
14138: douta=16'h7c96;
14139: douta=16'h7455;
14140: douta=16'h9559;
14141: douta=16'h9559;
14142: douta=16'h8d39;
14143: douta=16'h7cb7;
14144: douta=16'h7496;
14145: douta=16'h8d59;
14146: douta=16'h7c75;
14147: douta=16'h8d39;
14148: douta=16'h7c97;
14149: douta=16'h7496;
14150: douta=16'h7477;
14151: douta=16'h7c77;
14152: douta=16'h8519;
14153: douta=16'h8d3a;
14154: douta=16'h8519;
14155: douta=16'h8519;
14156: douta=16'h8539;
14157: douta=16'h8d3a;
14158: douta=16'h8539;
14159: douta=16'h8519;
14160: douta=16'h7497;
14161: douta=16'h959a;
14162: douta=16'h959a;
14163: douta=16'h8d7a;
14164: douta=16'h7cb7;
14165: douta=16'h8519;
14166: douta=16'h8519;
14167: douta=16'h8d39;
14168: douta=16'h959a;
14169: douta=16'h959b;
14170: douta=16'h9ddb;
14171: douta=16'h8559;
14172: douta=16'h959b;
14173: douta=16'h959a;
14174: douta=16'h8d18;
14175: douta=16'h9d9a;
14176: douta=16'hae7e;
14177: douta=16'h8474;
14178: douta=16'h62ec;
14179: douta=16'h6cb9;
14180: douta=16'h53f6;
14181: douta=16'h6457;
14182: douta=16'h5c37;
14183: douta=16'h74fb;
14184: douta=16'h4bd6;
14185: douta=16'h4374;
14186: douta=16'h5c17;
14187: douta=16'h64b8;
14188: douta=16'h62cc;
14189: douta=16'h7ac5;
14190: douta=16'h6a44;
14191: douta=16'h1082;
14192: douta=16'h1063;
14193: douta=16'h0000;
14194: douta=16'h7477;
14195: douta=16'h53f5;
14196: douta=16'h7aeb;
14197: douta=16'h85bd;
14198: douta=16'h1882;
14199: douta=16'h6478;
14200: douta=16'h6435;
14201: douta=16'h7497;
14202: douta=16'h9dba;
14203: douta=16'h5b2e;
14204: douta=16'h8472;
14205: douta=16'h9d14;
14206: douta=16'hc638;
14207: douta=16'ha5d8;
14208: douta=16'h526b;
14209: douta=16'h3966;
14210: douta=16'h3145;
14211: douta=16'h1882;
14212: douta=16'h4332;
14213: douta=16'h4333;
14214: douta=16'h3ad1;
14215: douta=16'h2a4f;
14216: douta=16'h5bb4;
14217: douta=16'h6436;
14218: douta=16'h63f5;
14219: douta=16'h6c35;
14220: douta=16'h6bf4;
14221: douta=16'h6bd3;
14222: douta=16'h8433;
14223: douta=16'h9cb5;
14224: douta=16'h8c73;
14225: douta=16'hb5b8;
14226: douta=16'hc551;
14227: douta=16'hc54f;
14228: douta=16'hc530;
14229: douta=16'hc551;
14230: douta=16'hd5d2;
14231: douta=16'hde15;
14232: douta=16'hde14;
14233: douta=16'heed7;
14234: douta=16'heeb6;
14235: douta=16'hee96;
14236: douta=16'hee96;
14237: douta=16'hd591;
14238: douta=16'hde34;
14239: douta=16'hde13;
14240: douta=16'hd5b2;
14241: douta=16'hbd11;
14242: douta=16'ha4b1;
14243: douta=16'h9450;
14244: douta=16'h9450;
14245: douta=16'h7b8f;
14246: douta=16'h838e;
14247: douta=16'h7baf;
14248: douta=16'h528a;
14249: douta=16'h3945;
14250: douta=16'hbc6a;
14251: douta=16'hc50e;
14252: douta=16'hd570;
14253: douta=16'hd56f;
14254: douta=16'he674;
14255: douta=16'hee74;
14256: douta=16'hee75;
14257: douta=16'he674;
14258: douta=16'hf6b6;
14259: douta=16'hddd2;
14260: douta=16'hdd91;
14261: douta=16'hcd71;
14262: douta=16'hb4cf;
14263: douta=16'hb4f2;
14264: douta=16'ha491;
14265: douta=16'h9c72;
14266: douta=16'h8412;
14267: douta=16'ha4b4;
14268: douta=16'h83f1;
14269: douta=16'h8c52;
14270: douta=16'h7bd1;
14271: douta=16'h6b2e;
14272: douta=16'h632e;
14273: douta=16'h4a4a;
14274: douta=16'h59a5;
14275: douta=16'ha3ea;
14276: douta=16'hc4cc;
14277: douta=16'hdd90;
14278: douta=16'he653;
14279: douta=16'he654;
14280: douta=16'he634;
14281: douta=16'hddf3;
14282: douta=16'hddd3;
14283: douta=16'hd591;
14284: douta=16'hb4af;
14285: douta=16'ha491;
14286: douta=16'hac92;
14287: douta=16'h8433;
14288: douta=16'h7c13;
14289: douta=16'h7c34;
14290: douta=16'h73f3;
14291: douta=16'h5bb2;
14292: douta=16'h5b71;
14293: douta=16'h4aef;
14294: douta=16'h3a6d;
14295: douta=16'h324d;
14296: douta=16'h3a8e;
14297: douta=16'h3aae;
14298: douta=16'h21ca;
14299: douta=16'h10a4;
14300: douta=16'h10e5;
14301: douta=16'h10c4;
14302: douta=16'h10c4;
14303: douta=16'h10c4;
14304: douta=16'h10c4;
14305: douta=16'h10c5;
14306: douta=16'h18e5;
14307: douta=16'h1905;
14308: douta=16'h10c5;
14309: douta=16'h0883;
14310: douta=16'h10a5;
14311: douta=16'h63b3;
14312: douta=16'h7412;
14313: douta=16'h52cd;
14314: douta=16'h736c;
14315: douta=16'h52cb;
14316: douta=16'h7bef;
14317: douta=16'h5aec;
14318: douta=16'h6391;
14319: douta=16'h84d8;
14320: douta=16'h84d8;
14321: douta=16'h8497;
14322: douta=16'h84f7;
14323: douta=16'h84d7;
14324: douta=16'h8d18;
14325: douta=16'ha5da;
14326: douta=16'h9d99;
14327: douta=16'h8cf7;
14328: douta=16'h84b6;
14329: douta=16'h8cf7;
14330: douta=16'h84b7;
14331: douta=16'h7c96;
14332: douta=16'h84d7;
14333: douta=16'h84d7;
14334: douta=16'h7c96;
14335: douta=16'h7476;
14336: douta=16'h8d39;
14337: douta=16'h8d39;
14338: douta=16'h7cd7;
14339: douta=16'ha5db;
14340: douta=16'ha5db;
14341: douta=16'h7476;
14342: douta=16'h7c96;
14343: douta=16'h8d18;
14344: douta=16'h84f8;
14345: douta=16'h7476;
14346: douta=16'h7456;
14347: douta=16'h8519;
14348: douta=16'h8519;
14349: douta=16'h7cd8;
14350: douta=16'h7cf9;
14351: douta=16'h8d5a;
14352: douta=16'h8d5a;
14353: douta=16'h8519;
14354: douta=16'h8519;
14355: douta=16'h7cf9;
14356: douta=16'h957b;
14357: douta=16'h959b;
14358: douta=16'h84f9;
14359: douta=16'h8d3a;
14360: douta=16'h74b8;
14361: douta=16'h6457;
14362: douta=16'h957a;
14363: douta=16'h959b;
14364: douta=16'h959a;
14365: douta=16'h959c;
14366: douta=16'h8d9c;
14367: douta=16'h8cf6;
14368: douta=16'h3a4c;
14369: douta=16'h3b12;
14370: douta=16'h4c16;
14371: douta=16'h6cf9;
14372: douta=16'h74b9;
14373: douta=16'h5c37;
14374: douta=16'h753b;
14375: douta=16'h3b13;
14376: douta=16'h4374;
14377: douta=16'h4b95;
14378: douta=16'h4395;
14379: douta=16'h7d5b;
14380: douta=16'h651c;
14381: douta=16'h732c;
14382: douta=16'h8329;
14383: douta=16'h28e3;
14384: douta=16'h0882;
14385: douta=16'h0862;
14386: douta=16'h5c16;
14387: douta=16'h6436;
14388: douta=16'h5418;
14389: douta=16'h40c0;
14390: douta=16'h5c57;
14391: douta=16'h7498;
14392: douta=16'h8d18;
14393: douta=16'h63b1;
14394: douta=16'h73f0;
14395: douta=16'hbdd6;
14396: douta=16'hadd7;
14397: douta=16'h8cb3;
14398: douta=16'h39a6;
14399: douta=16'h1840;
14400: douta=16'h5b0e;
14401: douta=16'h3986;
14402: douta=16'h3146;
14403: douta=16'h1883;
14404: douta=16'h326e;
14405: douta=16'h3ad1;
14406: douta=16'h4b53;
14407: douta=16'h3290;
14408: douta=16'h5bd5;
14409: douta=16'h7477;
14410: douta=16'h7455;
14411: douta=16'h63f4;
14412: douta=16'h8475;
14413: douta=16'h7c75;
14414: douta=16'h73f2;
14415: douta=16'had77;
14416: douta=16'h6bb1;
14417: douta=16'hc63a;
14418: douta=16'hc572;
14419: douta=16'hc570;
14420: douta=16'hcd90;
14421: douta=16'hcdb2;
14422: douta=16'hd5d3;
14423: douta=16'he656;
14424: douta=16'he655;
14425: douta=16'heed7;
14426: douta=16'heed7;
14427: douta=16'hee96;
14428: douta=16'heeb6;
14429: douta=16'hd5d2;
14430: douta=16'hc54f;
14431: douta=16'he674;
14432: douta=16'hc551;
14433: douta=16'ha4b1;
14434: douta=16'ha4b1;
14435: douta=16'h9c51;
14436: douta=16'h7baf;
14437: douta=16'h8c10;
14438: douta=16'h7b6e;
14439: douta=16'h734d;
14440: douta=16'h41a5;
14441: douta=16'h8ae8;
14442: douta=16'hbcec;
14443: douta=16'hcd4f;
14444: douta=16'hddd2;
14445: douta=16'hd5b1;
14446: douta=16'hee95;
14447: douta=16'he674;
14448: douta=16'he654;
14449: douta=16'hddf3;
14450: douta=16'hee95;
14451: douta=16'hde13;
14452: douta=16'hcd31;
14453: douta=16'hcd31;
14454: douta=16'hbd10;
14455: douta=16'ha4b2;
14456: douta=16'hacb2;
14457: douta=16'h9c93;
14458: douta=16'h7bf2;
14459: douta=16'h9cb3;
14460: douta=16'h9cb4;
14461: douta=16'h7bd0;
14462: douta=16'h8412;
14463: douta=16'h734f;
14464: douta=16'h41e8;
14465: douta=16'h28c3;
14466: douta=16'h9348;
14467: douta=16'hbc8b;
14468: douta=16'hddaf;
14469: douta=16'hddf2;
14470: douta=16'hee54;
14471: douta=16'he633;
14472: douta=16'he633;
14473: douta=16'hddf2;
14474: douta=16'hddd3;
14475: douta=16'hd570;
14476: douta=16'hb4b0;
14477: douta=16'hacb1;
14478: douta=16'ha491;
14479: douta=16'h8c53;
14480: douta=16'h7c13;
14481: douta=16'h7c34;
14482: douta=16'h7414;
14483: douta=16'h5b92;
14484: douta=16'h5b71;
14485: douta=16'h5330;
14486: douta=16'h42ae;
14487: douta=16'h3a6d;
14488: douta=16'h42ae;
14489: douta=16'h3a6d;
14490: douta=16'h21c9;
14491: douta=16'h4b0e;
14492: douta=16'h0862;
14493: douta=16'h1084;
14494: douta=16'h18e5;
14495: douta=16'h18e5;
14496: douta=16'h18e5;
14497: douta=16'h1905;
14498: douta=16'h1906;
14499: douta=16'h1905;
14500: douta=16'h1906;
14501: douta=16'h0883;
14502: douta=16'h0062;
14503: douta=16'h324c;
14504: douta=16'h42b0;
14505: douta=16'h7433;
14506: douta=16'hded7;
14507: douta=16'h738f;
14508: douta=16'h6b2c;
14509: douta=16'h4229;
14510: douta=16'h3187;
14511: douta=16'h5aeb;
14512: douta=16'h7cb7;
14513: douta=16'h8539;
14514: douta=16'hadfb;
14515: douta=16'h9559;
14516: douta=16'h7456;
14517: douta=16'h84f7;
14518: douta=16'h9559;
14519: douta=16'h84b7;
14520: douta=16'h84b7;
14521: douta=16'h84b7;
14522: douta=16'h8d18;
14523: douta=16'h8d38;
14524: douta=16'h7cb7;
14525: douta=16'h957a;
14526: douta=16'h6c35;
14527: douta=16'h6c55;
14528: douta=16'h63f4;
14529: douta=16'h8d39;
14530: douta=16'h8d39;
14531: douta=16'h8d39;
14532: douta=16'h8d39;
14533: douta=16'h6c55;
14534: douta=16'h7cb7;
14535: douta=16'h9559;
14536: douta=16'h6c14;
14537: douta=16'h8d39;
14538: douta=16'h9559;
14539: douta=16'h7455;
14540: douta=16'h7cb7;
14541: douta=16'h8d7a;
14542: douta=16'h7497;
14543: douta=16'h7cd8;
14544: douta=16'h84f9;
14545: douta=16'h8d7a;
14546: douta=16'h8d5a;
14547: douta=16'h8d5a;
14548: douta=16'h8519;
14549: douta=16'h8d59;
14550: douta=16'h8d39;
14551: douta=16'h8d7a;
14552: douta=16'h957a;
14553: douta=16'h7cb8;
14554: douta=16'h74d7;
14555: douta=16'h9ddb;
14556: douta=16'h9e1d;
14557: douta=16'h7c95;
14558: douta=16'h6bb1;
14559: douta=16'h42ae;
14560: douta=16'h3312;
14561: douta=16'h4394;
14562: douta=16'h3b11;
14563: douta=16'h6c99;
14564: douta=16'h4393;
14565: douta=16'h6479;
14566: douta=16'h6cda;
14567: douta=16'h4374;
14568: douta=16'h5c37;
14569: douta=16'h4b94;
14570: douta=16'h6cda;
14571: douta=16'h4354;
14572: douta=16'h4bd7;
14573: douta=16'h63f5;
14574: douta=16'h8b69;
14575: douta=16'h3123;
14576: douta=16'h1082;
14577: douta=16'h0862;
14578: douta=16'h6c99;
14579: douta=16'h5bf5;
14580: douta=16'h74f9;
14581: douta=16'h4942;
14582: douta=16'h5c37;
14583: douta=16'h751b;
14584: douta=16'h8493;
14585: douta=16'h94f3;
14586: douta=16'hbdd6;
14587: douta=16'ha576;
14588: douta=16'h6bcf;
14589: douta=16'h5aaa;
14590: douta=16'h1881;
14591: douta=16'h3124;
14592: douta=16'h6413;
14593: douta=16'h41a6;
14594: douta=16'h3945;
14595: douta=16'h20e4;
14596: douta=16'h3a6e;
14597: douta=16'h53d6;
14598: douta=16'h3ad0;
14599: douta=16'h4353;
14600: douta=16'h4b74;
14601: douta=16'h5bf5;
14602: douta=16'h63d4;
14603: douta=16'h63f4;
14604: douta=16'h6352;
14605: douta=16'h7434;
14606: douta=16'h8454;
14607: douta=16'ha516;
14608: douta=16'h9cf5;
14609: douta=16'hbdd9;
14610: douta=16'h9d37;
14611: douta=16'hd5f3;
14612: douta=16'hde14;
14613: douta=16'hde34;
14614: douta=16'hde34;
14615: douta=16'heed7;
14616: douta=16'heed7;
14617: douta=16'heeb7;
14618: douta=16'heeb7;
14619: douta=16'heeb6;
14620: douta=16'he655;
14621: douta=16'hde13;
14622: douta=16'hddf3;
14623: douta=16'hb4d0;
14624: douta=16'hacd1;
14625: douta=16'ha491;
14626: douta=16'h83d1;
14627: douta=16'h7bd0;
14628: douta=16'h6b4f;
14629: douta=16'h736e;
14630: douta=16'h734d;
14631: douta=16'h628a;
14632: douta=16'hb4ac;
14633: douta=16'hbcce;
14634: douta=16'hcd4e;
14635: douta=16'he633;
14636: douta=16'he654;
14637: douta=16'he634;
14638: douta=16'he653;
14639: douta=16'he654;
14640: douta=16'he613;
14641: douta=16'hd592;
14642: douta=16'hd591;
14643: douta=16'hddf2;
14644: douta=16'hc531;
14645: douta=16'hacb2;
14646: douta=16'ha4b2;
14647: douta=16'ha4d3;
14648: douta=16'h9c93;
14649: douta=16'h8c32;
14650: douta=16'h8412;
14651: douta=16'h73b0;
14652: douta=16'h734f;
14653: douta=16'h6b4f;
14654: douta=16'h5aec;
14655: douta=16'h59e5;
14656: douta=16'hac2a;
14657: douta=16'hc4eb;
14658: douta=16'he5d2;
14659: douta=16'he653;
14660: douta=16'hee75;
14661: douta=16'hee74;
14662: douta=16'he613;
14663: douta=16'hee74;
14664: douta=16'he633;
14665: douta=16'hddd1;
14666: douta=16'hcd50;
14667: douta=16'hc4f0;
14668: douta=16'hb4b0;
14669: douta=16'h9c51;
14670: douta=16'h9452;
14671: douta=16'h8c73;
14672: douta=16'h8453;
14673: douta=16'h8c95;
14674: douta=16'h73f3;
14675: douta=16'h73d2;
14676: douta=16'h7413;
14677: douta=16'h6bf3;
14678: douta=16'h5370;
14679: douta=16'h5b72;
14680: douta=16'h4b10;
14681: douta=16'h4b31;
14682: douta=16'h31ea;
14683: douta=16'h42ae;
14684: douta=16'h0884;
14685: douta=16'h1926;
14686: douta=16'h0842;
14687: douta=16'h0862;
14688: douta=16'h1084;
14689: douta=16'h10a4;
14690: douta=16'h1905;
14691: douta=16'h1926;
14692: douta=16'h1905;
14693: douta=16'h1926;
14694: douta=16'h1905;
14695: douta=16'h0000;
14696: douta=16'h0000;
14697: douta=16'h0001;
14698: douta=16'h84b7;
14699: douta=16'h0021;
14700: douta=16'h10e5;
14701: douta=16'h1106;
14702: douta=16'h31c8;
14703: douta=16'h8bed;
14704: douta=16'h5248;
14705: douta=16'h946f;
14706: douta=16'had31;
14707: douta=16'h83ce;
14708: douta=16'h3a2a;
14709: douta=16'h5b92;
14710: douta=16'h9dba;
14711: douta=16'h9d9a;
14712: douta=16'h8d17;
14713: douta=16'h8d18;
14714: douta=16'h84f8;
14715: douta=16'h8d59;
14716: douta=16'h7cb7;
14717: douta=16'h7c97;
14718: douta=16'h8d39;
14719: douta=16'h9dbb;
14720: douta=16'h8d39;
14721: douta=16'h7476;
14722: douta=16'h84d7;
14723: douta=16'h7456;
14724: douta=16'h6c14;
14725: douta=16'h8d59;
14726: douta=16'h9dbb;
14727: douta=16'h84d8;
14728: douta=16'h9d9a;
14729: douta=16'h9dba;
14730: douta=16'h9d9a;
14731: douta=16'h7497;
14732: douta=16'h6c15;
14733: douta=16'h5392;
14734: douta=16'h8d39;
14735: douta=16'h8519;
14736: douta=16'h8518;
14737: douta=16'h9dbb;
14738: douta=16'h959a;
14739: douta=16'h959a;
14740: douta=16'h84f9;
14741: douta=16'h7cf9;
14742: douta=16'h8d39;
14743: douta=16'h95dd;
14744: douta=16'h7476;
14745: douta=16'h5b92;
14746: douta=16'h5207;
14747: douta=16'h72a9;
14748: douta=16'h6248;
14749: douta=16'h62ec;
14750: douta=16'h3a2c;
14751: douta=16'h224e;
14752: douta=16'h2a6f;
14753: douta=16'h4c17;
14754: douta=16'h5438;
14755: douta=16'h3b54;
14756: douta=16'h4b94;
14757: douta=16'h4bb4;
14758: douta=16'h5c58;
14759: douta=16'h53b6;
14760: douta=16'h4b95;
14761: douta=16'h6457;
14762: douta=16'h53f6;
14763: douta=16'h53b6;
14764: douta=16'h3b33;
14765: douta=16'h5c17;
14766: douta=16'h6b0c;
14767: douta=16'h6a65;
14768: douta=16'h3144;
14769: douta=16'h20a2;
14770: douta=16'h1926;
14771: douta=16'h5c58;
14772: douta=16'h649a;
14773: douta=16'h6bd0;
14774: douta=16'hbdd4;
14775: douta=16'hdeb7;
14776: douta=16'had52;
14777: douta=16'h5aa8;
14778: douta=16'h28c2;
14779: douta=16'h3944;
14780: douta=16'h3964;
14781: douta=16'h4164;
14782: douta=16'h3964;
14783: douta=16'h49a6;
14784: douta=16'h6390;
14785: douta=16'h3986;
14786: douta=16'h3965;
14787: douta=16'h2904;
14788: douta=16'h424b;
14789: douta=16'h2a4e;
14790: douta=16'h4353;
14791: douta=16'h4374;
14792: douta=16'h3ad1;
14793: douta=16'h6457;
14794: douta=16'h7476;
14795: douta=16'h6c15;
14796: douta=16'h63d3;
14797: douta=16'h8496;
14798: douta=16'h73f3;
14799: douta=16'h8c74;
14800: douta=16'h8433;
14801: douta=16'had77;
14802: douta=16'hc638;
14803: douta=16'he613;
14804: douta=16'hee95;
14805: douta=16'he676;
14806: douta=16'he696;
14807: douta=16'heed8;
14808: douta=16'heed8;
14809: douta=16'heed7;
14810: douta=16'hee96;
14811: douta=16'heeb7;
14812: douta=16'he634;
14813: douta=16'hde13;
14814: douta=16'hd5b2;
14815: douta=16'hbd31;
14816: douta=16'h8c10;
14817: douta=16'h7bd1;
14818: douta=16'h7bb0;
14819: douta=16'h7390;
14820: douta=16'h7bb0;
14821: douta=16'h6b0d;
14822: douta=16'h4985;
14823: douta=16'h8328;
14824: douta=16'hbcac;
14825: douta=16'hd570;
14826: douta=16'he634;
14827: douta=16'hee75;
14828: douta=16'he633;
14829: douta=16'hddb1;
14830: douta=16'he654;
14831: douta=16'hde13;
14832: douta=16'hd5b1;
14833: douta=16'hcd71;
14834: douta=16'hc530;
14835: douta=16'hbd11;
14836: douta=16'hb4f1;
14837: douta=16'ha4b2;
14838: douta=16'ha4b2;
14839: douta=16'h8c12;
14840: douta=16'h9472;
14841: douta=16'h8412;
14842: douta=16'h732e;
14843: douta=16'h7bb0;
14844: douta=16'h7bb0;
14845: douta=16'h4a28;
14846: douta=16'h7a87;
14847: douta=16'h9b8a;
14848: douta=16'hcd2d;
14849: douta=16'hddd1;
14850: douta=16'he654;
14851: douta=16'hee74;
14852: douta=16'hee74;
14853: douta=16'hee74;
14854: douta=16'he653;
14855: douta=16'he632;
14856: douta=16'hddd0;
14857: douta=16'hcd30;
14858: douta=16'hbd0f;
14859: douta=16'hb48f;
14860: douta=16'ha470;
14861: douta=16'h9451;
14862: douta=16'h8c11;
14863: douta=16'h8c32;
14864: douta=16'h8c94;
14865: douta=16'h8454;
14866: douta=16'h8474;
14867: douta=16'h8475;
14868: douta=16'h7c13;
14869: douta=16'h73f3;
14870: douta=16'h63b2;
14871: douta=16'h5b50;
14872: douta=16'h3a2c;
14873: douta=16'h7b2d;
14874: douta=16'h4ace;
14875: douta=16'h4ace;
14876: douta=16'h3a8d;
14877: douta=16'h2167;
14878: douta=16'h428d;
14879: douta=16'h4acf;
14880: douta=16'h0883;
14881: douta=16'h10c4;
14882: douta=16'h18e5;
14883: douta=16'h10e5;
14884: douta=16'h10c4;
14885: douta=16'h10c4;
14886: douta=16'h10e5;
14887: douta=16'h1926;
14888: douta=16'h1926;
14889: douta=16'h0000;
14890: douta=16'h0000;
14891: douta=16'h1905;
14892: douta=16'h2126;
14893: douta=16'h1946;
14894: douta=16'h1926;
14895: douta=16'h3a08;
14896: douta=16'hbd51;
14897: douta=16'had11;
14898: douta=16'h7bad;
14899: douta=16'h4248;
14900: douta=16'h62eb;
14901: douta=16'h9c8f;
14902: douta=16'h6b0b;
14903: douta=16'h4208;
14904: douta=16'h428d;
14905: douta=16'h5b51;
14906: douta=16'h7476;
14907: douta=16'h9559;
14908: douta=16'h8d39;
14909: douta=16'h8d18;
14910: douta=16'h8cf8;
14911: douta=16'h8d39;
14912: douta=16'h9559;
14913: douta=16'h8d18;
14914: douta=16'h7cb7;
14915: douta=16'h8d39;
14916: douta=16'h9dbb;
14917: douta=16'h7cb7;
14918: douta=16'h6c76;
14919: douta=16'h959a;
14920: douta=16'h7cb7;
14921: douta=16'h8d39;
14922: douta=16'h8d39;
14923: douta=16'h9559;
14924: douta=16'h84f8;
14925: douta=16'h9ddc;
14926: douta=16'h6435;
14927: douta=16'h5371;
14928: douta=16'h5b52;
14929: douta=16'h7cf8;
14930: douta=16'h8539;
14931: douta=16'h74b7;
14932: douta=16'h7cb7;
14933: douta=16'h7496;
14934: douta=16'h63b3;
14935: douta=16'h3a2d;
14936: douta=16'h4310;
14937: douta=16'h5bb4;
14938: douta=16'h4b11;
14939: douta=16'h62ed;
14940: douta=16'h72a8;
14941: douta=16'h6248;
14942: douta=16'h6248;
14943: douta=16'h5a8a;
14944: douta=16'h11cd;
14945: douta=16'h4395;
14946: douta=16'h2ab0;
14947: douta=16'h43d6;
14948: douta=16'h3b33;
14949: douta=16'h4bd6;
14950: douta=16'h4bb5;
14951: douta=16'h4374;
14952: douta=16'h4b75;
14953: douta=16'h6458;
14954: douta=16'h53d6;
14955: douta=16'h6479;
14956: douta=16'h7d7c;
14957: douta=16'h5c37;
14958: douta=16'h5c78;
14959: douta=16'h8348;
14960: douta=16'h51c4;
14961: douta=16'h3144;
14962: douta=16'h0000;
14963: douta=16'h08e5;
14964: douta=16'h94d3;
14965: douta=16'hde75;
14966: douta=16'had10;
14967: douta=16'h6b4a;
14968: douta=16'h30c2;
14969: douta=16'h3944;
14970: douta=16'h3944;
14971: douta=16'h4185;
14972: douta=16'h41a5;
14973: douta=16'h4985;
14974: douta=16'h41a5;
14975: douta=16'h49c7;
14976: douta=16'h5b0e;
14977: douta=16'h3966;
14978: douta=16'h3945;
14979: douta=16'h2904;
14980: douta=16'h4a6c;
14981: douta=16'h21ca;
14982: douta=16'h4b95;
14983: douta=16'h53d6;
14984: douta=16'h4333;
14985: douta=16'h5c16;
14986: douta=16'h7455;
14987: douta=16'h7c97;
14988: douta=16'h6bf4;
14989: douta=16'h7c75;
14990: douta=16'h73f4;
14991: douta=16'h94b5;
14992: douta=16'h8c74;
14993: douta=16'hbdd8;
14994: douta=16'hc618;
14995: douta=16'hbd13;
14996: douta=16'hee94;
14997: douta=16'he696;
14998: douta=16'he696;
14999: douta=16'heed8;
15000: douta=16'heed8;
15001: douta=16'heeb7;
15002: douta=16'heeb7;
15003: douta=16'hee96;
15004: douta=16'he634;
15005: douta=16'hd5f3;
15006: douta=16'hcdb2;
15007: douta=16'ha4b1;
15008: douta=16'h9c71;
15009: douta=16'h83f1;
15010: douta=16'h738f;
15011: douta=16'h736f;
15012: douta=16'h6b4e;
15013: douta=16'h41c7;
15014: douta=16'h8b29;
15015: douta=16'hb48c;
15016: douta=16'hcd2e;
15017: douta=16'hde12;
15018: douta=16'he675;
15019: douta=16'he675;
15020: douta=16'he695;
15021: douta=16'he612;
15022: douta=16'he674;
15023: douta=16'hddb1;
15024: douta=16'hd591;
15025: douta=16'hcd50;
15026: douta=16'hc530;
15027: douta=16'hacb1;
15028: douta=16'hb4d2;
15029: douta=16'hacb2;
15030: douta=16'ha493;
15031: douta=16'h8c12;
15032: douta=16'h8c11;
15033: douta=16'h8c12;
15034: douta=16'h734e;
15035: douta=16'h730e;
15036: douta=16'h6b6f;
15037: douta=16'h4963;
15038: douta=16'habeb;
15039: douta=16'hac4a;
15040: douta=16'hdd8f;
15041: douta=16'he653;
15042: douta=16'hee95;
15043: douta=16'he674;
15044: douta=16'hee54;
15045: douta=16'hee74;
15046: douta=16'he653;
15047: douta=16'hddf2;
15048: douta=16'hd58f;
15049: douta=16'hbccf;
15050: douta=16'hb4af;
15051: douta=16'ha430;
15052: douta=16'h9c51;
15053: douta=16'h9452;
15054: douta=16'h8c32;
15055: douta=16'h8c33;
15056: douta=16'h8432;
15057: douta=16'h8453;
15058: douta=16'h8453;
15059: douta=16'h7bf3;
15060: douta=16'h7c13;
15061: douta=16'h6bd2;
15062: douta=16'h5b0e;
15063: douta=16'h52ae;
15064: douta=16'h9329;
15065: douta=16'he5b2;
15066: douta=16'h5351;
15067: douta=16'h4ace;
15068: douta=16'h3aad;
15069: douta=16'h1948;
15070: douta=16'h0884;
15071: douta=16'h2989;
15072: douta=16'h4aae;
15073: douta=16'h0883;
15074: douta=16'h10e5;
15075: douta=16'h10e5;
15076: douta=16'h10e5;
15077: douta=16'h10e5;
15078: douta=16'h10e5;
15079: douta=16'h10e5;
15080: douta=16'h1906;
15081: douta=16'h10c4;
15082: douta=16'h0000;
15083: douta=16'h0042;
15084: douta=16'h0883;
15085: douta=16'h2167;
15086: douta=16'h1947;
15087: douta=16'h08a5;
15088: douta=16'h738e;
15089: douta=16'h732b;
15090: douta=16'h3186;
15091: douta=16'hb512;
15092: douta=16'h2124;
15093: douta=16'ha4b0;
15094: douta=16'h5aa9;
15095: douta=16'h41e8;
15096: douta=16'h8bcd;
15097: douta=16'h4207;
15098: douta=16'h528b;
15099: douta=16'h5aed;
15100: douta=16'h5b92;
15101: douta=16'h7476;
15102: douta=16'h7cd7;
15103: douta=16'h959a;
15104: douta=16'h8d39;
15105: douta=16'h9559;
15106: douta=16'h957a;
15107: douta=16'h8518;
15108: douta=16'h8518;
15109: douta=16'h84d7;
15110: douta=16'h8538;
15111: douta=16'h8d18;
15112: douta=16'h8d59;
15113: douta=16'h7cd7;
15114: douta=16'h8d18;
15115: douta=16'h8519;
15116: douta=16'h9dfc;
15117: douta=16'ha63d;
15118: douta=16'hae7e;
15119: douta=16'ha65e;
15120: douta=16'h4b73;
15121: douta=16'h10e6;
15122: douta=16'h634f;
15123: douta=16'h3a2b;
15124: douta=16'h3a4c;
15125: douta=16'h2189;
15126: douta=16'h29ca;
15127: douta=16'h4b51;
15128: douta=16'h3a8e;
15129: douta=16'h3aaf;
15130: douta=16'h4b51;
15131: douta=16'h5bb3;
15132: douta=16'h734d;
15133: douta=16'h6aa9;
15134: douta=16'h6a89;
15135: douta=16'h6248;
15136: douta=16'h320b;
15137: douta=16'h118a;
15138: douta=16'h21ed;
15139: douta=16'h3333;
15140: douta=16'h32d2;
15141: douta=16'h2af2;
15142: douta=16'h3b12;
15143: douta=16'h4bb5;
15144: douta=16'h5417;
15145: douta=16'h5c17;
15146: douta=16'h6cb9;
15147: douta=16'h4374;
15148: douta=16'h7d7c;
15149: douta=16'h53f6;
15150: douta=16'h7dbf;
15151: douta=16'h8b69;
15152: douta=16'h6245;
15153: douta=16'h4164;
15154: douta=16'h2146;
15155: douta=16'h73ef;
15156: douta=16'hce13;
15157: douta=16'had2e;
15158: douta=16'h41a6;
15159: douta=16'h3923;
15160: douta=16'h3944;
15161: douta=16'h41a5;
15162: douta=16'h4185;
15163: douta=16'h49a6;
15164: douta=16'h49a6;
15165: douta=16'h41a6;
15166: douta=16'h41a7;
15167: douta=16'h4186;
15168: douta=16'h4144;
15169: douta=16'h3904;
15170: douta=16'h3965;
15171: douta=16'h2924;
15172: douta=16'h4a8d;
15173: douta=16'h42ce;
15174: douta=16'h2168;
15175: douta=16'h19eb;
15176: douta=16'h220d;
15177: douta=16'h4353;
15178: douta=16'h6c36;
15179: douta=16'h6c15;
15180: douta=16'h7cd8;
15181: douta=16'h7414;
15182: douta=16'h8cd7;
15183: douta=16'h94f6;
15184: douta=16'hb597;
15185: douta=16'h9cd5;
15186: douta=16'hc5f8;
15187: douta=16'h9492;
15188: douta=16'h7bf1;
15189: douta=16'he614;
15190: douta=16'he6b7;
15191: douta=16'heeb7;
15192: douta=16'heed7;
15193: douta=16'hee96;
15194: douta=16'he675;
15195: douta=16'he675;
15196: douta=16'hd5d3;
15197: douta=16'hc571;
15198: douta=16'hb4f1;
15199: douta=16'h8c31;
15200: douta=16'h8c11;
15201: douta=16'h83f1;
15202: douta=16'h6b0e;
15203: douta=16'h62ed;
15204: douta=16'h3945;
15205: douta=16'ha46c;
15206: douta=16'hac6c;
15207: douta=16'hbcee;
15208: douta=16'he655;
15209: douta=16'he634;
15210: douta=16'hee96;
15211: douta=16'he695;
15212: douta=16'he655;
15213: douta=16'hbcef;
15214: douta=16'hd550;
15215: douta=16'hcd50;
15216: douta=16'hbcd1;
15217: douta=16'hacd1;
15218: douta=16'ha4b1;
15219: douta=16'ha471;
15220: douta=16'h9452;
15221: douta=16'h83f1;
15222: douta=16'h7bd1;
15223: douta=16'h738f;
15224: douta=16'h734f;
15225: douta=16'h6b2d;
15226: douta=16'h62cd;
15227: douta=16'h4985;
15228: douta=16'h82e9;
15229: douta=16'hb48b;
15230: douta=16'hd54f;
15231: douta=16'heeb6;
15232: douta=16'heeb7;
15233: douta=16'heeb7;
15234: douta=16'hee95;
15235: douta=16'hee74;
15236: douta=16'he654;
15237: douta=16'he653;
15238: douta=16'hddb1;
15239: douta=16'hd530;
15240: douta=16'hb4d0;
15241: douta=16'ha472;
15242: douta=16'h9c71;
15243: douta=16'h9c52;
15244: douta=16'h9452;
15245: douta=16'h9432;
15246: douta=16'h8c32;
15247: douta=16'h7bd0;
15248: douta=16'h738f;
15249: douta=16'h7b90;
15250: douta=16'h73b0;
15251: douta=16'h734f;
15252: douta=16'h734f;
15253: douta=16'h5a6b;
15254: douta=16'h7a87;
15255: douta=16'hddd1;
15256: douta=16'hd5d2;
15257: douta=16'he614;
15258: douta=16'h9472;
15259: douta=16'h6b90;
15260: douta=16'h73f2;
15261: douta=16'h5b71;
15262: douta=16'h29cb;
15263: douta=16'h29eb;
15264: douta=16'h2147;
15265: douta=16'h0884;
15266: douta=16'h3a6d;
15267: douta=16'h326d;
15268: douta=16'h1083;
15269: douta=16'h18c5;
15270: douta=16'h1905;
15271: douta=16'h1926;
15272: douta=16'h1926;
15273: douta=16'h18e5;
15274: douta=16'h1926;
15275: douta=16'h2127;
15276: douta=16'h2146;
15277: douta=16'h0042;
15278: douta=16'h0001;
15279: douta=16'h0001;
15280: douta=16'h31c8;
15281: douta=16'h5bb3;
15282: douta=16'h5b93;
15283: douta=16'h0000;
15284: douta=16'h1106;
15285: douta=16'h73ad;
15286: douta=16'h9cb1;
15287: douta=16'h630b;
15288: douta=16'h5269;
15289: douta=16'h944f;
15290: douta=16'h2126;
15291: douta=16'h7bce;
15292: douta=16'h31a8;
15293: douta=16'h5aec;
15294: douta=16'h6b2d;
15295: douta=16'ha4d1;
15296: douta=16'h83ef;
15297: douta=16'h630c;
15298: douta=16'h7b8d;
15299: douta=16'h5acb;
15300: douta=16'h3187;
15301: douta=16'h39e7;
15302: douta=16'h31a6;
15303: douta=16'h5289;
15304: douta=16'h3186;
15305: douta=16'h20e4;
15306: douta=16'h1041;
15307: douta=16'h41e7;
15308: douta=16'h83ef;
15309: douta=16'hd54f;
15310: douta=16'hac0a;
15311: douta=16'hac2a;
15312: douta=16'ha3ca;
15313: douta=16'h2a4e;
15314: douta=16'h21a9;
15315: douta=16'h3a4c;
15316: douta=16'h4aad;
15317: douta=16'h4b0f;
15318: douta=16'h3a6d;
15319: douta=16'h530f;
15320: douta=16'h326e;
15321: douta=16'h328f;
15322: douta=16'h63d3;
15323: douta=16'h21ec;
15324: douta=16'h63b2;
15325: douta=16'h4310;
15326: douta=16'h6391;
15327: douta=16'h72eb;
15328: douta=16'h6289;
15329: douta=16'h5a48;
15330: douta=16'h6268;
15331: douta=16'h11cd;
15332: douta=16'h21ec;
15333: douta=16'h3333;
15334: douta=16'h5c7a;
15335: douta=16'h1a2e;
15336: douta=16'h3b54;
15337: douta=16'h6478;
15338: douta=16'h53f6;
15339: douta=16'h5c37;
15340: douta=16'h753b;
15341: douta=16'h6498;
15342: douta=16'h4b95;
15343: douta=16'h62aa;
15344: douta=16'h7aca;
15345: douta=16'h52aa;
15346: douta=16'h83cc;
15347: douta=16'h4985;
15348: douta=16'h28c2;
15349: douta=16'h4164;
15350: douta=16'h4164;
15351: douta=16'h4185;
15352: douta=16'h41a6;
15353: douta=16'h49e7;
15354: douta=16'h4a08;
15355: douta=16'h3966;
15356: douta=16'h39a6;
15357: douta=16'h41c7;
15358: douta=16'h41c7;
15359: douta=16'h39a6;
15360: douta=16'h3944;
15361: douta=16'h41a7;
15362: douta=16'h3945;
15363: douta=16'h3145;
15364: douta=16'h320a;
15365: douta=16'h4acf;
15366: douta=16'h21a9;
15367: douta=16'h3b12;
15368: douta=16'h3ad1;
15369: douta=16'h53b4;
15370: douta=16'h5373;
15371: douta=16'h5373;
15372: douta=16'h63f4;
15373: douta=16'h8518;
15374: douta=16'h4aef;
15375: douta=16'h5b30;
15376: douta=16'h6bd2;
15377: douta=16'h8411;
15378: douta=16'hadd9;
15379: douta=16'hce19;
15380: douta=16'hb5b7;
15381: douta=16'hde78;
15382: douta=16'he675;
15383: douta=16'hee96;
15384: douta=16'heeb7;
15385: douta=16'he696;
15386: douta=16'he675;
15387: douta=16'he634;
15388: douta=16'hcd72;
15389: douta=16'hc531;
15390: douta=16'hacd1;
15391: douta=16'h8c11;
15392: douta=16'h7b70;
15393: douta=16'h736e;
15394: douta=16'h526a;
15395: douta=16'h2904;
15396: douta=16'ha3eb;
15397: douta=16'hbc8d;
15398: douta=16'hd570;
15399: douta=16'hddd2;
15400: douta=16'he675;
15401: douta=16'he655;
15402: douta=16'hd591;
15403: douta=16'hee96;
15404: douta=16'hee75;
15405: douta=16'hee74;
15406: douta=16'h83ef;
15407: douta=16'ha491;
15408: douta=16'hb4b1;
15409: douta=16'h9431;
15410: douta=16'h9432;
15411: douta=16'h83f1;
15412: douta=16'h83d1;
15413: douta=16'h7bd1;
15414: douta=16'h83f1;
15415: douta=16'h736e;
15416: douta=16'h736f;
15417: douta=16'h630e;
15418: douta=16'h6a46;
15419: douta=16'ha40a;
15420: douta=16'hac0c;
15421: douta=16'hd590;
15422: douta=16'hee75;
15423: douta=16'hf6d7;
15424: douta=16'hf6b6;
15425: douta=16'hf6b6;
15426: douta=16'hee95;
15427: douta=16'he674;
15428: douta=16'hddd2;
15429: douta=16'hd590;
15430: douta=16'hb4d0;
15431: douta=16'hb4d1;
15432: douta=16'h9c72;
15433: douta=16'hacb2;
15434: douta=16'h9c72;
15435: douta=16'h9432;
15436: douta=16'h8c32;
15437: douta=16'h83f1;
15438: douta=16'h7bd1;
15439: douta=16'h83d1;
15440: douta=16'h7bb0;
15441: douta=16'h6b2d;
15442: douta=16'h732d;
15443: douta=16'h62cd;
15444: douta=16'h49e8;
15445: douta=16'hbc4b;
15446: douta=16'hddb0;
15447: douta=16'hddf3;
15448: douta=16'hd5b2;
15449: douta=16'hddb2;
15450: douta=16'h9c92;
15451: douta=16'h6bf3;
15452: douta=16'h6bd2;
15453: douta=16'h6bd2;
15454: douta=16'h42af;
15455: douta=16'h3a8e;
15456: douta=16'h3aae;
15457: douta=16'h21ec;
15458: douta=16'h2168;
15459: douta=16'h10a4;
15460: douta=16'h3a8e;
15461: douta=16'h2168;
15462: douta=16'h10c3;
15463: douta=16'h18e5;
15464: douta=16'h18e6;
15465: douta=16'h10e5;
15466: douta=16'h1906;
15467: douta=16'h1084;
15468: douta=16'h1083;
15469: douta=16'h1926;
15470: douta=16'h1926;
15471: douta=16'h2147;
15472: douta=16'h0000;
15473: douta=16'h0000;
15474: douta=16'h0000;
15475: douta=16'h10c4;
15476: douta=16'h2126;
15477: douta=16'h1926;
15478: douta=16'h0063;
15479: douta=16'h7bef;
15480: douta=16'h8c2f;
15481: douta=16'h31c8;
15482: douta=16'hde77;
15483: douta=16'had12;
15484: douta=16'h840f;
15485: douta=16'h2986;
15486: douta=16'h630b;
15487: douta=16'h6b2c;
15488: douta=16'ha4d2;
15489: douta=16'h4208;
15490: douta=16'h6b6d;
15491: douta=16'h52cb;
15492: douta=16'h8c4f;
15493: douta=16'h31a7;
15494: douta=16'h5acb;
15495: douta=16'h632c;
15496: douta=16'h39a6;
15497: douta=16'h39c7;
15498: douta=16'h62cb;
15499: douta=16'hc56f;
15500: douta=16'h9348;
15501: douta=16'ha3ea;
15502: douta=16'h6aca;
15503: douta=16'h31c9;
15504: douta=16'h2a2d;
15505: douta=16'h322b;
15506: douta=16'h42ae;
15507: douta=16'h3a6d;
15508: douta=16'h42ad;
15509: douta=16'h42ae;
15510: douta=16'h3a6c;
15511: douta=16'h3aae;
15512: douta=16'h6370;
15513: douta=16'h73f2;
15514: douta=16'h326d;
15515: douta=16'h5b91;
15516: douta=16'h42f0;
15517: douta=16'h5351;
15518: douta=16'h5b71;
15519: douta=16'h2a6f;
15520: douta=16'h5aaa;
15521: douta=16'h5a48;
15522: douta=16'h5a88;
15523: douta=16'h6289;
15524: douta=16'h4a8d;
15525: douta=16'h19ac;
15526: douta=16'h2b13;
15527: douta=16'h3334;
15528: douta=16'h3b75;
15529: douta=16'h3b12;
15530: douta=16'h4bd5;
15531: douta=16'h6cfa;
15532: douta=16'h4373;
15533: douta=16'h3af1;
15534: douta=16'h4bf8;
15535: douta=16'h7c51;
15536: douta=16'hb573;
15537: douta=16'h836c;
15538: douta=16'h4164;
15539: douta=16'h4985;
15540: douta=16'h4985;
15541: douta=16'h49a6;
15542: douta=16'h41a6;
15543: douta=16'h49c6;
15544: douta=16'h4166;
15545: douta=16'h49e7;
15546: douta=16'h39a6;
15547: douta=16'h41a7;
15548: douta=16'h41c7;
15549: douta=16'h41a7;
15550: douta=16'h41a7;
15551: douta=16'h41a7;
15552: douta=16'h4185;
15553: douta=16'h526b;
15554: douta=16'h3945;
15555: douta=16'h3124;
15556: douta=16'h320a;
15557: douta=16'h5b51;
15558: douta=16'h322b;
15559: douta=16'h4353;
15560: douta=16'h2a0e;
15561: douta=16'h53d4;
15562: douta=16'h6c77;
15563: douta=16'h5bf5;
15564: douta=16'h8539;
15565: douta=16'h7c55;
15566: douta=16'h9d59;
15567: douta=16'h8cd6;
15568: douta=16'h8495;
15569: douta=16'h630d;
15570: douta=16'hadfa;
15571: douta=16'hb597;
15572: douta=16'hc65a;
15573: douta=16'h83f0;
15574: douta=16'hee75;
15575: douta=16'he676;
15576: douta=16'hee96;
15577: douta=16'he675;
15578: douta=16'he675;
15579: douta=16'hde15;
15580: douta=16'hc552;
15581: douta=16'hacb1;
15582: douta=16'ha471;
15583: douta=16'h83d0;
15584: douta=16'h7b90;
15585: douta=16'h7b6f;
15586: douta=16'h2903;
15587: douta=16'h6a87;
15588: douta=16'ha46b;
15589: douta=16'hc52f;
15590: douta=16'hddf2;
15591: douta=16'he634;
15592: douta=16'he675;
15593: douta=16'hee95;
15594: douta=16'hcd2f;
15595: douta=16'hee75;
15596: douta=16'he675;
15597: douta=16'he654;
15598: douta=16'h7bae;
15599: douta=16'h7390;
15600: douta=16'h9c72;
15601: douta=16'h9431;
15602: douta=16'h8c31;
15603: douta=16'h8bf1;
15604: douta=16'h7bf1;
15605: douta=16'h7bd0;
15606: douta=16'h7bd1;
15607: douta=16'h7bb0;
15608: douta=16'h73b0;
15609: douta=16'h20c3;
15610: douta=16'h9bab;
15611: douta=16'hbc8c;
15612: douta=16'hcd0e;
15613: douta=16'he633;
15614: douta=16'hee96;
15615: douta=16'heeb7;
15616: douta=16'hee96;
15617: douta=16'hee75;
15618: douta=16'hee95;
15619: douta=16'hddd2;
15620: douta=16'hd591;
15621: douta=16'hc531;
15622: douta=16'h9c72;
15623: douta=16'ha492;
15624: douta=16'h9c93;
15625: douta=16'h9c93;
15626: douta=16'ha4b4;
15627: douta=16'h8c32;
15628: douta=16'h8412;
15629: douta=16'h7bd1;
15630: douta=16'h7bb0;
15631: douta=16'h7b6f;
15632: douta=16'h7b8f;
15633: douta=16'h736e;
15634: douta=16'h6aec;
15635: douta=16'h832b;
15636: douta=16'h82e9;
15637: douta=16'hdd90;
15638: douta=16'hee74;
15639: douta=16'he634;
15640: douta=16'hd5d3;
15641: douta=16'hc532;
15642: douta=16'h9472;
15643: douta=16'h7413;
15644: douta=16'h73f3;
15645: douta=16'h6bd2;
15646: douta=16'h5330;
15647: douta=16'h5351;
15648: douta=16'h42d0;
15649: douta=16'h324d;
15650: douta=16'h29eb;
15651: douta=16'h21a9;
15652: douta=16'h10c4;
15653: douta=16'h4af0;
15654: douta=16'h1906;
15655: douta=16'h1105;
15656: douta=16'h10e5;
15657: douta=16'h1926;
15658: douta=16'h10e5;
15659: douta=16'h10a4;
15660: douta=16'h10e6;
15661: douta=16'h2168;
15662: douta=16'h1948;
15663: douta=16'h2168;
15664: douta=16'h1926;
15665: douta=16'h0883;
15666: douta=16'h0000;
15667: douta=16'h0883;
15668: douta=16'h1106;
15669: douta=16'h1926;
15670: douta=16'h08a3;
15671: douta=16'h424d;
15672: douta=16'h8474;
15673: douta=16'h3a09;
15674: douta=16'h4a49;
15675: douta=16'h7b8d;
15676: douta=16'hacf2;
15677: douta=16'h738e;
15678: douta=16'h31c7;
15679: douta=16'h6b4c;
15680: douta=16'h8c2e;
15681: douta=16'h9cb1;
15682: douta=16'h52ab;
15683: douta=16'h5aab;
15684: douta=16'h6b6c;
15685: douta=16'h4a8a;
15686: douta=16'h4229;
15687: douta=16'h31a6;
15688: douta=16'h41e7;
15689: douta=16'h734b;
15690: douta=16'hbd30;
15691: douta=16'h9368;
15692: douta=16'ha3eb;
15693: douta=16'ha40b;
15694: douta=16'h1969;
15695: douta=16'h322c;
15696: douta=16'h530f;
15697: douta=16'h4aee;
15698: douta=16'h530f;
15699: douta=16'h2a0b;
15700: douta=16'h4ace;
15701: douta=16'h19aa;
15702: douta=16'h5b50;
15703: douta=16'h2a2b;
15704: douta=16'h530f;
15705: douta=16'h6b91;
15706: douta=16'h3a8e;
15707: douta=16'h5b71;
15708: douta=16'h3aaf;
15709: douta=16'h42d0;
15710: douta=16'h6c14;
15711: douta=16'h2a2c;
15712: douta=16'h5b92;
15713: douta=16'h6269;
15714: douta=16'h6227;
15715: douta=16'h5228;
15716: douta=16'h5a69;
15717: douta=16'h42af;
15718: douta=16'h3334;
15719: douta=16'h4c18;
15720: douta=16'h3b54;
15721: douta=16'h4bf7;
15722: douta=16'h4bf6;
15723: douta=16'h5c37;
15724: douta=16'h4332;
15725: douta=16'h4333;
15726: douta=16'h5418;
15727: douta=16'h944f;
15728: douta=16'h51e6;
15729: douta=16'h2060;
15730: douta=16'h49a5;
15731: douta=16'h49c6;
15732: douta=16'h49a6;
15733: douta=16'h49c6;
15734: douta=16'h49c7;
15735: douta=16'h49c8;
15736: douta=16'h49c7;
15737: douta=16'h49e7;
15738: douta=16'h41c7;
15739: douta=16'h41a7;
15740: douta=16'h41a6;
15741: douta=16'h49e7;
15742: douta=16'h49c7;
15743: douta=16'h3146;
15744: douta=16'h41a6;
15745: douta=16'h6391;
15746: douta=16'h3965;
15747: douta=16'h3124;
15748: douta=16'h2146;
15749: douta=16'h63d3;
15750: douta=16'h19a9;
15751: douta=16'h5394;
15752: douta=16'h6416;
15753: douta=16'h4b11;
15754: douta=16'h5393;
15755: douta=16'h4b11;
15756: douta=16'h7cb7;
15757: douta=16'h6bf4;
15758: douta=16'h9517;
15759: douta=16'h9517;
15760: douta=16'h8475;
15761: douta=16'h9d16;
15762: douta=16'had57;
15763: douta=16'hbdf9;
15764: douta=16'hb5b8;
15765: douta=16'ha4d4;
15766: douta=16'had57;
15767: douta=16'hd5f3;
15768: douta=16'he654;
15769: douta=16'hde55;
15770: douta=16'hd614;
15771: douta=16'hcd93;
15772: douta=16'hb4f3;
15773: douta=16'h9472;
15774: douta=16'h8c31;
15775: douta=16'h7b8f;
15776: douta=16'h6b4f;
15777: douta=16'h3124;
15778: douta=16'h9c4d;
15779: douta=16'hb48e;
15780: douta=16'hd5b1;
15781: douta=16'hde13;
15782: douta=16'he633;
15783: douta=16'hee75;
15784: douta=16'he675;
15785: douta=16'he655;
15786: douta=16'he614;
15787: douta=16'hcd50;
15788: douta=16'he614;
15789: douta=16'hde14;
15790: douta=16'hacd0;
15791: douta=16'h9471;
15792: douta=16'h8433;
15793: douta=16'h5b2f;
15794: douta=16'h52ee;
15795: douta=16'h7390;
15796: douta=16'h7bf1;
15797: douta=16'h8c11;
15798: douta=16'h7bd0;
15799: douta=16'h38e2;
15800: douta=16'h82c6;
15801: douta=16'hb44a;
15802: douta=16'he5b0;
15803: douta=16'hee75;
15804: douta=16'hee95;
15805: douta=16'heeb7;
15806: douta=16'hee96;
15807: douta=16'he655;
15808: douta=16'he654;
15809: douta=16'he654;
15810: douta=16'hddf3;
15811: douta=16'hc512;
15812: douta=16'hc532;
15813: douta=16'hcd52;
15814: douta=16'h9c92;
15815: douta=16'h8c53;
15816: douta=16'h8412;
15817: douta=16'h83f1;
15818: douta=16'h8412;
15819: douta=16'h8c32;
15820: douta=16'h83b0;
15821: douta=16'h7baf;
15822: douta=16'h7b4e;
15823: douta=16'h6b0d;
15824: douta=16'h628b;
15825: douta=16'hb46b;
15826: douta=16'he5f2;
15827: douta=16'hd5d2;
15828: douta=16'hee95;
15829: douta=16'hee75;
15830: douta=16'he654;
15831: douta=16'hddf3;
15832: douta=16'hbd11;
15833: douta=16'ha492;
15834: douta=16'h9c93;
15835: douta=16'h8c74;
15836: douta=16'h7c54;
15837: douta=16'h7433;
15838: douta=16'h6bf4;
15839: douta=16'h63d3;
15840: douta=16'h5b93;
15841: douta=16'h4b31;
15842: douta=16'h3ad0;
15843: douta=16'h42f0;
15844: douta=16'h3a6e;
15845: douta=16'h29ea;
15846: douta=16'h10e7;
15847: douta=16'h4b10;
15848: douta=16'h4b31;
15849: douta=16'h1969;
15850: douta=16'h2189;
15851: douta=16'h1926;
15852: douta=16'h1906;
15853: douta=16'h1105;
15854: douta=16'h1905;
15855: douta=16'h1106;
15856: douta=16'h29a9;
15857: douta=16'h1946;
15858: douta=16'h1926;
15859: douta=16'h1926;
15860: douta=16'h2127;
15861: douta=16'h10a4;
15862: douta=16'h0042;
15863: douta=16'h0000;
15864: douta=16'h1063;
15865: douta=16'h7413;
15866: douta=16'h0021;
15867: douta=16'h2127;
15868: douta=16'h1927;
15869: douta=16'h08a5;
15870: douta=16'h73d1;
15871: douta=16'h39e8;
15872: douta=16'h7bae;
15873: douta=16'h4a68;
15874: douta=16'h6b6c;
15875: douta=16'h31e8;
15876: douta=16'h2986;
15877: douta=16'h0042;
15878: douta=16'h0083;
15879: douta=16'h72ea;
15880: douta=16'ha3aa;
15881: douta=16'habeb;
15882: douta=16'hb44b;
15883: douta=16'h5249;
15884: douta=16'h21aa;
15885: douta=16'h1106;
15886: douta=16'h52cc;
15887: douta=16'h4acd;
15888: douta=16'h52ee;
15889: douta=16'h42cf;
15890: douta=16'h634f;
15891: douta=16'h4aad;
15892: douta=16'h4acf;
15893: douta=16'h322c;
15894: douta=16'h326c;
15895: douta=16'h530f;
15896: douta=16'h4ace;
15897: douta=16'h4ace;
15898: douta=16'h3a8d;
15899: douta=16'h31eb;
15900: douta=16'h63b1;
15901: douta=16'h3acf;
15902: douta=16'h3aaf;
15903: douta=16'h4b31;
15904: douta=16'h5350;
15905: douta=16'h4b30;
15906: douta=16'h430f;
15907: douta=16'h5a8b;
15908: douta=16'h51e7;
15909: douta=16'h4a08;
15910: douta=16'h5228;
15911: douta=16'h42cf;
15912: douta=16'h19ab;
15913: douta=16'h4c18;
15914: douta=16'h32f2;
15915: douta=16'h3b33;
15916: douta=16'h7c32;
15917: douta=16'h730a;
15918: douta=16'h30c2;
15919: douta=16'h4985;
15920: douta=16'h49c6;
15921: douta=16'h49a5;
15922: douta=16'h51e8;
15923: douta=16'h5a29;
15924: douta=16'h4a08;
15925: douta=16'h5229;
15926: douta=16'h41a7;
15927: douta=16'h41a7;
15928: douta=16'h41a6;
15929: douta=16'h41a7;
15930: douta=16'h49c7;
15931: douta=16'h41a7;
15932: douta=16'h41c7;
15933: douta=16'h3986;
15934: douta=16'h41a7;
15935: douta=16'h41a7;
15936: douta=16'h41a5;
15937: douta=16'h6390;
15938: douta=16'h3103;
15939: douta=16'h3145;
15940: douta=16'h2945;
15941: douta=16'h31a9;
15942: douta=16'h328e;
15943: douta=16'h2168;
15944: douta=16'h3a2c;
15945: douta=16'h4acf;
15946: douta=16'h8c31;
15947: douta=16'h9cb4;
15948: douta=16'h8d39;
15949: douta=16'ha537;
15950: douta=16'hadb9;
15951: douta=16'h94f6;
15952: douta=16'h94f5;
15953: douta=16'h94d5;
15954: douta=16'hc5d7;
15955: douta=16'hc619;
15956: douta=16'h8431;
15957: douta=16'h5b0e;
15958: douta=16'had97;
15959: douta=16'hde79;
15960: douta=16'hd69a;
15961: douta=16'hde34;
15962: douta=16'hd5f3;
15963: douta=16'hc551;
15964: douta=16'h9451;
15965: douta=16'h8c11;
15966: douta=16'h7bb0;
15967: douta=16'h632f;
15968: douta=16'h28e3;
15969: douta=16'hb48d;
15970: douta=16'hc54f;
15971: douta=16'hd5b0;
15972: douta=16'he634;
15973: douta=16'he675;
15974: douta=16'hee75;
15975: douta=16'hddd2;
15976: douta=16'he654;
15977: douta=16'he654;
15978: douta=16'hde13;
15979: douta=16'hd5b2;
15980: douta=16'hc550;
15981: douta=16'hc531;
15982: douta=16'hbd12;
15983: douta=16'h9c92;
15984: douta=16'h8452;
15985: douta=16'h73b1;
15986: douta=16'h632f;
15987: douta=16'h632f;
15988: douta=16'h5ace;
15989: douta=16'h4aae;
15990: douta=16'h2947;
15991: douta=16'ha389;
15992: douta=16'he590;
15993: douta=16'he633;
15994: douta=16'heeb7;
15995: douta=16'hee96;
15996: douta=16'hf6d7;
15997: douta=16'he675;
15998: douta=16'heeb6;
15999: douta=16'he634;
16000: douta=16'hd5d3;
16001: douta=16'hcdb3;
16002: douta=16'hbd32;
16003: douta=16'hacb2;
16004: douta=16'h9452;
16005: douta=16'h9473;
16006: douta=16'h8c33;
16007: douta=16'h8432;
16008: douta=16'h7bb0;
16009: douta=16'h7b8f;
16010: douta=16'h736e;
16011: douta=16'h732d;
16012: douta=16'h72ec;
16013: douta=16'h732d;
16014: douta=16'h7b4d;
16015: douta=16'h936a;
16016: douta=16'hb44b;
16017: douta=16'ha3e9;
16018: douta=16'hb46b;
16019: douta=16'hcd0e;
16020: douta=16'hd590;
16021: douta=16'hddd2;
16022: douta=16'hcd92;
16023: douta=16'hcd32;
16024: douta=16'hac91;
16025: douta=16'ha492;
16026: douta=16'h9473;
16027: douta=16'h8cb5;
16028: douta=16'h7413;
16029: douta=16'h7413;
16030: douta=16'h6bf3;
16031: douta=16'h7413;
16032: douta=16'h6c14;
16033: douta=16'h63d4;
16034: douta=16'h5bd4;
16035: douta=16'h4b52;
16036: douta=16'h324d;
16037: douta=16'h29cb;
16038: douta=16'h320c;
16039: douta=16'h2189;
16040: douta=16'h08c5;
16041: douta=16'h320b;
16042: douta=16'h21a9;
16043: douta=16'h1106;
16044: douta=16'h0884;
16045: douta=16'h10e5;
16046: douta=16'h10e5;
16047: douta=16'h10c5;
16048: douta=16'h10e5;
16049: douta=16'h10e5;
16050: douta=16'h10e5;
16051: douta=16'h2147;
16052: douta=16'h1927;
16053: douta=16'h1947;
16054: douta=16'h1926;
16055: douta=16'h1927;
16056: douta=16'h1947;
16057: douta=16'h0000;
16058: douta=16'h0062;
16059: douta=16'h0062;
16060: douta=16'h1906;
16061: douta=16'h10e5;
16062: douta=16'h7c74;
16063: douta=16'h84b6;
16064: douta=16'h6c14;
16065: douta=16'h6393;
16066: douta=16'h1906;
16067: douta=16'h1905;
16068: douta=16'h18e5;
16069: douta=16'hc50f;
16070: douta=16'hd50d;
16071: douta=16'hb42b;
16072: douta=16'hb44b;
16073: douta=16'h4a4a;
16074: douta=16'h0086;
16075: douta=16'h634d;
16076: douta=16'h2168;
16077: douta=16'h3209;
16078: douta=16'h2188;
16079: douta=16'h4a8c;
16080: douta=16'h52ac;
16081: douta=16'h29ca;
16082: douta=16'h320b;
16083: douta=16'h52ee;
16084: douta=16'h42ae;
16085: douta=16'h4b10;
16086: douta=16'h29aa;
16087: douta=16'h4ace;
16088: douta=16'h4b0f;
16089: douta=16'h634f;
16090: douta=16'h3a4c;
16091: douta=16'h530f;
16092: douta=16'h428d;
16093: douta=16'h322d;
16094: douta=16'h5372;
16095: douta=16'h328e;
16096: douta=16'h4b51;
16097: douta=16'h42f0;
16098: douta=16'h4b0f;
16099: douta=16'h21a9;
16100: douta=16'h3a6c;
16101: douta=16'h41c7;
16102: douta=16'h4a08;
16103: douta=16'h49c7;
16104: douta=16'h5209;
16105: douta=16'h328f;
16106: douta=16'h32f2;
16107: douta=16'h3a4b;
16108: douta=16'h3922;
16109: douta=16'h4185;
16110: douta=16'h51c5;
16111: douta=16'h49a6;
16112: douta=16'h49a6;
16113: douta=16'h49c6;
16114: douta=16'h3966;
16115: douta=16'h4186;
16116: douta=16'h49e7;
16117: douta=16'h49e8;
16118: douta=16'h49c7;
16119: douta=16'h49e8;
16120: douta=16'h49e7;
16121: douta=16'h39a6;
16122: douta=16'h41a7;
16123: douta=16'h49e7;
16124: douta=16'h49e8;
16125: douta=16'h49c7;
16126: douta=16'h4a08;
16127: douta=16'h49e7;
16128: douta=16'h41a5;
16129: douta=16'h632e;
16130: douta=16'h3103;
16131: douta=16'h3125;
16132: douta=16'h3146;
16133: douta=16'h2967;
16134: douta=16'h430f;
16135: douta=16'h21a9;
16136: douta=16'h1946;
16137: douta=16'h1926;
16138: douta=16'h836d;
16139: douta=16'hac71;
16140: douta=16'h9c30;
16141: douta=16'ha46f;
16142: douta=16'hbcf1;
16143: douta=16'ha46f;
16144: douta=16'had34;
16145: douta=16'h8c73;
16146: douta=16'h632e;
16147: douta=16'ha514;
16148: douta=16'hb535;
16149: douta=16'h9492;
16150: douta=16'ha535;
16151: douta=16'hef1a;
16152: douta=16'he6fb;
16153: douta=16'hee74;
16154: douta=16'hde13;
16155: douta=16'hc552;
16156: douta=16'h9410;
16157: douta=16'h7b90;
16158: douta=16'h7b90;
16159: douta=16'h39e9;
16160: douta=16'h936a;
16161: douta=16'hac8d;
16162: douta=16'hd591;
16163: douta=16'hddd2;
16164: douta=16'he634;
16165: douta=16'he654;
16166: douta=16'hee96;
16167: douta=16'he634;
16168: douta=16'hddd2;
16169: douta=16'hddf3;
16170: douta=16'hde13;
16171: douta=16'hc531;
16172: douta=16'hbcf0;
16173: douta=16'hb4d1;
16174: douta=16'h9c91;
16175: douta=16'h9c93;
16176: douta=16'h8433;
16177: douta=16'h7c12;
16178: douta=16'h73b0;
16179: douta=16'h630d;
16180: douta=16'h6b71;
16181: douta=16'h3145;
16182: douta=16'h40e2;
16183: douta=16'hc4ae;
16184: douta=16'hee53;
16185: douta=16'heeb6;
16186: douta=16'heeb6;
16187: douta=16'hee95;
16188: douta=16'hee96;
16189: douta=16'he655;
16190: douta=16'hee75;
16191: douta=16'hddf3;
16192: douta=16'hd5b3;
16193: douta=16'hcd73;
16194: douta=16'hbd32;
16195: douta=16'ha4b2;
16196: douta=16'h8c52;
16197: douta=16'h8c32;
16198: douta=16'h8c53;
16199: douta=16'h8411;
16200: douta=16'h7b6f;
16201: douta=16'h7b6e;
16202: douta=16'h736d;
16203: douta=16'h732c;
16204: douta=16'h732d;
16205: douta=16'h72eb;
16206: douta=16'h6227;
16207: douta=16'h9b6a;
16208: douta=16'hb42a;
16209: douta=16'hddd0;
16210: douta=16'hd570;
16211: douta=16'hddb1;
16212: douta=16'hddd1;
16213: douta=16'hddf3;
16214: douta=16'hd5b2;
16215: douta=16'hc532;
16216: douta=16'hacd2;
16217: douta=16'ha4b2;
16218: douta=16'h9473;
16219: douta=16'h94b5;
16220: douta=16'h8454;
16221: douta=16'h7c34;
16222: douta=16'h6bf2;
16223: douta=16'h6bf3;
16224: douta=16'h6bf3;
16225: douta=16'h63d3;
16226: douta=16'h5b93;
16227: douta=16'h4b31;
16228: douta=16'h3a6e;
16229: douta=16'h2a0c;
16230: douta=16'h29eb;
16231: douta=16'h218a;
16232: douta=16'h29aa;
16233: douta=16'h1927;
16234: douta=16'h29a9;
16235: douta=16'h320c;
16236: douta=16'h322c;
16237: douta=16'h10c4;
16238: douta=16'h10e5;
16239: douta=16'h10e5;
16240: douta=16'h18e5;
16241: douta=16'h10c5;
16242: douta=16'h10e5;
16243: douta=16'h1967;
16244: douta=16'h2147;
16245: douta=16'h2147;
16246: douta=16'h1927;
16247: douta=16'h1927;
16248: douta=16'h1946;
16249: douta=16'h1926;
16250: douta=16'h10e5;
16251: douta=16'h0883;
16252: douta=16'h0042;
16253: douta=16'h0041;
16254: douta=16'h10a4;
16255: douta=16'h4acc;
16256: douta=16'h6370;
16257: douta=16'h7c14;
16258: douta=16'h2147;
16259: douta=16'h1906;
16260: douta=16'h18e5;
16261: douta=16'h73b0;
16262: douta=16'h734d;
16263: douta=16'h834b;
16264: douta=16'h5228;
16265: douta=16'h29eb;
16266: douta=16'h422c;
16267: douta=16'h634e;
16268: douta=16'h422b;
16269: douta=16'h52ed;
16270: douta=16'h08a6;
16271: douta=16'h1968;
16272: douta=16'h52ee;
16273: douta=16'h6b8f;
16274: douta=16'h426c;
16275: douta=16'h320c;
16276: douta=16'h5b2f;
16277: douta=16'h4aae;
16278: douta=16'h530f;
16279: douta=16'h42af;
16280: douta=16'h320b;
16281: douta=16'h320b;
16282: douta=16'h6b90;
16283: douta=16'h63b1;
16284: douta=16'h21aa;
16285: douta=16'h530f;
16286: douta=16'h42ef;
16287: douta=16'h5b92;
16288: douta=16'h3aaf;
16289: douta=16'h5352;
16290: douta=16'h29ea;
16291: douta=16'h21aa;
16292: douta=16'h31ea;
16293: douta=16'h840f;
16294: douta=16'h5229;
16295: douta=16'h49c7;
16296: douta=16'h49c6;
16297: douta=16'h4396;
16298: douta=16'h3166;
16299: douta=16'h38e1;
16300: douta=16'h49c6;
16301: douta=16'h51e7;
16302: douta=16'h49c6;
16303: douta=16'h51e7;
16304: douta=16'h51e7;
16305: douta=16'h49c7;
16306: douta=16'h41c7;
16307: douta=16'h4186;
16308: douta=16'h49e8;
16309: douta=16'h41a7;
16310: douta=16'h49e8;
16311: douta=16'h49e7;
16312: douta=16'h49e7;
16313: douta=16'h41a7;
16314: douta=16'h41c7;
16315: douta=16'h49c7;
16316: douta=16'h41a7;
16317: douta=16'h41a7;
16318: douta=16'h41c7;
16319: douta=16'h49e7;
16320: douta=16'h4185;
16321: douta=16'h3966;
16322: douta=16'h4228;
16323: douta=16'h3145;
16324: douta=16'h3145;
16325: douta=16'h20e4;
16326: douta=16'h4b50;
16327: douta=16'h29a9;
16328: douta=16'h29a9;
16329: douta=16'h2167;
16330: douta=16'h5a6a;
16331: douta=16'hac2e;
16332: douta=16'ha40e;
16333: douta=16'ha40e;
16334: douta=16'ha3ee;
16335: douta=16'hac4e;
16336: douta=16'h940e;
16337: douta=16'h630d;
16338: douta=16'h6b6f;
16339: douta=16'h73d0;
16340: douta=16'h73f0;
16341: douta=16'h73d1;
16342: douta=16'h73d1;
16343: douta=16'h6bb1;
16344: douta=16'h6370;
16345: douta=16'h6390;
16346: douta=16'h3aab;
16347: douta=16'hbcf1;
16348: douta=16'h736e;
16349: douta=16'h62ad;
16350: douta=16'h41a8;
16351: douta=16'hc50d;
16352: douta=16'hd590;
16353: douta=16'hd5d2;
16354: douta=16'he694;
16355: douta=16'hee96;
16356: douta=16'hee75;
16357: douta=16'hee75;
16358: douta=16'he654;
16359: douta=16'he654;
16360: douta=16'hd591;
16361: douta=16'hcd91;
16362: douta=16'hc531;
16363: douta=16'hcd93;
16364: douta=16'ha4d3;
16365: douta=16'h9c93;
16366: douta=16'h8c32;
16367: douta=16'h7bd1;
16368: douta=16'h734e;
16369: douta=16'h732e;
16370: douta=16'h6b4e;
16371: douta=16'h5acc;
16372: douta=16'h82c6;
16373: douta=16'hac0b;
16374: douta=16'hc4ac;
16375: douta=16'hff18;
16376: douta=16'he674;
16377: douta=16'h7b2d;
16378: douta=16'heeb6;
16379: douta=16'he653;
16380: douta=16'he654;
16381: douta=16'hddf3;
16382: douta=16'hc552;
16383: douta=16'hc533;
16384: douta=16'ha4d3;
16385: douta=16'hacd3;
16386: douta=16'ha4b3;
16387: douta=16'h9452;
16388: douta=16'h8c32;
16389: douta=16'h8c11;
16390: douta=16'h736e;
16391: douta=16'h7b8f;
16392: douta=16'h7b8f;
16393: douta=16'h7b6e;
16394: douta=16'h7b8e;
16395: douta=16'h6268;
16396: douta=16'hbc6d;
16397: douta=16'hc50e;
16398: douta=16'hddb0;
16399: douta=16'hee96;
16400: douta=16'he695;
16401: douta=16'hee96;
16402: douta=16'he655;
16403: douta=16'hde13;
16404: douta=16'hd5f2;
16405: douta=16'hbcb1;
16406: douta=16'ha472;
16407: douta=16'h9c72;
16408: douta=16'h9431;
16409: douta=16'h7bf1;
16410: douta=16'h7bd1;
16411: douta=16'h7bf2;
16412: douta=16'h7c12;
16413: douta=16'h7c13;
16414: douta=16'h6bb2;
16415: douta=16'h73d2;
16416: douta=16'h5b50;
16417: douta=16'h6392;
16418: douta=16'h63f4;
16419: douta=16'h6435;
16420: douta=16'h4af0;
16421: douta=16'h4af0;
16422: douta=16'h5374;
16423: douta=16'h42cf;
16424: douta=16'h2189;
16425: douta=16'h5310;
16426: douta=16'h3a8e;
16427: douta=16'h324e;
16428: douta=16'h328e;
16429: douta=16'h0882;
16430: douta=16'h18e5;
16431: douta=16'h32ae;
16432: douta=16'h10e6;
16433: douta=16'h1948;
16434: douta=16'h1947;
16435: douta=16'h1927;
16436: douta=16'h1906;
16437: douta=16'h1927;
16438: douta=16'h1927;
16439: douta=16'h1947;
16440: douta=16'h1946;
16441: douta=16'h1926;
16442: douta=16'h10c5;
16443: douta=16'h10e5;
16444: douta=16'h1926;
16445: douta=16'h1926;
16446: douta=16'h1926;
16447: douta=16'h1926;
16448: douta=16'h2127;
16449: douta=16'h2147;
16450: douta=16'h18e5;
16451: douta=16'h0883;
16452: douta=16'h0863;
16453: douta=16'h0000;
16454: douta=16'h10a2;
16455: douta=16'h426d;
16456: douta=16'h10e5;
16457: douta=16'h1927;
16458: douta=16'h1906;
16459: douta=16'h52ad;
16460: douta=16'h634e;
16461: douta=16'h424b;
16462: douta=16'h73d0;
16463: douta=16'h5b2e;
16464: douta=16'h3a0a;
16465: douta=16'h4aad;
16466: douta=16'h08e5;
16467: douta=16'h426b;
16468: douta=16'h6b90;
16469: douta=16'h532e;
16470: douta=16'h5b50;
16471: douta=16'h6390;
16472: douta=16'h3a4c;
16473: douta=16'h636f;
16474: douta=16'h5b2f;
16475: douta=16'h320b;
16476: douta=16'h5b50;
16477: douta=16'h4acd;
16478: douta=16'h29e9;
16479: douta=16'h31a8;
16480: douta=16'h29aa;
16481: douta=16'h31e9;
16482: douta=16'h4a6a;
16483: douta=16'h49a7;
16484: douta=16'h5207;
16485: douta=16'h5208;
16486: douta=16'h53f5;
16487: douta=16'h21a9;
16488: douta=16'h5207;
16489: douta=16'h5a25;
16490: douta=16'h6227;
16491: douta=16'h49a5;
16492: douta=16'h6228;
16493: douta=16'h5207;
16494: douta=16'h4186;
16495: douta=16'h4187;
16496: douta=16'h41a7;
16497: douta=16'h3966;
16498: douta=16'h49c7;
16499: douta=16'h49c7;
16500: douta=16'h49c7;
16501: douta=16'h49e8;
16502: douta=16'h49c7;
16503: douta=16'h49e7;
16504: douta=16'h41c7;
16505: douta=16'h41c7;
16506: douta=16'h41c7;
16507: douta=16'h41a7;
16508: douta=16'h41c7;
16509: douta=16'h49e8;
16510: douta=16'h41c7;
16511: douta=16'h41c7;
16512: douta=16'h3924;
16513: douta=16'h30e3;
16514: douta=16'h5b2e;
16515: douta=16'h3145;
16516: douta=16'h3125;
16517: douta=16'h2904;
16518: douta=16'h4a6b;
16519: douta=16'h2168;
16520: douta=16'h29c9;
16521: douta=16'h2188;
16522: douta=16'h522a;
16523: douta=16'ha3ed;
16524: douta=16'ha42e;
16525: douta=16'ha42e;
16526: douta=16'h9bed;
16527: douta=16'hac4e;
16528: douta=16'h83ae;
16529: douta=16'h52cd;
16530: douta=16'h632e;
16531: douta=16'h73cf;
16532: douta=16'h6baf;
16533: douta=16'h636e;
16534: douta=16'h6baf;
16535: douta=16'h6bb0;
16536: douta=16'h6bd0;
16537: douta=16'h6bd0;
16538: douta=16'h636f;
16539: douta=16'h63af;
16540: douta=16'h7bef;
16541: douta=16'hbc8d;
16542: douta=16'hdd8f;
16543: douta=16'hddd2;
16544: douta=16'hde53;
16545: douta=16'he674;
16546: douta=16'heeb6;
16547: douta=16'heeb6;
16548: douta=16'he634;
16549: douta=16'he654;
16550: douta=16'he674;
16551: douta=16'he654;
16552: douta=16'hc552;
16553: douta=16'hbd11;
16554: douta=16'ha493;
16555: douta=16'ha4d2;
16556: douta=16'h9c92;
16557: douta=16'h9472;
16558: douta=16'h7bf1;
16559: douta=16'h7b70;
16560: douta=16'h736f;
16561: douta=16'h736f;
16562: douta=16'h5a6a;
16563: douta=16'h6245;
16564: douta=16'hb44a;
16565: douta=16'he5d0;
16566: douta=16'hee75;
16567: douta=16'heeb6;
16568: douta=16'hf6f7;
16569: douta=16'h93ee;
16570: douta=16'hc4ef;
16571: douta=16'he613;
16572: douta=16'hddd2;
16573: douta=16'hb4f2;
16574: douta=16'hacb2;
16575: douta=16'ha4b3;
16576: douta=16'h9c72;
16577: douta=16'h9452;
16578: douta=16'h9452;
16579: douta=16'h8c10;
16580: douta=16'h83d0;
16581: douta=16'h7b8e;
16582: douta=16'h732d;
16583: douta=16'h732d;
16584: douta=16'h6b0c;
16585: douta=16'h4165;
16586: douta=16'h51a5;
16587: douta=16'h834a;
16588: douta=16'hbc8c;
16589: douta=16'hd58f;
16590: douta=16'hde12;
16591: douta=16'he655;
16592: douta=16'he675;
16593: douta=16'he613;
16594: douta=16'hddf3;
16595: douta=16'hddd2;
16596: douta=16'hd5b3;
16597: douta=16'hbd12;
16598: douta=16'hb4d2;
16599: douta=16'h9c72;
16600: douta=16'h9c72;
16601: douta=16'h9452;
16602: douta=16'h8412;
16603: douta=16'h7bf2;
16604: douta=16'h6b4f;
16605: douta=16'h6b70;
16606: douta=16'h6b91;
16607: douta=16'h6b91;
16608: douta=16'h73d2;
16609: douta=16'h6371;
16610: douta=16'h5b10;
16611: douta=16'h5b10;
16612: douta=16'h4ace;
16613: douta=16'h5aee;
16614: douta=16'hbcef;
16615: douta=16'h5331;
16616: douta=16'h3a4d;
16617: douta=16'h3a4d;
16618: douta=16'h5351;
16619: douta=16'h3aae;
16620: douta=16'h42af;
16621: douta=16'h322d;
16622: douta=16'h29cb;
16623: douta=16'h1106;
16624: douta=16'h29ca;
16625: douta=16'h322d;
16626: douta=16'h2989;
16627: douta=16'h1926;
16628: douta=16'h1907;
16629: douta=16'h1926;
16630: douta=16'h1946;
16631: douta=16'h1927;
16632: douta=16'h1906;
16633: douta=16'h1105;
16634: douta=16'h10e5;
16635: douta=16'h10e6;
16636: douta=16'h1906;
16637: douta=16'h1105;
16638: douta=16'h10e6;
16639: douta=16'h10e5;
16640: douta=16'h10e5;
16641: douta=16'h18e5;
16642: douta=16'h1905;
16643: douta=16'h1926;
16644: douta=16'h1926;
16645: douta=16'h2168;
16646: douta=16'h2988;
16647: douta=16'h2147;
16648: douta=16'h0862;
16649: douta=16'h0000;
16650: douta=16'h0862;
16651: douta=16'h4aad;
16652: douta=16'h5373;
16653: douta=16'h4b0f;
16654: douta=16'h5b2f;
16655: douta=16'h6b90;
16656: douta=16'h8410;
16657: douta=16'h31ea;
16658: douta=16'h5b0e;
16659: douta=16'h6b70;
16660: douta=16'h634f;
16661: douta=16'h5b70;
16662: douta=16'h322b;
16663: douta=16'h3a2b;
16664: douta=16'h5b50;
16665: douta=16'h6370;
16666: douta=16'h428d;
16667: douta=16'h5330;
16668: douta=16'h322b;
16669: douta=16'h1906;
16670: douta=16'h29a8;
16671: douta=16'h4229;
16672: douta=16'ha48d;
16673: douta=16'h6268;
16674: douta=16'h5a48;
16675: douta=16'h52ac;
16676: douta=16'h4aaf;
16677: douta=16'h2a4e;
16678: douta=16'h5248;
16679: douta=16'h6a66;
16680: douta=16'h6246;
16681: douta=16'h51e6;
16682: douta=16'h51e6;
16683: douta=16'h5a28;
16684: douta=16'h41a7;
16685: douta=16'h49c8;
16686: douta=16'h49c8;
16687: douta=16'h49c8;
16688: douta=16'h49e8;
16689: douta=16'h41a7;
16690: douta=16'h49c7;
16691: douta=16'h41a7;
16692: douta=16'h41a7;
16693: douta=16'h49c7;
16694: douta=16'h49c7;
16695: douta=16'h49c8;
16696: douta=16'h49e8;
16697: douta=16'h49c7;
16698: douta=16'h49e8;
16699: douta=16'h49e8;
16700: douta=16'h49e8;
16701: douta=16'h41a6;
16702: douta=16'h41a7;
16703: douta=16'h41c7;
16704: douta=16'h3105;
16705: douta=16'h3903;
16706: douta=16'h5b4f;
16707: douta=16'h3124;
16708: douta=16'h3125;
16709: douta=16'h2924;
16710: douta=16'h4a2a;
16711: douta=16'h2189;
16712: douta=16'h29c9;
16713: douta=16'h2988;
16714: douta=16'h3188;
16715: douta=16'h936c;
16716: douta=16'hac6e;
16717: douta=16'ha3ed;
16718: douta=16'h9bee;
16719: douta=16'hb46e;
16720: douta=16'h838e;
16721: douta=16'h52ac;
16722: douta=16'h634e;
16723: douta=16'h73d0;
16724: douta=16'h6baf;
16725: douta=16'h634e;
16726: douta=16'h636e;
16727: douta=16'h73d0;
16728: douta=16'h6bd0;
16729: douta=16'h6bf0;
16730: douta=16'h6b8f;
16731: douta=16'h6bae;
16732: douta=16'h5b8e;
16733: douta=16'hee33;
16734: douta=16'heeb5;
16735: douta=16'he633;
16736: douta=16'he654;
16737: douta=16'he674;
16738: douta=16'hee96;
16739: douta=16'heeb6;
16740: douta=16'he634;
16741: douta=16'he654;
16742: douta=16'hde13;
16743: douta=16'he614;
16744: douta=16'hc532;
16745: douta=16'hb4d2;
16746: douta=16'h9c92;
16747: douta=16'h9c93;
16748: douta=16'h8c52;
16749: douta=16'h8c52;
16750: douta=16'h7bf1;
16751: douta=16'h738f;
16752: douta=16'h732e;
16753: douta=16'h5249;
16754: douta=16'h41a5;
16755: douta=16'ha3ca;
16756: douta=16'hcced;
16757: douta=16'hee74;
16758: douta=16'heeb6;
16759: douta=16'hee96;
16760: douta=16'heeb6;
16761: douta=16'hcd92;
16762: douta=16'h7b4d;
16763: douta=16'hc531;
16764: douta=16'hd592;
16765: douta=16'hb4f2;
16766: douta=16'hb4d3;
16767: douta=16'ha493;
16768: douta=16'h8c52;
16769: douta=16'h8c11;
16770: douta=16'h83f1;
16771: douta=16'h8410;
16772: douta=16'h7b8f;
16773: douta=16'h736d;
16774: douta=16'h7b6d;
16775: douta=16'h732d;
16776: douta=16'h6b2c;
16777: douta=16'h6a87;
16778: douta=16'h8b29;
16779: douta=16'hbcad;
16780: douta=16'he5f3;
16781: douta=16'he613;
16782: douta=16'he633;
16783: douta=16'he612;
16784: douta=16'he633;
16785: douta=16'he654;
16786: douta=16'hcd51;
16787: douta=16'hc510;
16788: douta=16'hc531;
16789: douta=16'hbcd2;
16790: douta=16'hac92;
16791: douta=16'h9452;
16792: douta=16'h83f1;
16793: douta=16'h8412;
16794: douta=16'h7bd1;
16795: douta=16'h6b4f;
16796: douta=16'h6b4f;
16797: douta=16'h6b91;
16798: douta=16'h6bb2;
16799: douta=16'h73b1;
16800: douta=16'h6bd2;
16801: douta=16'h6391;
16802: douta=16'h6370;
16803: douta=16'h5b0f;
16804: douta=16'h4a2d;
16805: douta=16'hd591;
16806: douta=16'ha4f4;
16807: douta=16'h6351;
16808: douta=16'h42ce;
16809: douta=16'h322c;
16810: douta=16'h5b92;
16811: douta=16'h3a8e;
16812: douta=16'h3aae;
16813: douta=16'h42af;
16814: douta=16'h42af;
16815: douta=16'h2a0c;
16816: douta=16'h0884;
16817: douta=16'h29aa;
16818: douta=16'h3a6f;
16819: douta=16'h18e6;
16820: douta=16'h1947;
16821: douta=16'h2148;
16822: douta=16'h1906;
16823: douta=16'h1106;
16824: douta=16'h1906;
16825: douta=16'h1926;
16826: douta=16'h10e5;
16827: douta=16'h1906;
16828: douta=16'h1906;
16829: douta=16'h1905;
16830: douta=16'h10e5;
16831: douta=16'h10e5;
16832: douta=16'h10c5;
16833: douta=16'h1905;
16834: douta=16'h1905;
16835: douta=16'h1906;
16836: douta=16'h1906;
16837: douta=16'h1906;
16838: douta=16'h10e6;
16839: douta=16'h2168;
16840: douta=16'h2168;
16841: douta=16'h10e4;
16842: douta=16'h0062;
16843: douta=16'h2987;
16844: douta=16'h7c97;
16845: douta=16'h6c76;
16846: douta=16'h2126;
16847: douta=16'h4acd;
16848: douta=16'h7bf1;
16849: douta=16'h4aad;
16850: douta=16'h6b6f;
16851: douta=16'h4acc;
16852: douta=16'h634f;
16853: douta=16'h3a2c;
16854: douta=16'h94b3;
16855: douta=16'h29ea;
16856: douta=16'h21aa;
16857: douta=16'h6390;
16858: douta=16'h428c;
16859: douta=16'h5b71;
16860: douta=16'h2146;
16861: douta=16'h3a4a;
16862: douta=16'h29c9;
16863: douta=16'hbd11;
16864: douta=16'h59e7;
16865: douta=16'h6a88;
16866: douta=16'h6a67;
16867: douta=16'h4b11;
16868: douta=16'h4312;
16869: douta=16'h63f6;
16870: douta=16'h82c6;
16871: douta=16'h6247;
16872: douta=16'h6246;
16873: douta=16'h51e6;
16874: douta=16'h5a48;
16875: douta=16'h51e7;
16876: douta=16'h41a7;
16877: douta=16'h41a7;
16878: douta=16'h49e8;
16879: douta=16'h49c8;
16880: douta=16'h49e8;
16881: douta=16'h49e8;
16882: douta=16'h49c7;
16883: douta=16'h41c7;
16884: douta=16'h4186;
16885: douta=16'h49e8;
16886: douta=16'h49c7;
16887: douta=16'h49c7;
16888: douta=16'h49e8;
16889: douta=16'h5249;
16890: douta=16'h49e8;
16891: douta=16'h49e7;
16892: douta=16'h41a7;
16893: douta=16'h41a6;
16894: douta=16'h41a6;
16895: douta=16'h41a7;
16896: douta=16'h41c5;
16897: douta=16'h4165;
16898: douta=16'h5b0e;
16899: douta=16'h30e2;
16900: douta=16'h3145;
16901: douta=16'h3945;
16902: douta=16'h41c7;
16903: douta=16'h2168;
16904: douta=16'h2188;
16905: douta=16'h29a9;
16906: douta=16'h2147;
16907: douta=16'h6aab;
16908: douta=16'hac2e;
16909: douta=16'h93cd;
16910: douta=16'h9bed;
16911: douta=16'hb46f;
16912: douta=16'h736d;
16913: douta=16'h4a8c;
16914: douta=16'h6bb0;
16915: douta=16'h634e;
16916: douta=16'h6b6f;
16917: douta=16'h634e;
16918: douta=16'h6bd0;
16919: douta=16'h6bd0;
16920: douta=16'h6bb0;
16921: douta=16'h6bd0;
16922: douta=16'h638e;
16923: douta=16'h6bcf;
16924: douta=16'h6bd0;
16925: douta=16'h63b0;
16926: douta=16'h5b6e;
16927: douta=16'he6b5;
16928: douta=16'he675;
16929: douta=16'he655;
16930: douta=16'he675;
16931: douta=16'hee96;
16932: douta=16'hde34;
16933: douta=16'hcd92;
16934: douta=16'hc552;
16935: douta=16'hc552;
16936: douta=16'h9451;
16937: douta=16'h9431;
16938: douta=16'h9472;
16939: douta=16'h7bf2;
16940: douta=16'h738f;
16941: douta=16'h734f;
16942: douta=16'h6b2f;
16943: douta=16'h7bb0;
16944: douta=16'h4985;
16945: douta=16'hac2a;
16946: douta=16'hc4ad;
16947: douta=16'hd5b1;
16948: douta=16'heeb6;
16949: douta=16'hf6b6;
16950: douta=16'hee95;
16951: douta=16'hee95;
16952: douta=16'he635;
16953: douta=16'hd592;
16954: douta=16'hbd33;
16955: douta=16'ha491;
16956: douta=16'h83af;
16957: douta=16'h62ed;
16958: douta=16'h7370;
16959: douta=16'h9453;
16960: douta=16'h9452;
16961: douta=16'h8411;
16962: douta=16'h83f0;
16963: douta=16'h83cf;
16964: douta=16'h83d0;
16965: douta=16'h83af;
16966: douta=16'h62cb;
16967: douta=16'h5a26;
16968: douta=16'hbc4b;
16969: douta=16'hddf2;
16970: douta=16'hf6d6;
16971: douta=16'hddf2;
16972: douta=16'he634;
16973: douta=16'hee95;
16974: douta=16'he654;
16975: douta=16'he5d3;
16976: douta=16'hd591;
16977: douta=16'hcd52;
16978: douta=16'hc4f1;
16979: douta=16'hb4d1;
16980: douta=16'hacb1;
16981: douta=16'ha493;
16982: douta=16'h9432;
16983: douta=16'h7bb0;
16984: douta=16'h7b6f;
16985: douta=16'h734e;
16986: douta=16'h734e;
16987: douta=16'h6b0e;
16988: douta=16'h732e;
16989: douta=16'h732e;
16990: douta=16'h6b0e;
16991: douta=16'h734e;
16992: douta=16'h5acd;
16993: douta=16'h732c;
16994: douta=16'hccad;
16995: douta=16'hd54f;
16996: douta=16'hddf3;
16997: douta=16'hbd12;
16998: douta=16'h9472;
16999: douta=16'h6371;
17000: douta=16'h5b11;
17001: douta=16'h428e;
17002: douta=16'h63b3;
17003: douta=16'h5b72;
17004: douta=16'h5331;
17005: douta=16'h42af;
17006: douta=16'h42af;
17007: douta=16'h4af0;
17008: douta=16'h3a8e;
17009: douta=16'h29aa;
17010: douta=16'h322d;
17011: douta=16'h21aa;
17012: douta=16'h3a6d;
17013: douta=16'h21a8;
17014: douta=16'h21c9;
17015: douta=16'h29ca;
17016: douta=16'h2168;
17017: douta=16'h10c4;
17018: douta=16'h10e5;
17019: douta=16'h1906;
17020: douta=16'h10e5;
17021: douta=16'h10e5;
17022: douta=16'h10e5;
17023: douta=16'h10e5;
17024: douta=16'h10c5;
17025: douta=16'h1905;
17026: douta=16'h1926;
17027: douta=16'h18e5;
17028: douta=16'h10e5;
17029: douta=16'h1905;
17030: douta=16'h1905;
17031: douta=16'h18e5;
17032: douta=16'h10c5;
17033: douta=16'h10e5;
17034: douta=16'h10e5;
17035: douta=16'h1906;
17036: douta=16'h29a9;
17037: douta=16'h0001;
17038: douta=16'h2147;
17039: douta=16'h2188;
17040: douta=16'h1948;
17041: douta=16'h324c;
17042: douta=16'h73d1;
17043: douta=16'h4aad;
17044: douta=16'h5b0d;
17045: douta=16'h428c;
17046: douta=16'h6b8e;
17047: douta=16'h94b4;
17048: douta=16'h4aed;
17049: douta=16'h530f;
17050: douta=16'h1906;
17051: douta=16'h8c31;
17052: douta=16'hb4ef;
17053: douta=16'h61e6;
17054: douta=16'h6247;
17055: douta=16'h6a66;
17056: douta=16'h1149;
17057: douta=16'h21cb;
17058: douta=16'h29eb;
17059: douta=16'h63d4;
17060: douta=16'h4b31;
17061: douta=16'h3ad1;
17062: douta=16'h6a67;
17063: douta=16'h6a69;
17064: douta=16'h6a88;
17065: douta=16'h5208;
17066: douta=16'h5208;
17067: douta=16'h5229;
17068: douta=16'h49e8;
17069: douta=16'h49e8;
17070: douta=16'h49e8;
17071: douta=16'h49e8;
17072: douta=16'h41a7;
17073: douta=16'h41a7;
17074: douta=16'h41a7;
17075: douta=16'h41a7;
17076: douta=16'h41c7;
17077: douta=16'h49c7;
17078: douta=16'h49e8;
17079: douta=16'h49e8;
17080: douta=16'h49e8;
17081: douta=16'h41a7;
17082: douta=16'h49e7;
17083: douta=16'h41a7;
17084: douta=16'h3986;
17085: douta=16'h49e7;
17086: douta=16'h41c7;
17087: douta=16'h41a7;
17088: douta=16'h8b88;
17089: douta=16'h4165;
17090: douta=16'h4a09;
17091: douta=16'h3124;
17092: douta=16'h3145;
17093: douta=16'h3124;
17094: douta=16'h3145;
17095: douta=16'h2168;
17096: douta=16'h29a9;
17097: douta=16'h29c9;
17098: douta=16'h39e9;
17099: douta=16'h7b4c;
17100: douta=16'h8b8d;
17101: douta=16'h8bad;
17102: douta=16'hac4e;
17103: douta=16'hac4e;
17104: douta=16'h6b2d;
17105: douta=16'h5aed;
17106: douta=16'h634e;
17107: douta=16'h6b8f;
17108: douta=16'h636e;
17109: douta=16'h6bb0;
17110: douta=16'h6bd0;
17111: douta=16'h73d0;
17112: douta=16'h6bb0;
17113: douta=16'h6baf;
17114: douta=16'h636f;
17115: douta=16'h638f;
17116: douta=16'h6bcf;
17117: douta=16'h6baf;
17118: douta=16'h6bd0;
17119: douta=16'hc511;
17120: douta=16'hf6f6;
17121: douta=16'hee96;
17122: douta=16'hee96;
17123: douta=16'hde34;
17124: douta=16'hddf3;
17125: douta=16'hc552;
17126: douta=16'hb4d1;
17127: douta=16'hac91;
17128: douta=16'h9451;
17129: douta=16'h9431;
17130: douta=16'h7bf1;
17131: douta=16'h736f;
17132: douta=16'h6b4f;
17133: douta=16'h734f;
17134: douta=16'h62cd;
17135: douta=16'h51e5;
17136: douta=16'ha42b;
17137: douta=16'hc50f;
17138: douta=16'hd591;
17139: douta=16'he695;
17140: douta=16'hf6b6;
17141: douta=16'hee95;
17142: douta=16'hee75;
17143: douta=16'he613;
17144: douta=16'hd5d3;
17145: douta=16'hcd73;
17146: douta=16'hb4b2;
17147: douta=16'h9c93;
17148: douta=16'h9494;
17149: douta=16'h9474;
17150: douta=16'h8c54;
17151: douta=16'h7390;
17152: douta=16'h73d1;
17153: douta=16'h7bf2;
17154: douta=16'h7391;
17155: douta=16'h7390;
17156: douta=16'h5aef;
17157: douta=16'h520a;
17158: douta=16'h936a;
17159: douta=16'hcd0e;
17160: douta=16'he633;
17161: douta=16'he612;
17162: douta=16'hd570;
17163: douta=16'hee75;
17164: douta=16'he634;
17165: douta=16'hddf3;
17166: douta=16'he634;
17167: douta=16'hd591;
17168: douta=16'hcd50;
17169: douta=16'hacb1;
17170: douta=16'h9431;
17171: douta=16'h9411;
17172: douta=16'h9411;
17173: douta=16'h83b0;
17174: douta=16'h838f;
17175: douta=16'h732c;
17176: douta=16'h732d;
17177: douta=16'h730d;
17178: douta=16'h7b6e;
17179: douta=16'h734e;
17180: douta=16'h62cd;
17181: douta=16'h5acc;
17182: douta=16'h836d;
17183: douta=16'h734d;
17184: douta=16'ha3ec;
17185: douta=16'hf6b7;
17186: douta=16'heeb7;
17187: douta=16'he675;
17188: douta=16'hcd93;
17189: douta=16'ha4b2;
17190: douta=16'ha4b3;
17191: douta=16'h6b91;
17192: douta=16'h5b50;
17193: douta=16'h5310;
17194: douta=16'h6392;
17195: douta=16'h5b72;
17196: douta=16'h5331;
17197: douta=16'h42af;
17198: douta=16'h4acf;
17199: douta=16'h4acf;
17200: douta=16'h320c;
17201: douta=16'h42af;
17202: douta=16'h42cf;
17203: douta=16'h3a2d;
17204: douta=16'h21aa;
17205: douta=16'h3a6d;
17206: douta=16'h2189;
17207: douta=16'h10a5;
17208: douta=16'h10e5;
17209: douta=16'h2189;
17210: douta=16'h29ca;
17211: douta=16'h21a9;
17212: douta=16'h08c4;
17213: douta=16'h10e5;
17214: douta=16'h1905;
17215: douta=16'h10c5;
17216: douta=16'h18e5;
17217: douta=16'h10e5;
17218: douta=16'h18e5;
17219: douta=16'h1905;
17220: douta=16'h10e5;
17221: douta=16'h1906;
17222: douta=16'h1906;
17223: douta=16'h1905;
17224: douta=16'h10c5;
17225: douta=16'h1905;
17226: douta=16'h1905;
17227: douta=16'h1905;
17228: douta=16'h18e5;
17229: douta=16'h18e5;
17230: douta=16'h1927;
17231: douta=16'h0884;
17232: douta=16'h08a3;
17233: douta=16'h7477;
17234: douta=16'h3a8d;
17235: douta=16'h530f;
17236: douta=16'h6b90;
17237: douta=16'h5b0e;
17238: douta=16'h94d3;
17239: douta=16'h2166;
17240: douta=16'h4a4a;
17241: douta=16'h322a;
17242: douta=16'hc530;
17243: douta=16'h7aa8;
17244: douta=16'h7aa6;
17245: douta=16'h5229;
17246: douta=16'h29a9;
17247: douta=16'h2a4c;
17248: douta=16'h3a4c;
17249: douta=16'h5b51;
17250: douta=16'h3aae;
17251: douta=16'h3a6e;
17252: douta=16'h322d;
17253: douta=16'h222e;
17254: douta=16'h72a9;
17255: douta=16'h6a68;
17256: douta=16'h6249;
17257: douta=16'h5228;
17258: douta=16'h5a49;
17259: douta=16'h5208;
17260: douta=16'h5229;
17261: douta=16'h5249;
17262: douta=16'h49e8;
17263: douta=16'h49e8;
17264: douta=16'h49c7;
17265: douta=16'h41a7;
17266: douta=16'h41a7;
17267: douta=16'h41a7;
17268: douta=16'h41a7;
17269: douta=16'h39a6;
17270: douta=16'h49e8;
17271: douta=16'h49e8;
17272: douta=16'h41a7;
17273: douta=16'h49e7;
17274: douta=16'h41c7;
17275: douta=16'h41a7;
17276: douta=16'h41a7;
17277: douta=16'h41a7;
17278: douta=16'h49e7;
17279: douta=16'h41a7;
17280: douta=16'hac69;
17281: douta=16'h4165;
17282: douta=16'h4186;
17283: douta=16'h39a6;
17284: douta=16'h3125;
17285: douta=16'h3145;
17286: douta=16'h2925;
17287: douta=16'h2188;
17288: douta=16'h2969;
17289: douta=16'h2168;
17290: douta=16'h526b;
17291: douta=16'h7b2c;
17292: douta=16'h732c;
17293: douta=16'h834c;
17294: douta=16'ha40d;
17295: douta=16'h9bed;
17296: douta=16'h52cc;
17297: douta=16'h52cd;
17298: douta=16'h636f;
17299: douta=16'h636e;
17300: douta=16'h634e;
17301: douta=16'h73d0;
17302: douta=16'h7411;
17303: douta=16'h73f1;
17304: douta=16'h7c11;
17305: douta=16'h63af;
17306: douta=16'h5b4e;
17307: douta=16'h5b4e;
17308: douta=16'h6baf;
17309: douta=16'h6bcf;
17310: douta=16'h6bd0;
17311: douta=16'h5b4e;
17312: douta=16'hfeb5;
17313: douta=16'hee96;
17314: douta=16'he675;
17315: douta=16'he655;
17316: douta=16'hd5b2;
17317: douta=16'hc531;
17318: douta=16'ha490;
17319: douta=16'ha471;
17320: douta=16'h9c72;
17321: douta=16'h9432;
17322: douta=16'h73b0;
17323: douta=16'h738f;
17324: douta=16'h6b4f;
17325: douta=16'h734e;
17326: douta=16'h4187;
17327: douta=16'ha3ea;
17328: douta=16'hbcad;
17329: douta=16'hddf3;
17330: douta=16'he654;
17331: douta=16'hf6d7;
17332: douta=16'heeb7;
17333: douta=16'hee95;
17334: douta=16'hee75;
17335: douta=16'hd5d2;
17336: douta=16'hd591;
17337: douta=16'hbcf2;
17338: douta=16'hacd3;
17339: douta=16'h9494;
17340: douta=16'h8c54;
17341: douta=16'h8c54;
17342: douta=16'h8c53;
17343: douta=16'h8c73;
17344: douta=16'h6b90;
17345: douta=16'h6370;
17346: douta=16'h6330;
17347: douta=16'h6b2e;
17348: douta=16'h49e7;
17349: douta=16'h59e6;
17350: douta=16'hb42b;
17351: douta=16'hbcee;
17352: douta=16'hff17;
17353: douta=16'heeb6;
17354: douta=16'he654;
17355: douta=16'hac0c;
17356: douta=16'he673;
17357: douta=16'hcd30;
17358: douta=16'hddd1;
17359: douta=16'hac70;
17360: douta=16'hb4d1;
17361: douta=16'ha472;
17362: douta=16'h9c31;
17363: douta=16'h8c10;
17364: douta=16'h8bf1;
17365: douta=16'h8c11;
17366: douta=16'h7b8f;
17367: douta=16'h7b6e;
17368: douta=16'h730c;
17369: douta=16'h6aeb;
17370: douta=16'h734d;
17371: douta=16'h732d;
17372: douta=16'h41ea;
17373: douta=16'h298a;
17374: douta=16'hc50f;
17375: douta=16'hcd71;
17376: douta=16'hb48e;
17377: douta=16'he696;
17378: douta=16'hde35;
17379: douta=16'hd5f4;
17380: douta=16'hacb3;
17381: douta=16'h9c94;
17382: douta=16'h9493;
17383: douta=16'h6371;
17384: douta=16'h530f;
17385: douta=16'h5330;
17386: douta=16'h6392;
17387: douta=16'h5351;
17388: douta=16'h5330;
17389: douta=16'h42ae;
17390: douta=16'h428e;
17391: douta=16'h42af;
17392: douta=16'h42ae;
17393: douta=16'h4ad0;
17394: douta=16'h4b10;
17395: douta=16'h734d;
17396: douta=16'h218a;
17397: douta=16'h4b10;
17398: douta=16'h324d;
17399: douta=16'h2988;
17400: douta=16'h2147;
17401: douta=16'h1084;
17402: douta=16'h10e5;
17403: douta=16'h2147;
17404: douta=16'h2167;
17405: douta=16'h1926;
17406: douta=16'h10e5;
17407: douta=16'h10e5;
17408: douta=16'h18e5;
17409: douta=16'h18e5;
17410: douta=16'h1905;
17411: douta=16'h10c4;
17412: douta=16'h10e5;
17413: douta=16'h1905;
17414: douta=16'h18e5;
17415: douta=16'h10e5;
17416: douta=16'h10e5;
17417: douta=16'h1926;
17418: douta=16'h1905;
17419: douta=16'h1905;
17420: douta=16'h1905;
17421: douta=16'h1905;
17422: douta=16'h1926;
17423: douta=16'h2147;
17424: douta=16'h0021;
17425: douta=16'h530f;
17426: douta=16'h6c14;
17427: douta=16'h6391;
17428: douta=16'h7411;
17429: douta=16'h636f;
17430: douta=16'h6b8e;
17431: douta=16'h4aab;
17432: douta=16'ha4d2;
17433: douta=16'hc5b3;
17434: douta=16'h7ac7;
17435: douta=16'h7aa7;
17436: douta=16'h6227;
17437: douta=16'h2a0c;
17438: douta=16'h2a2c;
17439: douta=16'h3aae;
17440: douta=16'h4aee;
17441: douta=16'h4acf;
17442: douta=16'h42ad;
17443: douta=16'h3a4c;
17444: douta=16'h31eb;
17445: douta=16'h4b52;
17446: douta=16'h6a88;
17447: douta=16'h6a69;
17448: douta=16'h5228;
17449: douta=16'h5228;
17450: douta=16'h5228;
17451: douta=16'h49e7;
17452: douta=16'h5249;
17453: douta=16'h5249;
17454: douta=16'h5209;
17455: douta=16'h49c7;
17456: douta=16'h41c7;
17457: douta=16'h4186;
17458: douta=16'h41c7;
17459: douta=16'h41c7;
17460: douta=16'h41c7;
17461: douta=16'h3987;
17462: douta=16'h49c7;
17463: douta=16'h49c8;
17464: douta=16'h49e7;
17465: douta=16'h49c7;
17466: douta=16'h49e7;
17467: douta=16'h3986;
17468: douta=16'h41a7;
17469: douta=16'h49e7;
17470: douta=16'h49e7;
17471: douta=16'h49e7;
17472: douta=16'hf5cb;
17473: douta=16'h4185;
17474: douta=16'h38e3;
17475: douta=16'h52ed;
17476: douta=16'h3124;
17477: douta=16'h3124;
17478: douta=16'h2904;
17479: douta=16'h2168;
17480: douta=16'h2188;
17481: douta=16'h2188;
17482: douta=16'h5aac;
17483: douta=16'h5a8b;
17484: douta=16'h62cc;
17485: douta=16'h72ec;
17486: douta=16'h6aec;
17487: douta=16'h730d;
17488: douta=16'h4a8b;
17489: douta=16'h4aad;
17490: douta=16'h52ee;
17491: douta=16'h636f;
17492: douta=16'h6b8f;
17493: douta=16'h6bb0;
17494: douta=16'h6bb0;
17495: douta=16'h6bd0;
17496: douta=16'h7411;
17497: douta=16'h73f1;
17498: douta=16'h6bcf;
17499: douta=16'h638f;
17500: douta=16'h6baf;
17501: douta=16'h638f;
17502: douta=16'h6bcf;
17503: douta=16'h6bf0;
17504: douta=16'h6bd0;
17505: douta=16'h5b0d;
17506: douta=16'he634;
17507: douta=16'hd5d3;
17508: douta=16'hd5b2;
17509: douta=16'ha450;
17510: douta=16'ha4b1;
17511: douta=16'hb4d2;
17512: douta=16'h6b2f;
17513: douta=16'h6b2e;
17514: douta=16'h7370;
17515: douta=16'h734f;
17516: douta=16'h420a;
17517: douta=16'h4187;
17518: douta=16'hcd2e;
17519: douta=16'hd5b0;
17520: douta=16'heeb6;
17521: douta=16'heed7;
17522: douta=16'heeb6;
17523: douta=16'heeb6;
17524: douta=16'hee96;
17525: douta=16'he634;
17526: douta=16'hd5f3;
17527: douta=16'hbcf2;
17528: douta=16'hacb3;
17529: douta=16'h9cb4;
17530: douta=16'h8455;
17531: douta=16'h8455;
17532: douta=16'h8454;
17533: douta=16'h7bd1;
17534: douta=16'h7bd1;
17535: douta=16'h7b90;
17536: douta=16'h62ed;
17537: douta=16'h632e;
17538: douta=16'h528b;
17539: douta=16'h72a8;
17540: douta=16'hc4ac;
17541: douta=16'hcd0e;
17542: douta=16'heed7;
17543: douta=16'hee95;
17544: douta=16'hd591;
17545: douta=16'he654;
17546: douta=16'hee95;
17547: douta=16'hee94;
17548: douta=16'h93cd;
17549: douta=16'hac70;
17550: douta=16'hac90;
17551: douta=16'h8c10;
17552: douta=16'h8bf0;
17553: douta=16'h838e;
17554: douta=16'h838e;
17555: douta=16'h7b4d;
17556: douta=16'h730c;
17557: douta=16'h730c;
17558: douta=16'h732c;
17559: douta=16'h838e;
17560: douta=16'h7b4d;
17561: douta=16'h6acb;
17562: douta=16'h628b;
17563: douta=16'hee75;
17564: douta=16'hd5d4;
17565: douta=16'hde15;
17566: douta=16'heeb8;
17567: douta=16'hee97;
17568: douta=16'hd5f5;
17569: douta=16'hbd54;
17570: douta=16'had14;
17571: douta=16'had15;
17572: douta=16'ha4b4;
17573: douta=16'h9c94;
17574: douta=16'h9494;
17575: douta=16'h7bf2;
17576: douta=16'h73b1;
17577: douta=16'h6350;
17578: douta=16'h5b30;
17579: douta=16'h530f;
17580: douta=16'h4acf;
17581: douta=16'h532f;
17582: douta=16'h5330;
17583: douta=16'h5b50;
17584: douta=16'h4af0;
17585: douta=16'h630e;
17586: douta=16'hc4f0;
17587: douta=16'h5bb2;
17588: douta=16'h3a6e;
17589: douta=16'h63b2;
17590: douta=16'h42af;
17591: douta=16'h4af0;
17592: douta=16'h328e;
17593: douta=16'h322c;
17594: douta=16'h2189;
17595: douta=16'h21aa;
17596: douta=16'h1927;
17597: douta=16'h1927;
17598: douta=16'h1947;
17599: douta=16'h3aaf;
17600: douta=16'h2a2c;
17601: douta=16'h2148;
17602: douta=16'h2167;
17603: douta=16'h29a9;
17604: douta=16'h29a9;
17605: douta=16'h18e5;
17606: douta=16'h10e4;
17607: douta=16'h10c4;
17608: douta=16'h1947;
17609: douta=16'h1926;
17610: douta=16'h10c5;
17611: douta=16'h18e5;
17612: douta=16'h18e5;
17613: douta=16'h10e5;
17614: douta=16'h10c4;
17615: douta=16'h10a4;
17616: douta=16'h1905;
17617: douta=16'h10e5;
17618: douta=16'h0042;
17619: douta=16'h0000;
17620: douta=16'h2146;
17621: douta=16'h10c6;
17622: douta=16'hcd92;
17623: douta=16'h8267;
17624: douta=16'h9327;
17625: douta=16'h82e9;
17626: douta=16'h324d;
17627: douta=16'h6391;
17628: douta=16'h29cb;
17629: douta=16'h4aad;
17630: douta=16'h29eb;
17631: douta=16'h5b50;
17632: douta=16'h4b0f;
17633: douta=16'h5330;
17634: douta=16'h5b71;
17635: douta=16'h328f;
17636: douta=16'h4b10;
17637: douta=16'h6bf4;
17638: douta=16'h6acc;
17639: douta=16'h6268;
17640: douta=16'h6289;
17641: douta=16'h5229;
17642: douta=16'h5228;
17643: douta=16'h5249;
17644: douta=16'h49e8;
17645: douta=16'h41a7;
17646: douta=16'h41a7;
17647: douta=16'h41a7;
17648: douta=16'h41a7;
17649: douta=16'h41c7;
17650: douta=16'h41c7;
17651: douta=16'h41c7;
17652: douta=16'h41a7;
17653: douta=16'h41a6;
17654: douta=16'h41a7;
17655: douta=16'h41c7;
17656: douta=16'h39a6;
17657: douta=16'h41a6;
17658: douta=16'h41c7;
17659: douta=16'h41c7;
17660: douta=16'h41a7;
17661: douta=16'h49c7;
17662: douta=16'h49c8;
17663: douta=16'h41a7;
17664: douta=16'hed8b;
17665: douta=16'h3124;
17666: douta=16'h3944;
17667: douta=16'h634f;
17668: douta=16'h3144;
17669: douta=16'h3124;
17670: douta=16'h3124;
17671: douta=16'h29ca;
17672: douta=16'h29a8;
17673: douta=16'h29a9;
17674: douta=16'h52ac;
17675: douta=16'h4a4a;
17676: douta=16'h5a8b;
17677: douta=16'h526a;
17678: douta=16'h5aac;
17679: douta=16'h5acd;
17680: douta=16'h426b;
17681: douta=16'h52cd;
17682: douta=16'h530e;
17683: douta=16'h634e;
17684: douta=16'h636f;
17685: douta=16'h6bd0;
17686: douta=16'h73f1;
17687: douta=16'h6bd0;
17688: douta=16'h73f0;
17689: douta=16'h73f1;
17690: douta=16'h6bcf;
17691: douta=16'h6bd0;
17692: douta=16'h6baf;
17693: douta=16'h638f;
17694: douta=16'h6baf;
17695: douta=16'h6bcf;
17696: douta=16'h6bd0;
17697: douta=16'h634e;
17698: douta=16'h736e;
17699: douta=16'hc531;
17700: douta=16'hcd52;
17701: douta=16'hac90;
17702: douta=16'h8bcf;
17703: douta=16'h8bf0;
17704: douta=16'h7bd0;
17705: douta=16'h7b6f;
17706: douta=16'h734e;
17707: douta=16'h3a2b;
17708: douta=16'h9b6a;
17709: douta=16'hbc4b;
17710: douta=16'hd5d2;
17711: douta=16'hee96;
17712: douta=16'heeb6;
17713: douta=16'heeb7;
17714: douta=16'heeb7;
17715: douta=16'he676;
17716: douta=16'he634;
17717: douta=16'hd5b3;
17718: douta=16'hbd32;
17719: douta=16'h9c93;
17720: douta=16'h9474;
17721: douta=16'h8c53;
17722: douta=16'h8454;
17723: douta=16'h7bd1;
17724: douta=16'h7390;
17725: douta=16'h6b4e;
17726: douta=16'h6b2e;
17727: douta=16'h6b0e;
17728: douta=16'h62cd;
17729: douta=16'h49a7;
17730: douta=16'h7287;
17731: douta=16'h8b28;
17732: douta=16'hee75;
17733: douta=16'hee75;
17734: douta=16'hbcac;
17735: douta=16'hf6d7;
17736: douta=16'ha470;
17737: douta=16'hee54;
17738: douta=16'he674;
17739: douta=16'hcd71;
17740: douta=16'ha490;
17741: douta=16'ha471;
17742: douta=16'h9431;
17743: douta=16'h83cf;
17744: douta=16'h7baf;
17745: douta=16'h734e;
17746: douta=16'h730d;
17747: douta=16'h7b6e;
17748: douta=16'h838e;
17749: douta=16'h62aa;
17750: douta=16'h5249;
17751: douta=16'h41e8;
17752: douta=16'h832b;
17753: douta=16'hbc8f;
17754: douta=16'hc531;
17755: douta=16'hac6d;
17756: douta=16'hd5d4;
17757: douta=16'hc573;
17758: douta=16'hd5d4;
17759: douta=16'hcdd5;
17760: douta=16'hcdb5;
17761: douta=16'hbd55;
17762: douta=16'hb535;
17763: douta=16'had15;
17764: douta=16'h9cd5;
17765: douta=16'h9494;
17766: douta=16'h8c93;
17767: douta=16'h8433;
17768: douta=16'h73d1;
17769: douta=16'h73b1;
17770: douta=16'h6350;
17771: douta=16'h5b30;
17772: douta=16'h5b0f;
17773: douta=16'h52ee;
17774: douta=16'h4ace;
17775: douta=16'h4ace;
17776: douta=16'hcd11;
17777: douta=16'hddd3;
17778: douta=16'hee35;
17779: douta=16'h6bf3;
17780: douta=16'h5350;
17781: douta=16'h6bd3;
17782: douta=16'h5310;
17783: douta=16'h4af0;
17784: douta=16'h3a8e;
17785: douta=16'h322c;
17786: douta=16'h29ca;
17787: douta=16'h29ca;
17788: douta=16'h1947;
17789: douta=16'h1927;
17790: douta=16'h29ca;
17791: douta=16'h29cb;
17792: douta=16'h42d0;
17793: douta=16'h29cb;
17794: douta=16'h10e5;
17795: douta=16'h2147;
17796: douta=16'h1927;
17797: douta=16'h2168;
17798: douta=16'h2169;
17799: douta=16'h29aa;
17800: douta=16'h29eb;
17801: douta=16'h29aa;
17802: douta=16'h1906;
17803: douta=16'h10c3;
17804: douta=16'h10e5;
17805: douta=16'h10e5;
17806: douta=16'h10e5;
17807: douta=16'h10e5;
17808: douta=16'h1905;
17809: douta=16'h0884;
17810: douta=16'h10c4;
17811: douta=16'h1905;
17812: douta=16'h08a3;
17813: douta=16'h10e5;
17814: douta=16'h08c6;
17815: douta=16'h7b2b;
17816: douta=16'h3a4d;
17817: douta=16'h320c;
17818: douta=16'h7413;
17819: douta=16'h428e;
17820: douta=16'h320c;
17821: douta=16'h4aad;
17822: douta=16'h7c13;
17823: douta=16'h5b71;
17824: douta=16'h5b71;
17825: douta=16'h5330;
17826: douta=16'h42af;
17827: douta=16'h4b0f;
17828: douta=16'h73f4;
17829: douta=16'h3a8e;
17830: douta=16'h4b31;
17831: douta=16'had34;
17832: douta=16'h6248;
17833: douta=16'h5229;
17834: douta=16'h5249;
17835: douta=16'h5208;
17836: douta=16'h49c8;
17837: douta=16'h49c7;
17838: douta=16'h41a7;
17839: douta=16'h41a7;
17840: douta=16'h49c7;
17841: douta=16'h49e8;
17842: douta=16'h3986;
17843: douta=16'h39a6;
17844: douta=16'h49c7;
17845: douta=16'h41a7;
17846: douta=16'h4186;
17847: douta=16'h4186;
17848: douta=16'h41a6;
17849: douta=16'h3986;
17850: douta=16'h39a6;
17851: douta=16'h41a7;
17852: douta=16'h41a7;
17853: douta=16'h49e7;
17854: douta=16'h4187;
17855: douta=16'h49e8;
17856: douta=16'he52a;
17857: douta=16'h28e3;
17858: douta=16'h3965;
17859: douta=16'h632f;
17860: douta=16'h3145;
17861: douta=16'h3124;
17862: douta=16'h3124;
17863: douta=16'h3a6c;
17864: douta=16'h2168;
17865: douta=16'h2168;
17866: douta=16'h528b;
17867: douta=16'h422a;
17868: douta=16'h4a0a;
17869: douta=16'h4209;
17870: douta=16'h528b;
17871: douta=16'h52cc;
17872: douta=16'h426b;
17873: douta=16'h52ce;
17874: douta=16'h5b0e;
17875: douta=16'h634f;
17876: douta=16'h6390;
17877: douta=16'h6b90;
17878: douta=16'h6bd0;
17879: douta=16'h73f1;
17880: douta=16'h73f1;
17881: douta=16'h7411;
17882: douta=16'h6bd0;
17883: douta=16'h6baf;
17884: douta=16'h6bcf;
17885: douta=16'h638f;
17886: douta=16'h63af;
17887: douta=16'h6bcf;
17888: douta=16'h636e;
17889: douta=16'h5b0d;
17890: douta=16'h3a6b;
17891: douta=16'h426b;
17892: douta=16'hddb2;
17893: douta=16'hac90;
17894: douta=16'h93ef;
17895: douta=16'h7b6e;
17896: douta=16'h734e;
17897: douta=16'h6b0d;
17898: douta=16'h5aab;
17899: douta=16'h3987;
17900: douta=16'hcd0e;
17901: douta=16'hc50c;
17902: douta=16'hde13;
17903: douta=16'heeb6;
17904: douta=16'heed7;
17905: douta=16'heeb7;
17906: douta=16'hee96;
17907: douta=16'he655;
17908: douta=16'hd5d3;
17909: douta=16'hc552;
17910: douta=16'hb513;
17911: douta=16'h8c74;
17912: douta=16'h8454;
17913: douta=16'h8413;
17914: douta=16'h8412;
17915: douta=16'h73b0;
17916: douta=16'h6b6f;
17917: douta=16'h6b4e;
17918: douta=16'h6b0d;
17919: douta=16'h62cd;
17920: douta=16'h49a6;
17921: douta=16'h59c6;
17922: douta=16'h9348;
17923: douta=16'hd570;
17924: douta=16'hee75;
17925: douta=16'hee96;
17926: douta=16'he633;
17927: douta=16'hee75;
17928: douta=16'hee73;
17929: douta=16'h8b6b;
17930: douta=16'hac6e;
17931: douta=16'hc511;
17932: douta=16'ha491;
17933: douta=16'h9431;
17934: douta=16'h9411;
17935: douta=16'h7b90;
17936: douta=16'h734e;
17937: douta=16'h732d;
17938: douta=16'h6acc;
17939: douta=16'h6aec;
17940: douta=16'h732c;
17941: douta=16'h7b4d;
17942: douta=16'h62cc;
17943: douta=16'h62aa;
17944: douta=16'hd52e;
17945: douta=16'hddd1;
17946: douta=16'hf6b6;
17947: douta=16'hd5f4;
17948: douta=16'hddf4;
17949: douta=16'he655;
17950: douta=16'hcd93;
17951: douta=16'hc594;
17952: douta=16'hacd3;
17953: douta=16'hb535;
17954: douta=16'had15;
17955: douta=16'ha4f5;
17956: douta=16'h9cd4;
17957: douta=16'h94b4;
17958: douta=16'h8c73;
17959: douta=16'h7bf1;
17960: douta=16'h7bf2;
17961: douta=16'h7390;
17962: douta=16'h634f;
17963: douta=16'h5b0e;
17964: douta=16'h5aee;
17965: douta=16'h4aae;
17966: douta=16'h4a8d;
17967: douta=16'h93ee;
17968: douta=16'he655;
17969: douta=16'hcdb5;
17970: douta=16'ha4b3;
17971: douta=16'h6371;
17972: douta=16'h4acf;
17973: douta=16'h5b50;
17974: douta=16'h4ad0;
17975: douta=16'h4aef;
17976: douta=16'h428e;
17977: douta=16'h3a4d;
17978: douta=16'h29aa;
17979: douta=16'h29aa;
17980: douta=16'h2168;
17981: douta=16'h29a9;
17982: douta=16'h1127;
17983: douta=16'h21aa;
17984: douta=16'h5311;
17985: douta=16'h21aa;
17986: douta=16'h1967;
17987: douta=16'h29cb;
17988: douta=16'h3a4e;
17989: douta=16'h1989;
17990: douta=16'h21a9;
17991: douta=16'h2189;
17992: douta=16'h2a0b;
17993: douta=16'h218a;
17994: douta=16'h29cb;
17995: douta=16'h29a9;
17996: douta=16'h1906;
17997: douta=16'h10e4;
17998: douta=16'h10e5;
17999: douta=16'h10e5;
18000: douta=16'h1905;
18001: douta=16'h1084;
18002: douta=16'h08a4;
18003: douta=16'h10e5;
18004: douta=16'h1105;
18005: douta=16'h10c4;
18006: douta=16'h1906;
18007: douta=16'h428e;
18008: douta=16'h29eb;
18009: douta=16'h428d;
18010: douta=16'h5b30;
18011: douta=16'h52ef;
18012: douta=16'h5b50;
18013: douta=16'h6bd2;
18014: douta=16'h6b71;
18015: douta=16'h5b30;
18016: douta=16'h6371;
18017: douta=16'h4b10;
18018: douta=16'h5b93;
18019: douta=16'h5b92;
18020: douta=16'h5351;
18021: douta=16'h5351;
18022: douta=16'h6c14;
18023: douta=16'hc67b;
18024: douta=16'hb5b7;
18025: douta=16'h5a28;
18026: douta=16'h49e8;
18027: douta=16'h5228;
18028: douta=16'h49c8;
18029: douta=16'h41a7;
18030: douta=16'h41a7;
18031: douta=16'h41c7;
18032: douta=16'h41a7;
18033: douta=16'h41c7;
18034: douta=16'h41a7;
18035: douta=16'h41a7;
18036: douta=16'h41a7;
18037: douta=16'h41a7;
18038: douta=16'h41a6;
18039: douta=16'h41a7;
18040: douta=16'h3986;
18041: douta=16'h41a7;
18042: douta=16'h3986;
18043: douta=16'h39a6;
18044: douta=16'h41a7;
18045: douta=16'h49c8;
18046: douta=16'h41a7;
18047: douta=16'h41a7;
18048: douta=16'hdd2a;
18049: douta=16'h51e5;
18050: douta=16'h3945;
18051: douta=16'h41a6;
18052: douta=16'h2904;
18053: douta=16'h2924;
18054: douta=16'h3124;
18055: douta=16'h320a;
18056: douta=16'h2188;
18057: douta=16'h1967;
18058: douta=16'h424b;
18059: douta=16'h422b;
18060: douta=16'h3a0a;
18061: douta=16'h31a8;
18062: douta=16'h3a2a;
18063: douta=16'h4a8c;
18064: douta=16'h428c;
18065: douta=16'h4acd;
18066: douta=16'h4acd;
18067: douta=16'h5b4f;
18068: douta=16'h6390;
18069: douta=16'h63b0;
18070: douta=16'h6bb1;
18071: douta=16'h6bb0;
18072: douta=16'h6bb0;
18073: douta=16'h73f1;
18074: douta=16'h5b6f;
18075: douta=16'h5b6e;
18076: douta=16'h638f;
18077: douta=16'h6baf;
18078: douta=16'h6bcf;
18079: douta=16'h638f;
18080: douta=16'h6bcf;
18081: douta=16'h6bd0;
18082: douta=16'h63af;
18083: douta=16'h5b2d;
18084: douta=16'h5b4d;
18085: douta=16'h6b6e;
18086: douta=16'ha470;
18087: douta=16'h9c50;
18088: douta=16'h6b0d;
18089: douta=16'h62ec;
18090: douta=16'h398a;
18091: douta=16'he675;
18092: douta=16'hde34;
18093: douta=16'he696;
18094: douta=16'he655;
18095: douta=16'heed7;
18096: douta=16'he655;
18097: douta=16'hde34;
18098: douta=16'he634;
18099: douta=16'hcdb3;
18100: douta=16'hbd54;
18101: douta=16'hbd73;
18102: douta=16'hb533;
18103: douta=16'h8c54;
18104: douta=16'h8433;
18105: douta=16'h7c12;
18106: douta=16'h738f;
18107: douta=16'h7390;
18108: douta=16'h7390;
18109: douta=16'h632e;
18110: douta=16'h6aed;
18111: douta=16'h4146;
18112: douta=16'hccee;
18113: douta=16'hdd90;
18114: douta=16'hee95;
18115: douta=16'hd5d2;
18116: douta=16'hac4e;
18117: douta=16'hf694;
18118: douta=16'he5f3;
18119: douta=16'hb511;
18120: douta=16'hb4b1;
18121: douta=16'ha472;
18122: douta=16'ha492;
18123: douta=16'h9472;
18124: douta=16'h736f;
18125: douta=16'h7b8f;
18126: douta=16'h9411;
18127: douta=16'h7b90;
18128: douta=16'h83af;
18129: douta=16'h8bf0;
18130: douta=16'h7b4d;
18131: douta=16'h7b2d;
18132: douta=16'h6aec;
18133: douta=16'hb40c;
18134: douta=16'he632;
18135: douta=16'hd591;
18136: douta=16'hd5b3;
18137: douta=16'hde13;
18138: douta=16'hde14;
18139: douta=16'hb533;
18140: douta=16'hb4f4;
18141: douta=16'hacd4;
18142: douta=16'hbd74;
18143: douta=16'hbd54;
18144: douta=16'hbd54;
18145: douta=16'hb513;
18146: douta=16'h9cb3;
18147: douta=16'h9452;
18148: douta=16'h8c31;
18149: douta=16'h8411;
18150: douta=16'h83f1;
18151: douta=16'h7bd1;
18152: douta=16'h7bb0;
18153: douta=16'h736f;
18154: douta=16'h6b4f;
18155: douta=16'h528d;
18156: douta=16'h6aed;
18157: douta=16'hd592;
18158: douta=16'hde14;
18159: douta=16'hd5b3;
18160: douta=16'ha4d4;
18161: douta=16'h8c74;
18162: douta=16'h7c33;
18163: douta=16'h6370;
18164: douta=16'h52ce;
18165: douta=16'h5b0f;
18166: douta=16'h4aae;
18167: douta=16'h4aad;
18168: douta=16'h426c;
18169: douta=16'h3a2c;
18170: douta=16'h39ea;
18171: douta=16'h31eb;
18172: douta=16'h4a4b;
18173: douta=16'hac70;
18174: douta=16'h9494;
18175: douta=16'h424d;
18176: douta=16'h7414;
18177: douta=16'h42ae;
18178: douta=16'h3a6d;
18179: douta=16'h3a4e;
18180: douta=16'h3a8e;
18181: douta=16'h29cb;
18182: douta=16'h2a0b;
18183: douta=16'h324e;
18184: douta=16'h7414;
18185: douta=16'h1948;
18186: douta=16'h322c;
18187: douta=16'h2189;
18188: douta=16'h29ca;
18189: douta=16'h1907;
18190: douta=16'h2147;
18191: douta=16'h1968;
18192: douta=16'h10a4;
18193: douta=16'h10a4;
18194: douta=16'h10e5;
18195: douta=16'h1906;
18196: douta=16'h10c5;
18197: douta=16'h10e5;
18198: douta=16'h10e5;
18199: douta=16'h3a4c;
18200: douta=16'h63b3;
18201: douta=16'h4aef;
18202: douta=16'h5b31;
18203: douta=16'h428d;
18204: douta=16'h6391;
18205: douta=16'h6bd2;
18206: douta=16'h8454;
18207: douta=16'h5b71;
18208: douta=16'h5372;
18209: douta=16'h63d3;
18210: douta=16'h63b3;
18211: douta=16'h328e;
18212: douta=16'h4b31;
18213: douta=16'h42f0;
18214: douta=16'h5bb3;
18215: douta=16'h4332;
18216: douta=16'h5352;
18217: douta=16'hae3b;
18218: douta=16'h3189;
18219: douta=16'h628a;
18220: douta=16'h49e7;
18221: douta=16'h41a7;
18222: douta=16'h41e7;
18223: douta=16'h41a7;
18224: douta=16'h49c7;
18225: douta=16'h41a7;
18226: douta=16'h41a7;
18227: douta=16'h41c7;
18228: douta=16'h41a7;
18229: douta=16'h39a6;
18230: douta=16'h41a7;
18231: douta=16'h49e7;
18232: douta=16'h39a6;
18233: douta=16'h41a7;
18234: douta=16'h49e8;
18235: douta=16'h49c8;
18236: douta=16'h49c8;
18237: douta=16'h49e8;
18238: douta=16'h49c8;
18239: douta=16'h49e8;
18240: douta=16'hdd2b;
18241: douta=16'h8ba8;
18242: douta=16'h3965;
18243: douta=16'h30e3;
18244: douta=16'h28c2;
18245: douta=16'h3124;
18246: douta=16'h3145;
18247: douta=16'h3a2b;
18248: douta=16'h2187;
18249: douta=16'h1967;
18250: douta=16'h3a2b;
18251: douta=16'h3a0a;
18252: douta=16'h31e9;
18253: douta=16'h31a8;
18254: douta=16'h422a;
18255: douta=16'h3a2a;
18256: douta=16'h424b;
18257: douta=16'h4aac;
18258: douta=16'h52cd;
18259: douta=16'h636f;
18260: douta=16'h6390;
18261: douta=16'h6370;
18262: douta=16'h636f;
18263: douta=16'h6bd0;
18264: douta=16'h6bb0;
18265: douta=16'h6bf1;
18266: douta=16'h5b2e;
18267: douta=16'h636f;
18268: douta=16'h636e;
18269: douta=16'h5b6e;
18270: douta=16'h5b6e;
18271: douta=16'h638f;
18272: douta=16'h638e;
18273: douta=16'h638e;
18274: douta=16'h5b2d;
18275: douta=16'h530c;
18276: douta=16'h530d;
18277: douta=16'h4acb;
18278: douta=16'h4acb;
18279: douta=16'h4acb;
18280: douta=16'h736e;
18281: douta=16'h4a8c;
18282: douta=16'hff37;
18283: douta=16'heeb6;
18284: douta=16'heeb6;
18285: douta=16'heeb7;
18286: douta=16'heeb6;
18287: douta=16'heed7;
18288: douta=16'hcd93;
18289: douta=16'hd5d4;
18290: douta=16'hc573;
18291: douta=16'hb4f3;
18292: douta=16'hb514;
18293: douta=16'had14;
18294: douta=16'ha4f4;
18295: douta=16'h8433;
18296: douta=16'h8412;
18297: douta=16'h7bd1;
18298: douta=16'h6b4f;
18299: douta=16'h6b2e;
18300: douta=16'h630d;
18301: douta=16'h62cd;
18302: douta=16'h72ca;
18303: douta=16'hc50d;
18304: douta=16'he633;
18305: douta=16'hddf2;
18306: douta=16'heeb6;
18307: douta=16'hddf2;
18308: douta=16'h83d0;
18309: douta=16'h5aee;
18310: douta=16'hb490;
18311: douta=16'h9c91;
18312: douta=16'h83d1;
18313: douta=16'h83f2;
18314: douta=16'h83d1;
18315: douta=16'h8c11;
18316: douta=16'h83af;
18317: douta=16'h7b8f;
18318: douta=16'h736e;
18319: douta=16'h6aec;
18320: douta=16'h62ed;
18321: douta=16'h422a;
18322: douta=16'h524c;
18323: douta=16'h9bec;
18324: douta=16'hc4ae;
18325: douta=16'hee96;
18326: douta=16'hf6d7;
18327: douta=16'hcd51;
18328: douta=16'hde35;
18329: douta=16'hde13;
18330: douta=16'hd592;
18331: douta=16'h8c53;
18332: douta=16'h9453;
18333: douta=16'h9c93;
18334: douta=16'h9432;
18335: douta=16'h9452;
18336: douta=16'h8c32;
18337: douta=16'h8c31;
18338: douta=16'h9472;
18339: douta=16'ha4d4;
18340: douta=16'h8c11;
18341: douta=16'h8432;
18342: douta=16'h9453;
18343: douta=16'h7bcf;
18344: douta=16'h736e;
18345: douta=16'h6aee;
18346: douta=16'hd5b3;
18347: douta=16'heeb5;
18348: douta=16'he655;
18349: douta=16'hbd34;
18350: douta=16'hacd4;
18351: douta=16'h9494;
18352: douta=16'h8c53;
18353: douta=16'h8433;
18354: douta=16'h73d1;
18355: douta=16'h5aee;
18356: douta=16'h630e;
18357: douta=16'h632f;
18358: douta=16'h4a8d;
18359: douta=16'h4a8d;
18360: douta=16'h4a8d;
18361: douta=16'h3a4c;
18362: douta=16'h29a9;
18363: douta=16'h39ea;
18364: douta=16'hacb2;
18365: douta=16'h7bd2;
18366: douta=16'h734f;
18367: douta=16'h6350;
18368: douta=16'h5b50;
18369: douta=16'h4ace;
18370: douta=16'h3a6c;
18371: douta=16'h3a4c;
18372: douta=16'h2a0c;
18373: douta=16'h2a0c;
18374: douta=16'h21cb;
18375: douta=16'h7bd1;
18376: douta=16'h5331;
18377: douta=16'h3a4d;
18378: douta=16'h4aef;
18379: douta=16'h42ce;
18380: douta=16'h320c;
18381: douta=16'h320c;
18382: douta=16'h2989;
18383: douta=16'h10e5;
18384: douta=16'h320b;
18385: douta=16'h29ca;
18386: douta=16'h10c4;
18387: douta=16'h18e5;
18388: douta=16'h10c5;
18389: douta=16'h10e5;
18390: douta=16'h1906;
18391: douta=16'h18e5;
18392: douta=16'h0884;
18393: douta=16'h5330;
18394: douta=16'h29a9;
18395: douta=16'h6bb1;
18396: douta=16'h42ce;
18397: douta=16'h6bf2;
18398: douta=16'h5b72;
18399: douta=16'h5b72;
18400: douta=16'h7c56;
18401: douta=16'h5b72;
18402: douta=16'h63b3;
18403: douta=16'h5bb3;
18404: douta=16'h4b31;
18405: douta=16'h6bd3;
18406: douta=16'h6c36;
18407: douta=16'h6c56;
18408: douta=16'h53f6;
18409: douta=16'h94f5;
18410: douta=16'hadda;
18411: douta=16'h11cb;
18412: douta=16'h5a27;
18413: douta=16'h5227;
18414: douta=16'h49c8;
18415: douta=16'h41a7;
18416: douta=16'h49c7;
18417: douta=16'h4186;
18418: douta=16'h41a7;
18419: douta=16'h41a7;
18420: douta=16'h41a7;
18421: douta=16'h39a6;
18422: douta=16'h41a7;
18423: douta=16'h41a7;
18424: douta=16'h49e7;
18425: douta=16'h4a08;
18426: douta=16'h49e8;
18427: douta=16'h49e8;
18428: douta=16'h49e8;
18429: douta=16'h49e8;
18430: douta=16'h49e8;
18431: douta=16'h5208;
18432: douta=16'hdd2b;
18433: douta=16'hac68;
18434: douta=16'h3944;
18435: douta=16'h30e3;
18436: douta=16'h30e2;
18437: douta=16'h3144;
18438: douta=16'h3124;
18439: douta=16'h3a0a;
18440: douta=16'h1946;
18441: douta=16'h2147;
18442: douta=16'h320b;
18443: douta=16'h3a0a;
18444: douta=16'h31c9;
18445: douta=16'h31a8;
18446: douta=16'h39e9;
18447: douta=16'h3a0a;
18448: douta=16'h426c;
18449: douta=16'h4aad;
18450: douta=16'h4aac;
18451: douta=16'h5b2f;
18452: douta=16'h636f;
18453: douta=16'h6370;
18454: douta=16'h6390;
18455: douta=16'h6bb1;
18456: douta=16'h6bd1;
18457: douta=16'h6390;
18458: douta=16'h532e;
18459: douta=16'h532e;
18460: douta=16'h5b2e;
18461: douta=16'h5b4e;
18462: douta=16'h532e;
18463: douta=16'h532d;
18464: douta=16'h5b4e;
18465: douta=16'h4aec;
18466: douta=16'h52ec;
18467: douta=16'h4acb;
18468: douta=16'h4acc;
18469: douta=16'h4acb;
18470: douta=16'h52ec;
18471: douta=16'h52ec;
18472: douta=16'h52ec;
18473: douta=16'h4aac;
18474: douta=16'hf696;
18475: douta=16'heeb7;
18476: douta=16'heed7;
18477: douta=16'heeb7;
18478: douta=16'heed7;
18479: douta=16'hee96;
18480: douta=16'hc572;
18481: douta=16'hd5b4;
18482: douta=16'hcd73;
18483: douta=16'had14;
18484: douta=16'h9c92;
18485: douta=16'h9cb4;
18486: douta=16'ha4f4;
18487: douta=16'h9473;
18488: douta=16'h8c74;
18489: douta=16'h8411;
18490: douta=16'h738f;
18491: douta=16'h734e;
18492: douta=16'h6b4e;
18493: douta=16'h4168;
18494: douta=16'hc4cc;
18495: douta=16'hddf3;
18496: douta=16'hf6d7;
18497: douta=16'he675;
18498: douta=16'he675;
18499: douta=16'hcd71;
18500: douta=16'h6b6e;
18501: douta=16'h6b70;
18502: douta=16'hc511;
18503: douta=16'h9452;
18504: douta=16'h9432;
18505: douta=16'h83f2;
18506: douta=16'h7bb0;
18507: douta=16'h83b0;
18508: douta=16'h83af;
18509: douta=16'h7b8f;
18510: douta=16'h7b8f;
18511: douta=16'h6aec;
18512: douta=16'h62ab;
18513: douta=16'h422b;
18514: douta=16'hac0d;
18515: douta=16'hddb0;
18516: douta=16'he633;
18517: douta=16'he696;
18518: douta=16'hcd72;
18519: douta=16'hd5f4;
18520: douta=16'hcd52;
18521: douta=16'hc554;
18522: douta=16'hc532;
18523: douta=16'ha4d3;
18524: douta=16'h8433;
18525: douta=16'h7bf2;
18526: douta=16'h9453;
18527: douta=16'h9451;
18528: douta=16'h9432;
18529: douta=16'h83d0;
18530: douta=16'h9451;
18531: douta=16'h9c52;
18532: douta=16'h9c93;
18533: douta=16'h8c30;
18534: douta=16'h8c11;
18535: douta=16'h6acc;
18536: douta=16'h7b6e;
18537: douta=16'hbd12;
18538: douta=16'heeb6;
18539: douta=16'hd5d4;
18540: douta=16'hd5d5;
18541: douta=16'hbd35;
18542: douta=16'hb515;
18543: douta=16'h94b5;
18544: douta=16'h8432;
18545: douta=16'h7bd1;
18546: douta=16'h7390;
18547: douta=16'h632e;
18548: douta=16'h630e;
18549: douta=16'h6b50;
18550: douta=16'h4aad;
18551: douta=16'h4aad;
18552: douta=16'h4a6d;
18553: douta=16'h3a0b;
18554: douta=16'h5aed;
18555: douta=16'h9c52;
18556: douta=16'h8c13;
18557: douta=16'h7bd2;
18558: douta=16'h736f;
18559: douta=16'h5b2f;
18560: douta=16'h530f;
18561: douta=16'h4aad;
18562: douta=16'h428d;
18563: douta=16'h3a2c;
18564: douta=16'h322b;
18565: douta=16'h21aa;
18566: douta=16'h630e;
18567: douta=16'hacd4;
18568: douta=16'h5351;
18569: douta=16'h4aaf;
18570: douta=16'h5310;
18571: douta=16'h4acf;
18572: douta=16'h324d;
18573: douta=16'h322c;
18574: douta=16'h2189;
18575: douta=16'h1947;
18576: douta=16'h21a9;
18577: douta=16'h4af0;
18578: douta=16'h10e5;
18579: douta=16'h1083;
18580: douta=16'h10c5;
18581: douta=16'h10e5;
18582: douta=16'h1905;
18583: douta=16'h10e5;
18584: douta=16'h10c4;
18585: douta=16'h1906;
18586: douta=16'h0884;
18587: douta=16'h8cd6;
18588: douta=16'h5b2f;
18589: douta=16'h7414;
18590: douta=16'h42ce;
18591: douta=16'h7414;
18592: douta=16'h73f4;
18593: douta=16'h428f;
18594: douta=16'h5b92;
18595: douta=16'h5352;
18596: douta=16'h5bd4;
18597: douta=16'h7456;
18598: douta=16'h5bd5;
18599: douta=16'h6c56;
18600: douta=16'h6c57;
18601: douta=16'h74f9;
18602: douta=16'hc67a;
18603: douta=16'h74f9;
18604: douta=16'h21ea;
18605: douta=16'h41c7;
18606: douta=16'h49e7;
18607: douta=16'h49c7;
18608: douta=16'h49e7;
18609: douta=16'h41a7;
18610: douta=16'h49a7;
18611: douta=16'h41c7;
18612: douta=16'h41a7;
18613: douta=16'h39a6;
18614: douta=16'h49e8;
18615: douta=16'h49e7;
18616: douta=16'h49e8;
18617: douta=16'h5229;
18618: douta=16'h49c8;
18619: douta=16'h49e8;
18620: douta=16'h49e8;
18621: douta=16'h49e8;
18622: douta=16'h49e8;
18623: douta=16'h5228;
18624: douta=16'hdd4c;
18625: douta=16'hf5ec;
18626: douta=16'h20a3;
18627: douta=16'h3965;
18628: douta=16'h52cb;
18629: douta=16'h30c2;
18630: douta=16'h3124;
18631: douta=16'h3125;
18632: douta=16'h1967;
18633: douta=16'h2167;
18634: douta=16'h29a9;
18635: douta=16'h29a9;
18636: douta=16'h2968;
18637: douta=16'h2988;
18638: douta=16'h29a8;
18639: douta=16'h2987;
18640: douta=16'h3a4b;
18641: douta=16'h426c;
18642: douta=16'h428c;
18643: douta=16'h4aad;
18644: douta=16'h52ee;
18645: douta=16'h5b4f;
18646: douta=16'h5b4f;
18647: douta=16'h636f;
18648: douta=16'h6bd1;
18649: douta=16'h6bf1;
18650: douta=16'h5b4e;
18651: douta=16'h5b4e;
18652: douta=16'h636f;
18653: douta=16'h5b2e;
18654: douta=16'h5b4e;
18655: douta=16'h5b6f;
18656: douta=16'h63af;
18657: douta=16'h532d;
18658: douta=16'h4aab;
18659: douta=16'h428b;
18660: douta=16'h4acb;
18661: douta=16'h5b2e;
18662: douta=16'h52ed;
18663: douta=16'h530d;
18664: douta=16'h4acc;
18665: douta=16'h530c;
18666: douta=16'h5b6e;
18667: douta=16'hddb4;
18668: douta=16'hee76;
18669: douta=16'hee96;
18670: douta=16'heeb6;
18671: douta=16'hde35;
18672: douta=16'hcdb3;
18673: douta=16'ha4b3;
18674: douta=16'hacd3;
18675: douta=16'hbd55;
18676: douta=16'ha4d5;
18677: douta=16'ha515;
18678: douta=16'ha4d5;
18679: douta=16'h7bd1;
18680: douta=16'h738f;
18681: douta=16'h738f;
18682: douta=16'h83f1;
18683: douta=16'h3146;
18684: douta=16'h59c5;
18685: douta=16'hee75;
18686: douta=16'hee76;
18687: douta=16'heed7;
18688: douta=16'he675;
18689: douta=16'he675;
18690: douta=16'hd5d3;
18691: douta=16'hd593;
18692: douta=16'ha4b2;
18693: douta=16'h8c53;
18694: douta=16'h3aaf;
18695: douta=16'h62cc;
18696: douta=16'h8c11;
18697: douta=16'h736f;
18698: douta=16'h736f;
18699: douta=16'h62ec;
18700: douta=16'h6b2d;
18701: douta=16'h62cc;
18702: douta=16'h6b0d;
18703: douta=16'h62cd;
18704: douta=16'h72eb;
18705: douta=16'hd52f;
18706: douta=16'he675;
18707: douta=16'hee98;
18708: douta=16'hee96;
18709: douta=16'hde35;
18710: douta=16'hcd94;
18711: douta=16'h8452;
18712: douta=16'ha4b3;
18713: douta=16'ha493;
18714: douta=16'ha4d4;
18715: douta=16'h8c32;
18716: douta=16'h9453;
18717: douta=16'h8c72;
18718: douta=16'h5330;
18719: douta=16'h5330;
18720: douta=16'h5b2f;
18721: douta=16'h736f;
18722: douta=16'h632d;
18723: douta=16'h528c;
18724: douta=16'h7b6d;
18725: douta=16'hac70;
18726: douta=16'hf6d6;
18727: douta=16'hee97;
18728: douta=16'hf6b6;
18729: douta=16'hddf5;
18730: douta=16'h9c94;
18731: douta=16'h9473;
18732: douta=16'h9454;
18733: douta=16'h9474;
18734: douta=16'h8c53;
18735: douta=16'h8412;
18736: douta=16'h7bd1;
18737: douta=16'h7b90;
18738: douta=16'h736f;
18739: douta=16'h732e;
18740: douta=16'h630d;
18741: douta=16'h630e;
18742: douta=16'h426b;
18743: douta=16'h528c;
18744: douta=16'h9432;
18745: douta=16'hb4f4;
18746: douta=16'h9452;
18747: douta=16'h8c32;
18748: douta=16'h7390;
18749: douta=16'h7390;
18750: douta=16'h630e;
18751: douta=16'h5aee;
18752: douta=16'h52cd;
18753: douta=16'h4aad;
18754: douta=16'h428d;
18755: douta=16'h320b;
18756: douta=16'h3a2b;
18757: douta=16'h8433;
18758: douta=16'h7c12;
18759: douta=16'h7bd2;
18760: douta=16'h5b0f;
18761: douta=16'h4ace;
18762: douta=16'h42ce;
18763: douta=16'h428e;
18764: douta=16'h3a6d;
18765: douta=16'h322c;
18766: douta=16'h29a9;
18767: douta=16'h2188;
18768: douta=16'h42ae;
18769: douta=16'h426d;
18770: douta=16'h29eb;
18771: douta=16'h29ca;
18772: douta=16'h10e5;
18773: douta=16'h10e5;
18774: douta=16'h10c4;
18775: douta=16'h10e5;
18776: douta=16'h10c4;
18777: douta=16'h10c4;
18778: douta=16'h1906;
18779: douta=16'h10e6;
18780: douta=16'h4acd;
18781: douta=16'h7414;
18782: douta=16'h7c75;
18783: douta=16'h5b71;
18784: douta=16'h5351;
18785: douta=16'h84d8;
18786: douta=16'h7456;
18787: douta=16'h5bb4;
18788: douta=16'h63f5;
18789: douta=16'h6c15;
18790: douta=16'h5bd5;
18791: douta=16'h6c77;
18792: douta=16'h7cd9;
18793: douta=16'h6416;
18794: douta=16'h53d4;
18795: douta=16'h6c57;
18796: douta=16'h9579;
18797: douta=16'h7d39;
18798: douta=16'h8d9b;
18799: douta=16'h422a;
18800: douta=16'h4165;
18801: douta=16'h41a6;
18802: douta=16'h41a6;
18803: douta=16'h49a7;
18804: douta=16'h41a7;
18805: douta=16'h49e7;
18806: douta=16'h5208;
18807: douta=16'h5208;
18808: douta=16'h5208;
18809: douta=16'h5229;
18810: douta=16'h5208;
18811: douta=16'h5228;
18812: douta=16'h5249;
18813: douta=16'h4a08;
18814: douta=16'h5229;
18815: douta=16'h5229;
18816: douta=16'hdd4b;
18817: douta=16'hed8b;
18818: douta=16'h41c5;
18819: douta=16'h3945;
18820: douta=16'h6b90;
18821: douta=16'h3124;
18822: douta=16'h3124;
18823: douta=16'h2904;
18824: douta=16'h2168;
18825: douta=16'h1926;
18826: douta=16'h29a9;
18827: douta=16'h29a9;
18828: douta=16'h29c9;
18829: douta=16'h2968;
18830: douta=16'h320b;
18831: douta=16'h3a4c;
18832: douta=16'h3a4c;
18833: douta=16'h3a4b;
18834: douta=16'h426c;
18835: douta=16'h52ee;
18836: douta=16'h5b2f;
18837: douta=16'h530e;
18838: douta=16'h530e;
18839: douta=16'h4aed;
18840: douta=16'h530e;
18841: douta=16'h5b4f;
18842: douta=16'h532e;
18843: douta=16'h5b4e;
18844: douta=16'h534e;
18845: douta=16'h5b4e;
18846: douta=16'h5b4e;
18847: douta=16'h5b6f;
18848: douta=16'h638f;
18849: douta=16'h5b6f;
18850: douta=16'h530d;
18851: douta=16'h4acc;
18852: douta=16'h4acc;
18853: douta=16'h4acc;
18854: douta=16'h530d;
18855: douta=16'h428b;
18856: douta=16'h52ec;
18857: douta=16'h530c;
18858: douta=16'h530d;
18859: douta=16'h530c;
18860: douta=16'hacb1;
18861: douta=16'he614;
18862: douta=16'hde35;
18863: douta=16'hd5f4;
18864: douta=16'hc5b4;
18865: douta=16'hb514;
18866: douta=16'ha4d4;
18867: douta=16'h9cb5;
18868: douta=16'ha515;
18869: douta=16'h9cd4;
18870: douta=16'h94b4;
18871: douta=16'h738e;
18872: douta=16'h734e;
18873: douta=16'h734e;
18874: douta=16'h49a5;
18875: douta=16'he5d1;
18876: douta=16'hcd0d;
18877: douta=16'he613;
18878: douta=16'heed7;
18879: douta=16'heeb7;
18880: douta=16'hde34;
18881: douta=16'he635;
18882: douta=16'hcd73;
18883: douta=16'hbd52;
18884: douta=16'h9cb3;
18885: douta=16'h8c73;
18886: douta=16'h8473;
18887: douta=16'h6bd3;
18888: douta=16'h31ea;
18889: douta=16'h732d;
18890: douta=16'h6b0d;
18891: douta=16'h6b0d;
18892: douta=16'h62cc;
18893: douta=16'h5a8b;
18894: douta=16'h4a2a;
18895: douta=16'hd52e;
18896: douta=16'he612;
18897: douta=16'heeb6;
18898: douta=16'hac70;
18899: douta=16'hee96;
18900: douta=16'hde54;
18901: douta=16'hbd54;
18902: douta=16'hb514;
18903: douta=16'hb515;
18904: douta=16'h9473;
18905: douta=16'hacd4;
18906: douta=16'ha4b4;
18907: douta=16'h8411;
18908: douta=16'h8412;
18909: douta=16'h8c12;
18910: douta=16'h7b8f;
18911: douta=16'h7baf;
18912: douta=16'h734e;
18913: douta=16'h62ed;
18914: douta=16'h93ee;
18915: douta=16'hb4b1;
18916: douta=16'hb4d3;
18917: douta=16'hc553;
18918: douta=16'hd5f4;
18919: douta=16'hacd3;
18920: douta=16'h9c53;
18921: douta=16'h9453;
18922: douta=16'h9c93;
18923: douta=16'ha4d4;
18924: douta=16'ha4b4;
18925: douta=16'h8432;
18926: douta=16'h8432;
18927: douta=16'h83f1;
18928: douta=16'h7bb0;
18929: douta=16'h734e;
18930: douta=16'h6b0d;
18931: douta=16'h6b0e;
18932: douta=16'h62ac;
18933: douta=16'h6aed;
18934: douta=16'ha4b4;
18935: douta=16'ha493;
18936: douta=16'h9cb3;
18937: douta=16'h9453;
18938: douta=16'h83d1;
18939: douta=16'h83d0;
18940: douta=16'h736f;
18941: douta=16'h630e;
18942: douta=16'h630e;
18943: douta=16'h5acd;
18944: douta=16'h52ad;
18945: douta=16'h4a8c;
18946: douta=16'h630d;
18947: douta=16'hacd4;
18948: douta=16'ha4b5;
18949: douta=16'h8c33;
18950: douta=16'h8452;
18951: douta=16'h8413;
18952: douta=16'h632f;
18953: douta=16'h4a8d;
18954: douta=16'h4a8d;
18955: douta=16'h4aad;
18956: douta=16'h3a4d;
18957: douta=16'h320b;
18958: douta=16'h3a2b;
18959: douta=16'h5b72;
18960: douta=16'h6b4e;
18961: douta=16'h3a4e;
18962: douta=16'h530f;
18963: douta=16'h5310;
18964: douta=16'h2168;
18965: douta=16'h29aa;
18966: douta=16'h18e6;
18967: douta=16'h18e5;
18968: douta=16'h08c4;
18969: douta=16'h10e5;
18970: douta=16'h10e5;
18971: douta=16'h10e6;
18972: douta=16'h1107;
18973: douta=16'h6bb3;
18974: douta=16'h6bf3;
18975: douta=16'h7c75;
18976: douta=16'h9d59;
18977: douta=16'h7435;
18978: douta=16'h63f5;
18979: douta=16'h63f5;
18980: douta=16'h6c56;
18981: douta=16'h7456;
18982: douta=16'h5bf5;
18983: douta=16'h7497;
18984: douta=16'h5bd4;
18985: douta=16'h6c77;
18986: douta=16'h5bd4;
18987: douta=16'h53b4;
18988: douta=16'h6436;
18989: douta=16'h74b8;
18990: douta=16'h53f6;
18991: douta=16'h7c97;
18992: douta=16'h959c;
18993: douta=16'h73f3;
18994: douta=16'h49e7;
18995: douta=16'h49e7;
18996: douta=16'h49e7;
18997: douta=16'h5228;
18998: douta=16'h5208;
18999: douta=16'h5229;
19000: douta=16'h5228;
19001: douta=16'h5208;
19002: douta=16'h5228;
19003: douta=16'h5208;
19004: douta=16'h5208;
19005: douta=16'h5208;
19006: douta=16'h5208;
19007: douta=16'h5228;
19008: douta=16'hdd4c;
19009: douta=16'he54b;
19010: douta=16'h6265;
19011: douta=16'h3965;
19012: douta=16'h6b6f;
19013: douta=16'h41a6;
19014: douta=16'h3944;
19015: douta=16'h2904;
19016: douta=16'h2988;
19017: douta=16'h1946;
19018: douta=16'h29a9;
19019: douta=16'h2168;
19020: douta=16'h2988;
19021: douta=16'h2988;
19022: douta=16'h3a2c;
19023: douta=16'h3a6c;
19024: douta=16'h3a4c;
19025: douta=16'h322b;
19026: douta=16'h3a2b;
19027: douta=16'h530e;
19028: douta=16'h532e;
19029: douta=16'h530e;
19030: douta=16'h530e;
19031: douta=16'h4aed;
19032: douta=16'h532e;
19033: douta=16'h638f;
19034: douta=16'h530e;
19035: douta=16'h532d;
19036: douta=16'h534e;
19037: douta=16'h534e;
19038: douta=16'h5b4e;
19039: douta=16'h5b6f;
19040: douta=16'h638f;
19041: douta=16'h5b6e;
19042: douta=16'h5b4e;
19043: douta=16'h5b2d;
19044: douta=16'h4acc;
19045: douta=16'h530d;
19046: douta=16'h52ec;
19047: douta=16'h52ec;
19048: douta=16'h4aab;
19049: douta=16'h4acc;
19050: douta=16'h4acb;
19051: douta=16'h5b4d;
19052: douta=16'h4aed;
19053: douta=16'h7b8f;
19054: douta=16'hddf4;
19055: douta=16'hcdb3;
19056: douta=16'hb533;
19057: douta=16'hb535;
19058: douta=16'hacf4;
19059: douta=16'ha4d4;
19060: douta=16'h9453;
19061: douta=16'h9493;
19062: douta=16'h8c53;
19063: douta=16'h736e;
19064: douta=16'h736e;
19065: douta=16'h62cc;
19066: douta=16'h8ae7;
19067: douta=16'hee73;
19068: douta=16'hc50e;
19069: douta=16'hddb1;
19070: douta=16'heeb7;
19071: douta=16'he676;
19072: douta=16'hde35;
19073: douta=16'hd5f3;
19074: douta=16'hbd13;
19075: douta=16'hacd3;
19076: douta=16'h9473;
19077: douta=16'h8c53;
19078: douta=16'h8412;
19079: douta=16'h5b2e;
19080: douta=16'h424c;
19081: douta=16'h7b4e;
19082: douta=16'h7b6e;
19083: douta=16'h6b2c;
19084: douta=16'h6aec;
19085: douta=16'h524b;
19086: douta=16'h628b;
19087: douta=16'he614;
19088: douta=16'heeb6;
19089: douta=16'hde55;
19090: douta=16'ha4b3;
19091: douta=16'hde14;
19092: douta=16'hcd54;
19093: douta=16'had14;
19094: douta=16'hacf4;
19095: douta=16'had15;
19096: douta=16'h7bf1;
19097: douta=16'h8c33;
19098: douta=16'h9c93;
19099: douta=16'h83d1;
19100: douta=16'h83d0;
19101: douta=16'h83f1;
19102: douta=16'h736e;
19103: douta=16'h7b8f;
19104: douta=16'h736e;
19105: douta=16'h7b4d;
19106: douta=16'hf696;
19107: douta=16'hee96;
19108: douta=16'h9434;
19109: douta=16'hcd74;
19110: douta=16'hde15;
19111: douta=16'hbd55;
19112: douta=16'hb535;
19113: douta=16'h9452;
19114: douta=16'h8c11;
19115: douta=16'h8c11;
19116: douta=16'h8c11;
19117: douta=16'h83d0;
19118: douta=16'h7b90;
19119: douta=16'h7bb0;
19120: douta=16'h736f;
19121: douta=16'h7b6f;
19122: douta=16'h734e;
19123: douta=16'h528c;
19124: douta=16'h7b8f;
19125: douta=16'hacd4;
19126: douta=16'h9cb3;
19127: douta=16'h9472;
19128: douta=16'h8c32;
19129: douta=16'h8412;
19130: douta=16'h7bb0;
19131: douta=16'h7bb0;
19132: douta=16'h736f;
19133: douta=16'h6b2e;
19134: douta=16'h630e;
19135: douta=16'h52cd;
19136: douta=16'h52ad;
19137: douta=16'h528d;
19138: douta=16'hcd94;
19139: douta=16'ha4d3;
19140: douta=16'h9c94;
19141: douta=16'h8433;
19142: douta=16'h7bf2;
19143: douta=16'h7390;
19144: douta=16'h5b2f;
19145: douta=16'h52ce;
19146: douta=16'h4ace;
19147: douta=16'h426d;
19148: douta=16'h428d;
19149: douta=16'h428d;
19150: douta=16'h322d;
19151: douta=16'h426d;
19152: douta=16'hc5b7;
19153: douta=16'h428e;
19154: douta=16'h6bb1;
19155: douta=16'h5b30;
19156: douta=16'h29a9;
19157: douta=16'h2168;
19158: douta=16'h31ca;
19159: douta=16'h1083;
19160: douta=16'h10e5;
19161: douta=16'h18e5;
19162: douta=16'h1905;
19163: douta=16'h10e5;
19164: douta=16'h10e6;
19165: douta=16'h84b6;
19166: douta=16'h7c75;
19167: douta=16'h7435;
19168: douta=16'h63f4;
19169: douta=16'h5bb4;
19170: douta=16'h6c35;
19171: douta=16'h84b7;
19172: douta=16'h9559;
19173: douta=16'h63f4;
19174: douta=16'h84d8;
19175: douta=16'h4b73;
19176: douta=16'h5bd4;
19177: douta=16'h6415;
19178: douta=16'h5bd5;
19179: douta=16'h5394;
19180: douta=16'h6c56;
19181: douta=16'h6477;
19182: douta=16'h6cb9;
19183: douta=16'h1948;
19184: douta=16'h5b70;
19185: douta=16'h6c55;
19186: douta=16'h49c7;
19187: douta=16'h49e8;
19188: douta=16'h5208;
19189: douta=16'h5208;
19190: douta=16'h5229;
19191: douta=16'h5229;
19192: douta=16'h4a08;
19193: douta=16'h5228;
19194: douta=16'h49e8;
19195: douta=16'h49e8;
19196: douta=16'h5228;
19197: douta=16'h49e8;
19198: douta=16'h5208;
19199: douta=16'h5208;
19200: douta=16'he56c;
19201: douta=16'hdd4b;
19202: douta=16'hccea;
19203: douta=16'h3945;
19204: douta=16'h5acb;
19205: douta=16'h6b6f;
19206: douta=16'h3945;
19207: douta=16'h3124;
19208: douta=16'h10a3;
19209: douta=16'h10c4;
19210: douta=16'h1083;
19211: douta=16'h1083;
19212: douta=16'h10a3;
19213: douta=16'h1906;
19214: douta=16'h320b;
19215: douta=16'h31eb;
19216: douta=16'h3a2c;
19217: douta=16'h31ea;
19218: douta=16'h320b;
19219: douta=16'h428d;
19220: douta=16'h42ad;
19221: douta=16'h4aee;
19222: douta=16'h532f;
19223: douta=16'h532f;
19224: douta=16'h530e;
19225: douta=16'h532f;
19226: douta=16'h42cd;
19227: douta=16'h4aed;
19228: douta=16'h4b0d;
19229: douta=16'h532e;
19230: douta=16'h532e;
19231: douta=16'h532e;
19232: douta=16'h532e;
19233: douta=16'h4b0d;
19234: douta=16'h530d;
19235: douta=16'h4aac;
19236: douta=16'h52ed;
19237: douta=16'h530d;
19238: douta=16'h5b2e;
19239: douta=16'h5b4e;
19240: douta=16'h638f;
19241: douta=16'h638f;
19242: douta=16'h638f;
19243: douta=16'h636f;
19244: douta=16'h63d0;
19245: douta=16'h63b0;
19246: douta=16'h5bb0;
19247: douta=16'h638f;
19248: douta=16'h9c50;
19249: douta=16'ha491;
19250: douta=16'ha492;
19251: douta=16'h8c51;
19252: douta=16'h7bb0;
19253: douta=16'h736e;
19254: douta=16'h732e;
19255: douta=16'h4a0a;
19256: douta=16'h6a8a;
19257: douta=16'hd52f;
19258: douta=16'heeb7;
19259: douta=16'he634;
19260: douta=16'hf6f7;
19261: douta=16'hac4e;
19262: douta=16'hee75;
19263: douta=16'hcd92;
19264: douta=16'hcd73;
19265: douta=16'hc532;
19266: douta=16'hb514;
19267: douta=16'h9cb3;
19268: douta=16'h8c73;
19269: douta=16'h8452;
19270: douta=16'h73b0;
19271: douta=16'h6b6e;
19272: douta=16'h734e;
19273: douta=16'h6b0d;
19274: douta=16'h6acd;
19275: douta=16'h5aac;
19276: douta=16'ha3cb;
19277: douta=16'hddf3;
19278: douta=16'heeb6;
19279: douta=16'hee96;
19280: douta=16'hde14;
19281: douta=16'hbd74;
19282: douta=16'h8c34;
19283: douta=16'ha4f4;
19284: douta=16'hacf5;
19285: douta=16'h632f;
19286: douta=16'h8c31;
19287: douta=16'h83d0;
19288: douta=16'h8bf1;
19289: douta=16'h8bf1;
19290: douta=16'h732e;
19291: douta=16'h83f0;
19292: douta=16'h83b0;
19293: douta=16'h83d0;
19294: douta=16'h8bce;
19295: douta=16'hbcd0;
19296: douta=16'hf6b5;
19297: douta=16'he636;
19298: douta=16'hbd12;
19299: douta=16'hc533;
19300: douta=16'h8454;
19301: douta=16'h5b10;
19302: douta=16'ha4b3;
19303: douta=16'h8bf2;
19304: douta=16'h8bf1;
19305: douta=16'h8bf0;
19306: douta=16'h7b8e;
19307: douta=16'h7b8e;
19308: douta=16'h7b6e;
19309: douta=16'h732d;
19310: douta=16'h732d;
19311: douta=16'h6aec;
19312: douta=16'h8bd0;
19313: douta=16'had14;
19314: douta=16'hb535;
19315: douta=16'h83f1;
19316: douta=16'h8c32;
19317: douta=16'h8c32;
19318: douta=16'h83f1;
19319: douta=16'h7b90;
19320: douta=16'h7b90;
19321: douta=16'h736e;
19322: douta=16'h7bd0;
19323: douta=16'h7bb0;
19324: douta=16'h5ace;
19325: douta=16'h5aad;
19326: douta=16'h632e;
19327: douta=16'h9cb5;
19328: douta=16'h9474;
19329: douta=16'h8c53;
19330: douta=16'ha493;
19331: douta=16'h8c32;
19332: douta=16'h8c32;
19333: douta=16'h6b4e;
19334: douta=16'h6b4f;
19335: douta=16'h6b4f;
19336: douta=16'h630f;
19337: douta=16'h5aee;
19338: douta=16'h5acd;
19339: douta=16'h4a6c;
19340: douta=16'h4a8c;
19341: douta=16'h9451;
19342: douta=16'hb534;
19343: douta=16'h94b5;
19344: douta=16'h8434;
19345: douta=16'h7433;
19346: douta=16'h5330;
19347: douta=16'h4aae;
19348: douta=16'h29a9;
19349: douta=16'h320b;
19350: douta=16'h2189;
19351: douta=16'h18e5;
19352: douta=16'h428e;
19353: douta=16'h29c9;
19354: douta=16'h10e5;
19355: douta=16'h10e5;
19356: douta=16'h10e6;
19357: douta=16'h10c4;
19358: douta=16'h29a9;
19359: douta=16'h7496;
19360: douta=16'h9517;
19361: douta=16'h5394;
19362: douta=16'h6c15;
19363: douta=16'h63f4;
19364: douta=16'h6c55;
19365: douta=16'h9539;
19366: douta=16'h84b7;
19367: douta=16'h6c35;
19368: douta=16'h4b32;
19369: douta=16'h5bd4;
19370: douta=16'h7cb8;
19371: douta=16'h53d4;
19372: douta=16'h6457;
19373: douta=16'h6436;
19374: douta=16'h2188;
19375: douta=16'h29aa;
19376: douta=16'h29a9;
19377: douta=16'h29ca;
19378: douta=16'h2168;
19379: douta=16'h39e9;
19380: douta=16'h6aaa;
19381: douta=16'h5208;
19382: douta=16'h5a49;
19383: douta=16'h5229;
19384: douta=16'h49e8;
19385: douta=16'h5208;
19386: douta=16'h5249;
19387: douta=16'h4a08;
19388: douta=16'h5208;
19389: douta=16'h49e8;
19390: douta=16'h5208;
19391: douta=16'h49c7;
19392: douta=16'he56c;
19393: douta=16'he54c;
19394: douta=16'hedec;
19395: douta=16'h28e4;
19396: douta=16'h4985;
19397: douta=16'h7bd1;
19398: douta=16'h3903;
19399: douta=16'h28e3;
19400: douta=16'h10a3;
19401: douta=16'h10c4;
19402: douta=16'h2146;
19403: douta=16'h2146;
19404: douta=16'h2125;
19405: douta=16'h29ca;
19406: douta=16'h29ea;
19407: douta=16'h31eb;
19408: douta=16'h3a2b;
19409: douta=16'h29ea;
19410: douta=16'h3a4c;
19411: douta=16'h42ae;
19412: douta=16'h4ace;
19413: douta=16'h4aae;
19414: douta=16'h530f;
19415: douta=16'h530e;
19416: douta=16'h4aee;
19417: douta=16'h4b0e;
19418: douta=16'h3a6b;
19419: douta=16'h42ac;
19420: douta=16'h4b0d;
19421: douta=16'h530e;
19422: douta=16'h4b0d;
19423: douta=16'h534e;
19424: douta=16'h4aed;
19425: douta=16'h4b0d;
19426: douta=16'h52ed;
19427: douta=16'h4acc;
19428: douta=16'h4aac;
19429: douta=16'h4aac;
19430: douta=16'h4aac;
19431: douta=16'h52ed;
19432: douta=16'h5b4e;
19433: douta=16'h636f;
19434: douta=16'h638f;
19435: douta=16'h6bf0;
19436: douta=16'h63d0;
19437: douta=16'h63af;
19438: douta=16'h63d0;
19439: douta=16'h63d0;
19440: douta=16'h5bb0;
19441: douta=16'h6bb0;
19442: douta=16'h7bd0;
19443: douta=16'h9451;
19444: douta=16'h8c11;
19445: douta=16'h6b2d;
19446: douta=16'h6b2d;
19447: douta=16'hd54f;
19448: douta=16'hbcae;
19449: douta=16'hee95;
19450: douta=16'hcd50;
19451: douta=16'hf759;
19452: douta=16'heeb6;
19453: douta=16'h9410;
19454: douta=16'he675;
19455: douta=16'hc552;
19456: douta=16'ha4b3;
19457: douta=16'h9c93;
19458: douta=16'h83f2;
19459: douta=16'h7bf1;
19460: douta=16'h7bd1;
19461: douta=16'h7bb0;
19462: douta=16'h732e;
19463: douta=16'h6b2d;
19464: douta=16'h62ec;
19465: douta=16'h5aac;
19466: douta=16'h4a4b;
19467: douta=16'h9b6b;
19468: douta=16'hee76;
19469: douta=16'he674;
19470: douta=16'he635;
19471: douta=16'hbd53;
19472: douta=16'hbd54;
19473: douta=16'ha4d5;
19474: douta=16'ha516;
19475: douta=16'h8c94;
19476: douta=16'h7c33;
19477: douta=16'h94b3;
19478: douta=16'h632f;
19479: douta=16'h4ace;
19480: douta=16'h7b6f;
19481: douta=16'h838f;
19482: douta=16'h8bd0;
19483: douta=16'h62ed;
19484: douta=16'h5a6c;
19485: douta=16'h8b6d;
19486: douta=16'hacb2;
19487: douta=16'he655;
19488: douta=16'hcd93;
19489: douta=16'h5b50;
19490: douta=16'h8453;
19491: douta=16'h8c95;
19492: douta=16'h8454;
19493: douta=16'h6b91;
19494: douta=16'h5b50;
19495: douta=16'h83f1;
19496: douta=16'h9430;
19497: douta=16'h83ae;
19498: douta=16'h730d;
19499: douta=16'h6aec;
19500: douta=16'h6aec;
19501: douta=16'h8bf0;
19502: douta=16'h8c11;
19503: douta=16'h73d0;
19504: douta=16'h7bf2;
19505: douta=16'h8412;
19506: douta=16'h8bf1;
19507: douta=16'h83b0;
19508: douta=16'h736f;
19509: douta=16'h6b2f;
19510: douta=16'h83b0;
19511: douta=16'h7b8f;
19512: douta=16'h7b8f;
19513: douta=16'h62ee;
19514: douta=16'h6b4e;
19515: douta=16'h736f;
19516: douta=16'hc593;
19517: douta=16'hcdd4;
19518: douta=16'hbd35;
19519: douta=16'h9473;
19520: douta=16'h8c53;
19521: douta=16'h8433;
19522: douta=16'h9c94;
19523: douta=16'h8c52;
19524: douta=16'h8431;
19525: douta=16'h6b6f;
19526: douta=16'h7390;
19527: douta=16'h73b1;
19528: douta=16'h6b6f;
19529: douta=16'h632e;
19530: douta=16'h632e;
19531: douta=16'hacf3;
19532: douta=16'hd5d5;
19533: douta=16'hcdb5;
19534: douta=16'had15;
19535: douta=16'h9cf5;
19536: douta=16'h8c95;
19537: douta=16'h7c35;
19538: douta=16'h6bb2;
19539: douta=16'h6372;
19540: douta=16'h4af0;
19541: douta=16'h3a2c;
19542: douta=16'h42ae;
19543: douta=16'h29ca;
19544: douta=16'h2168;
19545: douta=16'h1948;
19546: douta=16'h29ca;
19547: douta=16'h2126;
19548: douta=16'h2147;
19549: douta=16'h10c5;
19550: douta=16'h1905;
19551: douta=16'h0000;
19552: douta=16'h7cb7;
19553: douta=16'h8cf6;
19554: douta=16'h9d79;
19555: douta=16'h9d59;
19556: douta=16'h8cf8;
19557: douta=16'h7cb7;
19558: douta=16'h5373;
19559: douta=16'h7c75;
19560: douta=16'h7cb7;
19561: douta=16'h5bb4;
19562: douta=16'h5bf5;
19563: douta=16'h8519;
19564: douta=16'h4311;
19565: douta=16'h1926;
19566: douta=16'h320b;
19567: douta=16'h29a9;
19568: douta=16'h21a9;
19569: douta=16'h2188;
19570: douta=16'h29c9;
19571: douta=16'h29c9;
19572: douta=16'h21aa;
19573: douta=16'h6aaa;
19574: douta=16'h49c7;
19575: douta=16'h49e8;
19576: douta=16'h5249;
19577: douta=16'h5229;
19578: douta=16'h5229;
19579: douta=16'h5208;
19580: douta=16'h49e8;
19581: douta=16'h5208;
19582: douta=16'h49e8;
19583: douta=16'h49e8;
19584: douta=16'he56c;
19585: douta=16'hdd4b;
19586: douta=16'hf5cc;
19587: douta=16'h28e4;
19588: douta=16'h3923;
19589: douta=16'h7b90;
19590: douta=16'h3923;
19591: douta=16'h20e4;
19592: douta=16'h0861;
19593: douta=16'h08a2;
19594: douta=16'h2105;
19595: douta=16'h10c4;
19596: douta=16'h1084;
19597: douta=16'h1948;
19598: douta=16'h320b;
19599: douta=16'h29ea;
19600: douta=16'h3a2c;
19601: douta=16'h29aa;
19602: douta=16'h320b;
19603: douta=16'h42ad;
19604: douta=16'h42ad;
19605: douta=16'h4aee;
19606: douta=16'h4b0e;
19607: douta=16'h4ace;
19608: douta=16'h4ace;
19609: douta=16'h4acd;
19610: douta=16'h3a6c;
19611: douta=16'h428c;
19612: douta=16'h4acd;
19613: douta=16'h4b0e;
19614: douta=16'h4aed;
19615: douta=16'h532e;
19616: douta=16'h4b0e;
19617: douta=16'h4acd;
19618: douta=16'h4aac;
19619: douta=16'h428b;
19620: douta=16'h52ed;
19621: douta=16'h4aac;
19622: douta=16'h4aac;
19623: douta=16'h426b;
19624: douta=16'h4acc;
19625: douta=16'h5b2e;
19626: douta=16'h5b2e;
19627: douta=16'h63f0;
19628: douta=16'h5b6f;
19629: douta=16'h63b0;
19630: douta=16'h63b0;
19631: douta=16'h63af;
19632: douta=16'h63b0;
19633: douta=16'h5b90;
19634: douta=16'h5b90;
19635: douta=16'h6b8f;
19636: douta=16'h8410;
19637: douta=16'h734e;
19638: douta=16'h422c;
19639: douta=16'hd613;
19640: douta=16'hac2b;
19641: douta=16'hf739;
19642: douta=16'hac6f;
19643: douta=16'hfef7;
19644: douta=16'hee75;
19645: douta=16'h8bf1;
19646: douta=16'hd5d3;
19647: douta=16'hbd51;
19648: douta=16'h9c93;
19649: douta=16'h8c53;
19650: douta=16'h73b0;
19651: douta=16'h736e;
19652: douta=16'h736f;
19653: douta=16'h734e;
19654: douta=16'h6b0d;
19655: douta=16'h6b2d;
19656: douta=16'h62ec;
19657: douta=16'h420a;
19658: douta=16'h832b;
19659: douta=16'hee12;
19660: douta=16'he614;
19661: douta=16'hcdd3;
19662: douta=16'hbd33;
19663: douta=16'hacf4;
19664: douta=16'hacf4;
19665: douta=16'ha515;
19666: douta=16'h9cd5;
19667: douta=16'h8474;
19668: douta=16'h8453;
19669: douta=16'h8432;
19670: douta=16'h83f1;
19671: douta=16'h5b0e;
19672: douta=16'h424c;
19673: douta=16'h4a8c;
19674: douta=16'h52ac;
19675: douta=16'h524b;
19676: douta=16'hd572;
19677: douta=16'hf674;
19678: douta=16'h73d2;
19679: douta=16'hb4f3;
19680: douta=16'had13;
19681: douta=16'h7c95;
19682: douta=16'h6b91;
19683: douta=16'h6bd2;
19684: douta=16'h7bd1;
19685: douta=16'h7b90;
19686: douta=16'h7390;
19687: douta=16'h5b2f;
19688: douta=16'h630e;
19689: douta=16'h734d;
19690: douta=16'h5aac;
19691: douta=16'h420a;
19692: douta=16'h39a8;
19693: douta=16'had15;
19694: douta=16'h9cb4;
19695: douta=16'h8454;
19696: douta=16'h7bf3;
19697: douta=16'h7bf2;
19698: douta=16'h8411;
19699: douta=16'h738f;
19700: douta=16'h7baf;
19701: douta=16'h6b2e;
19702: douta=16'h632e;
19703: douta=16'h6b4e;
19704: douta=16'h52ac;
19705: douta=16'h8bf0;
19706: douta=16'hb4f3;
19707: douta=16'hd5b4;
19708: douta=16'h73b1;
19709: douta=16'h83f1;
19710: douta=16'h9c73;
19711: douta=16'h9493;
19712: douta=16'h8452;
19713: douta=16'h83f2;
19714: douta=16'h9453;
19715: douta=16'h9453;
19716: douta=16'h8c12;
19717: douta=16'h6b4f;
19718: douta=16'h632e;
19719: douta=16'h632e;
19720: douta=16'h5aee;
19721: douta=16'h630d;
19722: douta=16'h62ed;
19723: douta=16'hac90;
19724: douta=16'hbd74;
19725: douta=16'hb534;
19726: douta=16'ha515;
19727: douta=16'h9cd5;
19728: douta=16'h8cb5;
19729: douta=16'h73f3;
19730: douta=16'h6392;
19731: douta=16'h5b71;
19732: douta=16'h4ad0;
19733: douta=16'h320c;
19734: douta=16'h4acf;
19735: douta=16'h21aa;
19736: douta=16'h29a9;
19737: douta=16'h29a9;
19738: douta=16'h6370;
19739: douta=16'h10e5;
19740: douta=16'h1927;
19741: douta=16'h1946;
19742: douta=16'h10e5;
19743: douta=16'h10e5;
19744: douta=16'h7455;
19745: douta=16'h7c96;
19746: douta=16'h6bf3;
19747: douta=16'h9518;
19748: douta=16'h84b6;
19749: douta=16'h84b7;
19750: douta=16'h7455;
19751: douta=16'h84d8;
19752: douta=16'h6c35;
19753: douta=16'h6c56;
19754: douta=16'h32b0;
19755: douta=16'h7497;
19756: douta=16'h31c9;
19757: douta=16'h2167;
19758: douta=16'h29c9;
19759: douta=16'h2188;
19760: douta=16'h29ca;
19761: douta=16'h29ea;
19762: douta=16'h320b;
19763: douta=16'h3a4c;
19764: douta=16'h3a4c;
19765: douta=16'h422a;
19766: douta=16'h5207;
19767: douta=16'h49e7;
19768: douta=16'h5208;
19769: douta=16'h5229;
19770: douta=16'h5208;
19771: douta=16'h5208;
19772: douta=16'h5229;
19773: douta=16'h5208;
19774: douta=16'h49e8;
19775: douta=16'h5208;
19776: douta=16'he56d;
19777: douta=16'hdd4c;
19778: douta=16'he54b;
19779: douta=16'h7b28;
19780: douta=16'h4985;
19781: douta=16'h51c6;
19782: douta=16'h5a6a;
19783: douta=16'h7391;
19784: douta=16'h8c13;
19785: douta=16'h73b0;
19786: douta=16'h5a6a;
19787: douta=16'h8b8e;
19788: douta=16'h9432;
19789: douta=16'had99;
19790: douta=16'h29ca;
19791: douta=16'h2169;
19792: douta=16'h322c;
19793: douta=16'h29a9;
19794: douta=16'h320b;
19795: douta=16'h3a8d;
19796: douta=16'h3a4c;
19797: douta=16'h42ae;
19798: douta=16'h3a8d;
19799: douta=16'h4b0f;
19800: douta=16'h4aee;
19801: douta=16'h428d;
19802: douta=16'h2a0a;
19803: douta=16'h324b;
19804: douta=16'h3a6b;
19805: douta=16'h3a6b;
19806: douta=16'h42ac;
19807: douta=16'h42ac;
19808: douta=16'h4acd;
19809: douta=16'h4b0e;
19810: douta=16'h42ac;
19811: douta=16'h3a6b;
19812: douta=16'h4a8c;
19813: douta=16'h428b;
19814: douta=16'h4aac;
19815: douta=16'h52ed;
19816: douta=16'h52ed;
19817: douta=16'h530d;
19818: douta=16'h5b4e;
19819: douta=16'h534e;
19820: douta=16'h532e;
19821: douta=16'h532e;
19822: douta=16'h63b0;
19823: douta=16'h5b6f;
19824: douta=16'h5b6f;
19825: douta=16'h6bd0;
19826: douta=16'h63b0;
19827: douta=16'h6390;
19828: douta=16'h7411;
19829: douta=16'h536f;
19830: douta=16'h73f0;
19831: douta=16'he675;
19832: douta=16'hd5b2;
19833: douta=16'hee96;
19834: douta=16'he675;
19835: douta=16'h93f0;
19836: douta=16'hc512;
19837: douta=16'hacd2;
19838: douta=16'h8432;
19839: douta=16'hb4f2;
19840: douta=16'h9453;
19841: douta=16'h8411;
19842: douta=16'h738f;
19843: douta=16'h62ec;
19844: douta=16'h732d;
19845: douta=16'h6b2c;
19846: douta=16'h5aaa;
19847: douta=16'h5a8b;
19848: douta=16'h836c;
19849: douta=16'hee96;
19850: douta=16'hde56;
19851: douta=16'hde15;
19852: douta=16'h7c13;
19853: douta=16'hbd54;
19854: douta=16'h9cd4;
19855: douta=16'h9495;
19856: douta=16'h94d5;
19857: douta=16'h94b5;
19858: douta=16'h7bf2;
19859: douta=16'h7bf1;
19860: douta=16'h7bb0;
19861: douta=16'h6b0d;
19862: douta=16'h6b2d;
19863: douta=16'h734f;
19864: douta=16'h528c;
19865: douta=16'h4a4c;
19866: douta=16'hb46f;
19867: douta=16'hcd51;
19868: douta=16'ha494;
19869: douta=16'ha4b4;
19870: douta=16'h8453;
19871: douta=16'h6bb1;
19872: douta=16'h9c93;
19873: douta=16'h7390;
19874: douta=16'h62ee;
19875: douta=16'h632f;
19876: douta=16'h4aad;
19877: douta=16'h6b2e;
19878: douta=16'h7b4e;
19879: douta=16'h5a6b;
19880: douta=16'h526b;
19881: douta=16'h5a8b;
19882: douta=16'h9c94;
19883: douta=16'h73d0;
19884: douta=16'h7b6f;
19885: douta=16'h734d;
19886: douta=16'h734d;
19887: douta=16'h732d;
19888: douta=16'h4a8b;
19889: douta=16'h52ac;
19890: douta=16'h5aed;
19891: douta=16'h7baf;
19892: douta=16'h732e;
19893: douta=16'h4a6c;
19894: douta=16'hbd32;
19895: douta=16'hee35;
19896: douta=16'h9493;
19897: douta=16'h8c32;
19898: douta=16'ha4d4;
19899: douta=16'h9c94;
19900: douta=16'h6b6f;
19901: douta=16'h6b4f;
19902: douta=16'h7bd1;
19903: douta=16'h5aee;
19904: douta=16'h52cd;
19905: douta=16'h632e;
19906: douta=16'h7bb0;
19907: douta=16'h734e;
19908: douta=16'h632e;
19909: douta=16'h7b8f;
19910: douta=16'h8c10;
19911: douta=16'h8bef;
19912: douta=16'hd616;
19913: douta=16'he678;
19914: douta=16'hde36;
19915: douta=16'hcdb5;
19916: douta=16'hbd74;
19917: douta=16'h94d5;
19918: douta=16'h8454;
19919: douta=16'h8454;
19920: douta=16'h73d1;
19921: douta=16'h6b91;
19922: douta=16'h6371;
19923: douta=16'h6371;
19924: douta=16'h5330;
19925: douta=16'h4acf;
19926: douta=16'h3a4d;
19927: douta=16'h3a6e;
19928: douta=16'h21aa;
19929: douta=16'h52ed;
19930: douta=16'h2148;
19931: douta=16'h428c;
19932: douta=16'h10e4;
19933: douta=16'h10c5;
19934: douta=16'h10c4;
19935: douta=16'h18e5;
19936: douta=16'h1927;
19937: douta=16'h7413;
19938: douta=16'h9d79;
19939: douta=16'h6bd4;
19940: douta=16'h7414;
19941: douta=16'h7434;
19942: douta=16'h63f5;
19943: douta=16'h8d18;
19944: douta=16'h8cf8;
19945: douta=16'ha5db;
19946: douta=16'h4b10;
19947: douta=16'h2126;
19948: douta=16'h3a2b;
19949: douta=16'h3a2b;
19950: douta=16'h424b;
19951: douta=16'h426c;
19952: douta=16'h5bb2;
19953: douta=16'h63d3;
19954: douta=16'h5bf4;
19955: douta=16'h6435;
19956: douta=16'h5bb3;
19957: douta=16'h5c36;
19958: douta=16'h42cf;
19959: douta=16'h5b92;
19960: douta=16'h49c6;
19961: douta=16'h3986;
19962: douta=16'h49c7;
19963: douta=16'h41c7;
19964: douta=16'h49e7;
19965: douta=16'h49e7;
19966: douta=16'h49e8;
19967: douta=16'h49c7;
19968: douta=16'he58d;
19969: douta=16'he56c;
19970: douta=16'hdd4b;
19971: douta=16'hc509;
19972: douta=16'h51c5;
19973: douta=16'h5164;
19974: douta=16'h83ad;
19975: douta=16'hbd98;
19976: douta=16'h83f2;
19977: douta=16'h7bf1;
19978: douta=16'h8b4d;
19979: douta=16'ha410;
19980: douta=16'had57;
19981: douta=16'h9d17;
19982: douta=16'h21ca;
19983: douta=16'h29eb;
19984: douta=16'h320c;
19985: douta=16'h2189;
19986: douta=16'h320b;
19987: douta=16'h42ae;
19988: douta=16'h3a6d;
19989: douta=16'h3a8d;
19990: douta=16'h3a6d;
19991: douta=16'h42ae;
19992: douta=16'h428d;
19993: douta=16'h42ad;
19994: douta=16'h324b;
19995: douta=16'h322a;
19996: douta=16'h3a4b;
19997: douta=16'h3a6b;
19998: douta=16'h3a8c;
19999: douta=16'h428c;
20000: douta=16'h3a6b;
20001: douta=16'h3a8c;
20002: douta=16'h4b0e;
20003: douta=16'h4b0e;
20004: douta=16'h3a6b;
20005: douta=16'h322a;
20006: douta=16'h4a8c;
20007: douta=16'h4aac;
20008: douta=16'h530d;
20009: douta=16'h530e;
20010: douta=16'h5b4e;
20011: douta=16'h5b6f;
20012: douta=16'h5b6f;
20013: douta=16'h534e;
20014: douta=16'h532e;
20015: douta=16'h5b6f;
20016: douta=16'h5b4f;
20017: douta=16'h6390;
20018: douta=16'h6390;
20019: douta=16'h63b0;
20020: douta=16'h6c11;
20021: douta=16'h5b70;
20022: douta=16'h63af;
20023: douta=16'hcd71;
20024: douta=16'hc510;
20025: douta=16'hd5b4;
20026: douta=16'hbd33;
20027: douta=16'hacb2;
20028: douta=16'h9c93;
20029: douta=16'hacd2;
20030: douta=16'h8432;
20031: douta=16'h9c93;
20032: douta=16'h7bf1;
20033: douta=16'h83d0;
20034: douta=16'h7baf;
20035: douta=16'h6b2e;
20036: douta=16'h6b0d;
20037: douta=16'h6b0c;
20038: douta=16'h62ed;
20039: douta=16'h8b29;
20040: douta=16'hd5f3;
20041: douta=16'he655;
20042: douta=16'hde35;
20043: douta=16'hbd75;
20044: douta=16'h84b5;
20045: douta=16'h8c74;
20046: douta=16'hb556;
20047: douta=16'h8454;
20048: douta=16'h8c94;
20049: douta=16'h8c94;
20050: douta=16'h7370;
20051: douta=16'h734e;
20052: douta=16'h734e;
20053: douta=16'h7b6f;
20054: douta=16'h8390;
20055: douta=16'h52ac;
20056: douta=16'hddb2;
20057: douta=16'hd5b3;
20058: douta=16'hd593;
20059: douta=16'hb533;
20060: douta=16'hbd55;
20061: douta=16'ha4b4;
20062: douta=16'h9495;
20063: douta=16'h8434;
20064: douta=16'h6371;
20065: douta=16'h7bb1;
20066: douta=16'h736f;
20067: douta=16'h62cd;
20068: douta=16'h31ca;
20069: douta=16'h420a;
20070: douta=16'h31a8;
20071: douta=16'h526c;
20072: douta=16'h7bb0;
20073: douta=16'ha4b5;
20074: douta=16'h7370;
20075: douta=16'h732e;
20076: douta=16'h62ed;
20077: douta=16'h732d;
20078: douta=16'h732d;
20079: douta=16'h734d;
20080: douta=16'h422a;
20081: douta=16'h31c9;
20082: douta=16'h31a8;
20083: douta=16'h420c;
20084: douta=16'hcdb4;
20085: douta=16'hd595;
20086: douta=16'ha4b4;
20087: douta=16'h9cb5;
20088: douta=16'h9474;
20089: douta=16'h8c74;
20090: douta=16'h7bd1;
20091: douta=16'h7b8f;
20092: douta=16'h734e;
20093: douta=16'h6b0e;
20094: douta=16'h5acc;
20095: douta=16'h630d;
20096: douta=16'h5aed;
20097: douta=16'h422b;
20098: douta=16'h3a2b;
20099: douta=16'h62ac;
20100: douta=16'h836d;
20101: douta=16'heeb7;
20102: douta=16'he697;
20103: douta=16'hde57;
20104: douta=16'hcdf6;
20105: douta=16'hc5b6;
20106: douta=16'hbd76;
20107: douta=16'had15;
20108: douta=16'had15;
20109: douta=16'h9c94;
20110: douta=16'h7bd1;
20111: douta=16'h6b91;
20112: douta=16'h6b91;
20113: douta=16'h6b90;
20114: douta=16'h6b91;
20115: douta=16'h6b91;
20116: douta=16'h52ef;
20117: douta=16'h4ace;
20118: douta=16'h4aae;
20119: douta=16'h62eb;
20120: douta=16'hc574;
20121: douta=16'h6b92;
20122: douta=16'h2168;
20123: douta=16'h18c5;
20124: douta=16'h5b50;
20125: douta=16'h10a4;
20126: douta=16'h10c4;
20127: douta=16'h18e5;
20128: douta=16'h10e5;
20129: douta=16'h0083;
20130: douta=16'h63b2;
20131: douta=16'h8cd7;
20132: douta=16'h9d58;
20133: douta=16'h6c15;
20134: douta=16'h6c16;
20135: douta=16'h9d58;
20136: douta=16'ha599;
20137: douta=16'h4b10;
20138: douta=16'h5330;
20139: douta=16'h63f2;
20140: douta=16'h6c34;
20141: douta=16'h6c14;
20142: douta=16'h7cf7;
20143: douta=16'h855a;
20144: douta=16'h6bf3;
20145: douta=16'h5b50;
20146: douta=16'h5a47;
20147: douta=16'h6247;
20148: douta=16'h6a25;
20149: douta=16'h69e4;
20150: douta=16'h61e4;
20151: douta=16'h61e4;
20152: douta=16'h6a47;
20153: douta=16'h5a28;
20154: douta=16'h41a7;
20155: douta=16'h49e7;
20156: douta=16'h41a7;
20157: douta=16'h49c7;
20158: douta=16'h49c7;
20159: douta=16'h41c7;
20160: douta=16'he58d;
20161: douta=16'he56d;
20162: douta=16'he56c;
20163: douta=16'he58c;
20164: douta=16'h59e6;
20165: douta=16'h51c5;
20166: douta=16'h8bae;
20167: douta=16'hb516;
20168: douta=16'h8c32;
20169: douta=16'h9452;
20170: douta=16'ha40f;
20171: douta=16'hac51;
20172: douta=16'hb557;
20173: douta=16'h9d17;
20174: douta=16'h2188;
20175: douta=16'h29ca;
20176: douta=16'h322c;
20177: douta=16'h2188;
20178: douta=16'h29aa;
20179: douta=16'h322c;
20180: douta=16'h3a4c;
20181: douta=16'h42ae;
20182: douta=16'h3a6d;
20183: douta=16'h3a8d;
20184: douta=16'h3a8d;
20185: douta=16'h428d;
20186: douta=16'h322a;
20187: douta=16'h322b;
20188: douta=16'h322a;
20189: douta=16'h324b;
20190: douta=16'h3a6b;
20191: douta=16'h3a6c;
20192: douta=16'h3a6c;
20193: douta=16'h428c;
20194: douta=16'h4b0e;
20195: douta=16'h4b2e;
20196: douta=16'h530e;
20197: douta=16'h3a2a;
20198: douta=16'h322a;
20199: douta=16'h3a4a;
20200: douta=16'h530d;
20201: douta=16'h4acd;
20202: douta=16'h5b6f;
20203: douta=16'h63b0;
20204: douta=16'h534e;
20205: douta=16'h4b0d;
20206: douta=16'h5b4f;
20207: douta=16'h5b4f;
20208: douta=16'h5b6f;
20209: douta=16'h6390;
20210: douta=16'h6390;
20211: douta=16'h6390;
20212: douta=16'h63b1;
20213: douta=16'h6390;
20214: douta=16'h638f;
20215: douta=16'h6b6f;
20216: douta=16'h7bce;
20217: douta=16'hbcf1;
20218: douta=16'hb4f2;
20219: douta=16'h9c51;
20220: douta=16'ha472;
20221: douta=16'hacd3;
20222: douta=16'h8433;
20223: douta=16'h8412;
20224: douta=16'h83f0;
20225: douta=16'h7bd0;
20226: douta=16'h7baf;
20227: douta=16'h7b6f;
20228: douta=16'h6b0c;
20229: douta=16'h6b0d;
20230: douta=16'h8bad;
20231: douta=16'hd591;
20232: douta=16'hd5d4;
20233: douta=16'hde15;
20234: douta=16'hcdb4;
20235: douta=16'had15;
20236: douta=16'h94d6;
20237: douta=16'h6371;
20238: douta=16'h9494;
20239: douta=16'h73d1;
20240: douta=16'h73d0;
20241: douta=16'h8453;
20242: douta=16'h7bb0;
20243: douta=16'h736e;
20244: douta=16'h736e;
20245: douta=16'h736e;
20246: douta=16'h62ed;
20247: douta=16'h8bce;
20248: douta=16'hee55;
20249: douta=16'hcdb4;
20250: douta=16'hacf3;
20251: douta=16'h6bb2;
20252: douta=16'h8413;
20253: douta=16'h8c53;
20254: douta=16'h8433;
20255: douta=16'h7bf3;
20256: douta=16'h6b91;
20257: douta=16'h6b6f;
20258: douta=16'h7391;
20259: douta=16'h7391;
20260: douta=16'h5a8b;
20261: douta=16'h4a2a;
20262: douta=16'h5a8b;
20263: douta=16'h6b71;
20264: douta=16'h6370;
20265: douta=16'h9432;
20266: douta=16'h7b90;
20267: douta=16'h6aec;
20268: douta=16'h62cc;
20269: douta=16'h526b;
20270: douta=16'h5a8b;
20271: douta=16'h732c;
20272: douta=16'h6acb;
20273: douta=16'h31c9;
20274: douta=16'h422a;
20275: douta=16'h8413;
20276: douta=16'hacd3;
20277: douta=16'hacf5;
20278: douta=16'h9cb5;
20279: douta=16'ha4d5;
20280: douta=16'h8c73;
20281: douta=16'h8433;
20282: douta=16'h8432;
20283: douta=16'h7bf2;
20284: douta=16'h6b0d;
20285: douta=16'h6aed;
20286: douta=16'h62cd;
20287: douta=16'h5acd;
20288: douta=16'h5aee;
20289: douta=16'h4a6c;
20290: douta=16'h838e;
20291: douta=16'h93ee;
20292: douta=16'hac6f;
20293: douta=16'hde36;
20294: douta=16'hd617;
20295: douta=16'hbd96;
20296: douta=16'hb536;
20297: douta=16'hb556;
20298: douta=16'hbd76;
20299: douta=16'had15;
20300: douta=16'h9494;
20301: douta=16'h8432;
20302: douta=16'h6b90;
20303: douta=16'h6b90;
20304: douta=16'h6b90;
20305: douta=16'h73f2;
20306: douta=16'h6b91;
20307: douta=16'h6350;
20308: douta=16'h52ce;
20309: douta=16'h52cf;
20310: douta=16'h31c9;
20311: douta=16'he634;
20312: douta=16'h8c52;
20313: douta=16'h4acf;
20314: douta=16'h39ea;
20315: douta=16'h1906;
20316: douta=16'h2987;
20317: douta=16'h0863;
20318: douta=16'h18c4;
20319: douta=16'h18e4;
20320: douta=16'h10e4;
20321: douta=16'h1947;
20322: douta=16'h42ce;
20323: douta=16'h84b6;
20324: douta=16'h7c96;
20325: douta=16'h84d7;
20326: douta=16'h84b7;
20327: douta=16'h9518;
20328: douta=16'h84b8;
20329: douta=16'h42ee;
20330: douta=16'h7cf8;
20331: douta=16'h7d19;
20332: douta=16'h7413;
20333: douta=16'h6390;
20334: douta=16'h73d0;
20335: douta=16'h6a47;
20336: douta=16'h6a25;
20337: douta=16'h7246;
20338: douta=16'h7224;
20339: douta=16'h6a25;
20340: douta=16'h6a25;
20341: douta=16'h6a26;
20342: douta=16'h6205;
20343: douta=16'h6205;
20344: douta=16'h59e5;
20345: douta=16'h728a;
20346: douta=16'h41c7;
20347: douta=16'h49e7;
20348: douta=16'h49e7;
20349: douta=16'h49e8;
20350: douta=16'h49e8;
20351: douta=16'h49e7;
20352: douta=16'hedae;
20353: douta=16'he56d;
20354: douta=16'he56c;
20355: douta=16'hedac;
20356: douta=16'h6226;
20357: douta=16'h7267;
20358: douta=16'h4964;
20359: douta=16'hbd13;
20360: douta=16'h9c72;
20361: douta=16'h9432;
20362: douta=16'hdd93;
20363: douta=16'hd5d5;
20364: douta=16'hbd97;
20365: douta=16'h73f3;
20366: douta=16'h6393;
20367: douta=16'h6c14;
20368: douta=16'h1927;
20369: douta=16'h2188;
20370: douta=16'h21a9;
20371: douta=16'h322c;
20372: douta=16'h2a0b;
20373: douta=16'h322c;
20374: douta=16'h3a4d;
20375: douta=16'h320b;
20376: douta=16'h320b;
20377: douta=16'h320b;
20378: douta=16'h29ca;
20379: douta=16'h3a4c;
20380: douta=16'h3a4c;
20381: douta=16'h322b;
20382: douta=16'h3a4c;
20383: douta=16'h3a8c;
20384: douta=16'h3a6b;
20385: douta=16'h3a6b;
20386: douta=16'h3a8c;
20387: douta=16'h42ad;
20388: douta=16'h42ac;
20389: douta=16'h530e;
20390: douta=16'h5b2e;
20391: douta=16'h5b2e;
20392: douta=16'h5b4f;
20393: douta=16'h5b2f;
20394: douta=16'h530e;
20395: douta=16'h532e;
20396: douta=16'h4aad;
20397: douta=16'h4aed;
20398: douta=16'h532e;
20399: douta=16'h530e;
20400: douta=16'h534f;
20401: douta=16'h63b0;
20402: douta=16'h5b6f;
20403: douta=16'h6390;
20404: douta=16'h6390;
20405: douta=16'h638f;
20406: douta=16'h6390;
20407: douta=16'h638f;
20408: douta=16'h638f;
20409: douta=16'h6bd0;
20410: douta=16'h73d0;
20411: douta=16'h8c0f;
20412: douta=16'h93ef;
20413: douta=16'h8bcf;
20414: douta=16'h83cf;
20415: douta=16'h7b8e;
20416: douta=16'h7bcf;
20417: douta=16'h7baf;
20418: douta=16'h6b2c;
20419: douta=16'h528b;
20420: douta=16'h7b0c;
20421: douta=16'hcd10;
20422: douta=16'hcdd4;
20423: douta=16'heeb7;
20424: douta=16'hbd74;
20425: douta=16'ha536;
20426: douta=16'ha537;
20427: douta=16'ha516;
20428: douta=16'h8c95;
20429: douta=16'h8c95;
20430: douta=16'h8413;
20431: douta=16'h9493;
20432: douta=16'h7bf1;
20433: douta=16'h6b6f;
20434: douta=16'h6b4f;
20435: douta=16'h630e;
20436: douta=16'h62ed;
20437: douta=16'ha3ee;
20438: douta=16'hee55;
20439: douta=16'hb4d1;
20440: douta=16'hacd3;
20441: douta=16'ha4f4;
20442: douta=16'h9cd5;
20443: douta=16'h9cf6;
20444: douta=16'h7413;
20445: douta=16'h634f;
20446: douta=16'h3a0a;
20447: douta=16'h52ac;
20448: douta=16'h7b4e;
20449: douta=16'h7b4d;
20450: douta=16'h62cb;
20451: douta=16'h4a09;
20452: douta=16'h8c32;
20453: douta=16'h5ace;
20454: douta=16'h9412;
20455: douta=16'h62ed;
20456: douta=16'h6b0e;
20457: douta=16'h5a8c;
20458: douta=16'h4a2b;
20459: douta=16'h6b0c;
20460: douta=16'h6aeb;
20461: douta=16'h41a8;
20462: douta=16'h3167;
20463: douta=16'h41e8;
20464: douta=16'hb556;
20465: douta=16'h8c74;
20466: douta=16'h9c94;
20467: douta=16'h8454;
20468: douta=16'h73d2;
20469: douta=16'h9c92;
20470: douta=16'h8432;
20471: douta=16'h8c52;
20472: douta=16'h73b0;
20473: douta=16'h7bd1;
20474: douta=16'h7bb0;
20475: douta=16'h736f;
20476: douta=16'h528c;
20477: douta=16'h528c;
20478: douta=16'h7b6d;
20479: douta=16'hee75;
20480: douta=16'hee96;
20481: douta=16'hcdb5;
20482: douta=16'hb535;
20483: douta=16'hbd75;
20484: douta=16'hc575;
20485: douta=16'ha4b2;
20486: douta=16'had14;
20487: douta=16'had15;
20488: douta=16'ha4f5;
20489: douta=16'h9473;
20490: douta=16'h8c73;
20491: douta=16'h8c53;
20492: douta=16'h8433;
20493: douta=16'h8432;
20494: douta=16'h8432;
20495: douta=16'h7c12;
20496: douta=16'h6b70;
20497: douta=16'h6b50;
20498: douta=16'h6350;
20499: douta=16'h52ad;
20500: douta=16'hac8e;
20501: douta=16'hcd92;
20502: douta=16'hde14;
20503: douta=16'hcd73;
20504: douta=16'h6371;
20505: douta=16'h324d;
20506: douta=16'h6350;
20507: douta=16'h322c;
20508: douta=16'h324c;
20509: douta=16'h18e5;
20510: douta=16'h3a4c;
20511: douta=16'h1083;
20512: douta=16'h2168;
20513: douta=16'h10e5;
20514: douta=16'h10e5;
20515: douta=16'h6c36;
20516: douta=16'h6c14;
20517: douta=16'h63b3;
20518: douta=16'h9558;
20519: douta=16'h20a2;
20520: douta=16'h1860;
20521: douta=16'h61c3;
20522: douta=16'h7a44;
20523: douta=16'h7a65;
20524: douta=16'h7245;
20525: douta=16'h7245;
20526: douta=16'h7245;
20527: douta=16'h6a04;
20528: douta=16'h6a24;
20529: douta=16'h6a25;
20530: douta=16'h6a25;
20531: douta=16'h6205;
20532: douta=16'h6a05;
20533: douta=16'h61e5;
20534: douta=16'h61e5;
20535: douta=16'h59e5;
20536: douta=16'h59c5;
20537: douta=16'h4964;
20538: douta=16'h8bf0;
20539: douta=16'h49e7;
20540: douta=16'h4a08;
20541: douta=16'h5209;
20542: douta=16'h41a7;
20543: douta=16'h41c7;
20544: douta=16'he5ae;
20545: douta=16'he56c;
20546: douta=16'he56c;
20547: douta=16'he56b;
20548: douta=16'h6205;
20549: douta=16'h7aa8;
20550: douta=16'h8aeb;
20551: douta=16'hb4b2;
20552: douta=16'hac92;
20553: douta=16'hac71;
20554: douta=16'hee77;
20555: douta=16'he676;
20556: douta=16'hb515;
20557: douta=16'h6bb3;
20558: douta=16'h7c55;
20559: douta=16'h7c76;
20560: douta=16'h322b;
20561: douta=16'h1927;
20562: douta=16'h31ea;
20563: douta=16'h322c;
20564: douta=16'h326d;
20565: douta=16'h326d;
20566: douta=16'h3a8d;
20567: douta=16'h3a8d;
20568: douta=16'h322c;
20569: douta=16'h3a6d;
20570: douta=16'h3a4c;
20571: douta=16'h29ca;
20572: douta=16'h2a0a;
20573: douta=16'h3a6c;
20574: douta=16'h3a4c;
20575: douta=16'h42ad;
20576: douta=16'h3a8c;
20577: douta=16'h3a8d;
20578: douta=16'h324b;
20579: douta=16'h3a6b;
20580: douta=16'h42cd;
20581: douta=16'h5b0e;
20582: douta=16'h636f;
20583: douta=16'h5b4e;
20584: douta=16'h6370;
20585: douta=16'h634f;
20586: douta=16'h534f;
20587: douta=16'h4b0e;
20588: douta=16'h532e;
20589: douta=16'h530e;
20590: douta=16'h532f;
20591: douta=16'h534f;
20592: douta=16'h532e;
20593: douta=16'h534f;
20594: douta=16'h5b4f;
20595: douta=16'h5b2f;
20596: douta=16'h5b6f;
20597: douta=16'h5b6f;
20598: douta=16'h5b4f;
20599: douta=16'h5b6f;
20600: douta=16'h638f;
20601: douta=16'h638f;
20602: douta=16'h6b90;
20603: douta=16'h6bd0;
20604: douta=16'h638f;
20605: douta=16'h6baf;
20606: douta=16'h736e;
20607: douta=16'h734c;
20608: douta=16'h732c;
20609: douta=16'h72cb;
20610: douta=16'h5a8a;
20611: douta=16'hddb3;
20612: douta=16'hde55;
20613: douta=16'heeb7;
20614: douta=16'he656;
20615: douta=16'hc574;
20616: douta=16'hb555;
20617: douta=16'had36;
20618: douta=16'h9d17;
20619: douta=16'h94b6;
20620: douta=16'h8c75;
20621: douta=16'h7bf2;
20622: douta=16'h7bd1;
20623: douta=16'h6b4f;
20624: douta=16'h7bf1;
20625: douta=16'h73b1;
20626: douta=16'h734f;
20627: douta=16'h4a6c;
20628: douta=16'h730d;
20629: douta=16'hddf4;
20630: douta=16'hd593;
20631: douta=16'h8c54;
20632: douta=16'h94b5;
20633: douta=16'h9cd5;
20634: douta=16'h8c95;
20635: douta=16'h7c12;
20636: douta=16'h6b90;
20637: douta=16'h6b6f;
20638: douta=16'h528c;
20639: douta=16'h3a2b;
20640: douta=16'h29ca;
20641: douta=16'h29aa;
20642: douta=16'h93f0;
20643: douta=16'hb4d4;
20644: douta=16'h73f2;
20645: douta=16'h424c;
20646: douta=16'h4a4c;
20647: douta=16'h734e;
20648: douta=16'h6b0c;
20649: douta=16'h6b0c;
20650: douta=16'h5aab;
20651: douta=16'h522a;
20652: douta=16'h39e9;
20653: douta=16'h732c;
20654: douta=16'hc511;
20655: douta=16'hd593;
20656: douta=16'ha4f6;
20657: douta=16'h73d2;
20658: douta=16'h6b91;
20659: douta=16'h8453;
20660: douta=16'h7bf2;
20661: douta=16'h73b1;
20662: douta=16'h5b0f;
20663: douta=16'h3a6d;
20664: douta=16'h52ce;
20665: douta=16'h734f;
20666: douta=16'h6b4e;
20667: douta=16'h630d;
20668: douta=16'hc552;
20669: douta=16'hd5d4;
20670: douta=16'hde77;
20671: douta=16'he676;
20672: douta=16'hde15;
20673: douta=16'hc595;
20674: douta=16'hb536;
20675: douta=16'h8c51;
20676: douta=16'h8c51;
20677: douta=16'h8c31;
20678: douta=16'h9c93;
20679: douta=16'had35;
20680: douta=16'h9cf5;
20681: douta=16'h9474;
20682: douta=16'h8c73;
20683: douta=16'h8c53;
20684: douta=16'h83f2;
20685: douta=16'h7390;
20686: douta=16'h73b0;
20687: douta=16'h6b90;
20688: douta=16'h6b90;
20689: douta=16'h528b;
20690: douta=16'h6aeb;
20691: douta=16'h8bee;
20692: douta=16'hcdb4;
20693: douta=16'hde34;
20694: douta=16'hddd4;
20695: douta=16'had14;
20696: douta=16'h7c13;
20697: douta=16'h530f;
20698: douta=16'h5b50;
20699: douta=16'h4aef;
20700: douta=16'h42cf;
20701: douta=16'h322d;
20702: douta=16'h29ca;
20703: douta=16'h3a4d;
20704: douta=16'h29a8;
20705: douta=16'h2988;
20706: douta=16'h2147;
20707: douta=16'h5371;
20708: douta=16'h9d59;
20709: douta=16'ha5da;
20710: douta=16'h1020;
20711: douta=16'h2904;
20712: douta=16'h59a4;
20713: douta=16'h7a44;
20714: douta=16'h7a44;
20715: douta=16'h7a65;
20716: douta=16'h7244;
20717: douta=16'h7245;
20718: douta=16'h7224;
20719: douta=16'h6a24;
20720: douta=16'h6a24;
20721: douta=16'h6a04;
20722: douta=16'h6205;
20723: douta=16'h6205;
20724: douta=16'h6205;
20725: douta=16'h59e5;
20726: douta=16'h61e5;
20727: douta=16'h59e5;
20728: douta=16'h59c5;
20729: douta=16'h51c6;
20730: douta=16'h4964;
20731: douta=16'h7b4e;
20732: douta=16'h5208;
20733: douta=16'h41a7;
20734: douta=16'h49e8;
20735: douta=16'h41c8;
20736: douta=16'hedae;
20737: douta=16'he58d;
20738: douta=16'he56c;
20739: douta=16'hdd6c;
20740: douta=16'h6a26;
20741: douta=16'h8ae8;
20742: douta=16'h9bae;
20743: douta=16'hb492;
20744: douta=16'hac91;
20745: douta=16'hb4b1;
20746: douta=16'hee56;
20747: douta=16'hee97;
20748: douta=16'hb514;
20749: douta=16'h63b2;
20750: douta=16'h7c76;
20751: douta=16'h84b7;
20752: douta=16'h1106;
20753: douta=16'h2168;
20754: douta=16'h2188;
20755: douta=16'h2a2b;
20756: douta=16'h322d;
20757: douta=16'h324d;
20758: douta=16'h3a8e;
20759: douta=16'h3a8e;
20760: douta=16'h3a8d;
20761: douta=16'h3a8d;
20762: douta=16'h324c;
20763: douta=16'h29ca;
20764: douta=16'h320b;
20765: douta=16'h320b;
20766: douta=16'h3a4c;
20767: douta=16'h42ad;
20768: douta=16'h428d;
20769: douta=16'h428d;
20770: douta=16'h42ad;
20771: douta=16'h4ace;
20772: douta=16'h42ad;
20773: douta=16'h4aad;
20774: douta=16'h4aac;
20775: douta=16'h4aac;
20776: douta=16'h4acd;
20777: douta=16'h4aed;
20778: douta=16'h534f;
20779: douta=16'h536f;
20780: douta=16'h534f;
20781: douta=16'h532f;
20782: douta=16'h532e;
20783: douta=16'h532e;
20784: douta=16'h5b4f;
20785: douta=16'h532f;
20786: douta=16'h5b4f;
20787: douta=16'h534f;
20788: douta=16'h5b4f;
20789: douta=16'h5b6e;
20790: douta=16'h5b6f;
20791: douta=16'h636f;
20792: douta=16'h638f;
20793: douta=16'h636f;
20794: douta=16'h634f;
20795: douta=16'h638f;
20796: douta=16'h638f;
20797: douta=16'h638f;
20798: douta=16'h6bd0;
20799: douta=16'h6b6e;
20800: douta=16'h7bae;
20801: douta=16'h738e;
20802: douta=16'h8bce;
20803: douta=16'heed7;
20804: douta=16'he676;
20805: douta=16'he6b7;
20806: douta=16'hc5b6;
20807: douta=16'hbd75;
20808: douta=16'hb556;
20809: douta=16'hb596;
20810: douta=16'h94f6;
20811: douta=16'h8c54;
20812: douta=16'h8433;
20813: douta=16'h6b6f;
20814: douta=16'h6b6f;
20815: douta=16'h734f;
20816: douta=16'h7b90;
20817: douta=16'h8412;
20818: douta=16'h632f;
20819: douta=16'h8b4c;
20820: douta=16'hdd92;
20821: douta=16'hddf3;
20822: douta=16'hc553;
20823: douta=16'h8c74;
20824: douta=16'h8c74;
20825: douta=16'h8c74;
20826: douta=16'h8454;
20827: douta=16'h7c12;
20828: douta=16'h73b0;
20829: douta=16'h6b6f;
20830: douta=16'h62cb;
20831: douta=16'h62ab;
20832: douta=16'h62ab;
20833: douta=16'h7b2c;
20834: douta=16'hb4f4;
20835: douta=16'h8c53;
20836: douta=16'h73b1;
20837: douta=16'h52ad;
20838: douta=16'h31eb;
20839: douta=16'h732d;
20840: douta=16'h7b6d;
20841: douta=16'h6aec;
20842: douta=16'h6aab;
20843: douta=16'h72ec;
20844: douta=16'h5a6a;
20845: douta=16'he5f4;
20846: douta=16'he5d4;
20847: douta=16'hbd54;
20848: douta=16'h9cd5;
20849: douta=16'h8454;
20850: douta=16'h6b72;
20851: douta=16'h8c32;
20852: douta=16'h7bf1;
20853: douta=16'h632f;
20854: douta=16'h83f2;
20855: douta=16'h6b4f;
20856: douta=16'h31ec;
20857: douta=16'h426d;
20858: douta=16'h4a8c;
20859: douta=16'h6b2d;
20860: douta=16'hde35;
20861: douta=16'hbd33;
20862: douta=16'hde35;
20863: douta=16'hc5b5;
20864: douta=16'hc595;
20865: douta=16'hbd76;
20866: douta=16'had36;
20867: douta=16'ha515;
20868: douta=16'h9cd4;
20869: douta=16'h9452;
20870: douta=16'h8c31;
20871: douta=16'h9cb3;
20872: douta=16'h9cd4;
20873: douta=16'h9494;
20874: douta=16'h8c73;
20875: douta=16'h7bd1;
20876: douta=16'h7bf2;
20877: douta=16'h7bd1;
20878: douta=16'h73d1;
20879: douta=16'h7bb1;
20880: douta=16'h5acc;
20881: douta=16'h6aeb;
20882: douta=16'hc531;
20883: douta=16'hd5d3;
20884: douta=16'he676;
20885: douta=16'hd5f4;
20886: douta=16'hc554;
20887: douta=16'h9cd5;
20888: douta=16'h8c95;
20889: douta=16'h7c54;
20890: douta=16'h5b50;
20891: douta=16'h5351;
20892: douta=16'h4b10;
20893: douta=16'h3a6e;
20894: douta=16'h324d;
20895: douta=16'h21a9;
20896: douta=16'h31a9;
20897: douta=16'h2167;
20898: douta=16'h1927;
20899: douta=16'h08a4;
20900: douta=16'h08a4;
20901: douta=16'h8cf7;
20902: douta=16'h1021;
20903: douta=16'h51a4;
20904: douta=16'h7a63;
20905: douta=16'h7a65;
20906: douta=16'h7a65;
20907: douta=16'h7a44;
20908: douta=16'h7244;
20909: douta=16'h7224;
20910: douta=16'h7224;
20911: douta=16'h6a04;
20912: douta=16'h6204;
20913: douta=16'h6205;
20914: douta=16'h61e4;
20915: douta=16'h6205;
20916: douta=16'h61e5;
20917: douta=16'h61e5;
20918: douta=16'h59e5;
20919: douta=16'h59c5;
20920: douta=16'h59c5;
20921: douta=16'h51c5;
20922: douta=16'h51a5;
20923: douta=16'h49a5;
20924: douta=16'h4986;
20925: douta=16'h49e8;
20926: douta=16'h3965;
20927: douta=16'h3966;
20928: douta=16'he5ad;
20929: douta=16'he58c;
20930: douta=16'he54c;
20931: douta=16'he54c;
20932: douta=16'ha3e8;
20933: douta=16'h7204;
20934: douta=16'hf698;
20935: douta=16'hcd12;
20936: douta=16'hc4f1;
20937: douta=16'hc4af;
20938: douta=16'hf718;
20939: douta=16'heed9;
20940: douta=16'hacf5;
20941: douta=16'h8496;
20942: douta=16'h8496;
20943: douta=16'h8d19;
20944: douta=16'h6370;
20945: douta=16'h6bd3;
20946: douta=16'h428e;
20947: douta=16'h2a0b;
20948: douta=16'h2a0b;
20949: douta=16'h2a0c;
20950: douta=16'h326d;
20951: douta=16'h3a8e;
20952: douta=16'h3a8d;
20953: douta=16'h3a8d;
20954: douta=16'h3aad;
20955: douta=16'h2189;
20956: douta=16'h2a0b;
20957: douta=16'h31eb;
20958: douta=16'h320b;
20959: douta=16'h322b;
20960: douta=16'h322b;
20961: douta=16'h29a7;
20962: douta=16'h18c4;
20963: douta=16'h18e4;
20964: douta=16'h2125;
20965: douta=16'h2966;
20966: douta=16'h3187;
20967: douta=16'h2967;
20968: douta=16'h2986;
20969: douta=16'h2966;
20970: douta=16'h2967;
20971: douta=16'h2126;
20972: douta=16'h1905;
20973: douta=16'h18e5;
20974: douta=16'h2147;
20975: douta=16'h3a6b;
20976: douta=16'h4b0e;
20977: douta=16'h4aee;
20978: douta=16'h4aee;
20979: douta=16'h5b6f;
20980: douta=16'h532e;
20981: douta=16'h5b4e;
20982: douta=16'h5b4f;
20983: douta=16'h5b4e;
20984: douta=16'h530e;
20985: douta=16'h5b2e;
20986: douta=16'h638f;
20987: douta=16'h636e;
20988: douta=16'h636f;
20989: douta=16'h638f;
20990: douta=16'h6bb0;
20991: douta=16'h6b90;
20992: douta=16'h6bb0;
20993: douta=16'h6bd0;
20994: douta=16'h6baf;
20995: douta=16'h530d;
20996: douta=16'h9471;
20997: douta=16'hbd34;
20998: douta=16'had36;
20999: douta=16'had35;
21000: douta=16'had35;
21001: douta=16'h9c94;
21002: douta=16'h94d5;
21003: douta=16'h8c73;
21004: douta=16'h8432;
21005: douta=16'h7bd1;
21006: douta=16'h7bd1;
21007: douta=16'h6b2e;
21008: douta=16'h630d;
21009: douta=16'h6acc;
21010: douta=16'hd5b3;
21011: douta=16'hcd94;
21012: douta=16'h9c94;
21013: douta=16'hacf5;
21014: douta=16'h9cd5;
21015: douta=16'h8453;
21016: douta=16'h8433;
21017: douta=16'h7c12;
21018: douta=16'h632f;
21019: douta=16'h632e;
21020: douta=16'h62ac;
21021: douta=16'h62cc;
21022: douta=16'h5229;
21023: douta=16'h72cb;
21024: douta=16'h52ef;
21025: douta=16'h9c31;
21026: douta=16'h8414;
21027: douta=16'h6b50;
21028: douta=16'h6b0d;
21029: douta=16'h5acc;
21030: douta=16'h62ac;
21031: douta=16'h524b;
21032: douta=16'h4a2a;
21033: douta=16'h41e8;
21034: douta=16'h5249;
21035: douta=16'hddf4;
21036: douta=16'hee55;
21037: douta=16'h6bb2;
21038: douta=16'h8c53;
21039: douta=16'h9495;
21040: douta=16'h7c32;
21041: douta=16'h73f2;
21042: douta=16'h73b1;
21043: douta=16'h632f;
21044: douta=16'h322c;
21045: douta=16'h424d;
21046: douta=16'h5aee;
21047: douta=16'h52ad;
21048: douta=16'h8bef;
21049: douta=16'hee97;
21050: douta=16'heed8;
21051: douta=16'heeb7;
21052: douta=16'hde37;
21053: douta=16'hcdf6;
21054: douta=16'hb555;
21055: douta=16'hbd96;
21056: douta=16'had15;
21057: douta=16'h9494;
21058: douta=16'ha515;
21059: douta=16'h9493;
21060: douta=16'h9473;
21061: douta=16'h8411;
21062: douta=16'h8412;
21063: douta=16'h7bf1;
21064: douta=16'h7c11;
21065: douta=16'h73b0;
21066: douta=16'h6b4f;
21067: douta=16'h73b1;
21068: douta=16'h630d;
21069: douta=16'h5249;
21070: douta=16'h5a8a;
21071: douta=16'h5a69;
21072: douta=16'h5a28;
21073: douta=16'hcd71;
21074: douta=16'he655;
21075: douta=16'hd5d3;
21076: douta=16'had34;
21077: douta=16'had14;
21078: douta=16'h9d15;
21079: douta=16'h94d5;
21080: douta=16'h7c54;
21081: douta=16'h7c54;
21082: douta=16'h7435;
21083: douta=16'h6392;
21084: douta=16'h4b10;
21085: douta=16'h42af;
21086: douta=16'h3a8e;
21087: douta=16'h29a9;
21088: douta=16'h6b91;
21089: douta=16'h31a8;
21090: douta=16'h0883;
21091: douta=16'h0884;
21092: douta=16'h10c5;
21093: douta=16'h29a9;
21094: douta=16'h6a24;
21095: douta=16'h8285;
21096: douta=16'h8285;
21097: douta=16'h7a84;
21098: douta=16'h7a65;
21099: douta=16'h7a44;
21100: douta=16'h7224;
21101: douta=16'h7224;
21102: douta=16'h7225;
21103: douta=16'h6a24;
21104: douta=16'h6204;
21105: douta=16'h6205;
21106: douta=16'h61e4;
21107: douta=16'h61e5;
21108: douta=16'h61e5;
21109: douta=16'h59e4;
21110: douta=16'h59c5;
21111: douta=16'h51a5;
21112: douta=16'h5144;
21113: douta=16'h4943;
21114: douta=16'h51a5;
21115: douta=16'h628a;
21116: douta=16'h62cb;
21117: douta=16'h736d;
21118: douta=16'h83f0;
21119: douta=16'h7c10;
21120: douta=16'hed8c;
21121: douta=16'he54b;
21122: douta=16'he54b;
21123: douta=16'hdd29;
21124: douta=16'hbc45;
21125: douta=16'h92c8;
21126: douta=16'he656;
21127: douta=16'hcd73;
21128: douta=16'hcd92;
21129: douta=16'hddd4;
21130: douta=16'he677;
21131: douta=16'hddf6;
21132: douta=16'h8433;
21133: douta=16'h7c55;
21134: douta=16'h84b7;
21135: douta=16'h8475;
21136: douta=16'h8496;
21137: douta=16'h8496;
21138: douta=16'h9d39;
21139: douta=16'h29eb;
21140: douta=16'h326d;
21141: douta=16'h3a8e;
21142: douta=16'h328e;
21143: douta=16'h3aae;
21144: douta=16'h3a8e;
21145: douta=16'h3aae;
21146: douta=16'h3a8d;
21147: douta=16'h21ca;
21148: douta=16'h29ea;
21149: douta=16'h29ea;
21150: douta=16'h29c9;
21151: douta=16'h18e4;
21152: douta=16'h10a3;
21153: douta=16'h18c4;
21154: douta=16'h2145;
21155: douta=16'h2967;
21156: douta=16'h31c9;
21157: douta=16'h422a;
21158: douta=16'h422a;
21159: douta=16'h4a4b;
21160: douta=16'h422a;
21161: douta=16'h39ea;
21162: douta=16'h31c9;
21163: douta=16'h29a8;
21164: douta=16'h2146;
21165: douta=16'h1905;
21166: douta=16'h10e6;
21167: douta=16'h10e5;
21168: douta=16'h0883;
21169: douta=16'h3a4c;
21170: douta=16'h42ee;
21171: douta=16'h4aed;
21172: douta=16'h532f;
21173: douta=16'h52ed;
21174: douta=16'h530d;
21175: douta=16'h5b2e;
21176: douta=16'h5b0e;
21177: douta=16'h636f;
21178: douta=16'h636f;
21179: douta=16'h638f;
21180: douta=16'h6bb0;
21181: douta=16'h6bd0;
21182: douta=16'h6bb0;
21183: douta=16'h636f;
21184: douta=16'h6b8f;
21185: douta=16'h6bb0;
21186: douta=16'h636f;
21187: douta=16'h5b4e;
21188: douta=16'h638f;
21189: douta=16'h636e;
21190: douta=16'h8410;
21191: douta=16'h9cb3;
21192: douta=16'h9cb3;
21193: douta=16'h9493;
21194: douta=16'h9493;
21195: douta=16'h8c32;
21196: douta=16'h83f1;
21197: douta=16'h7bf1;
21198: douta=16'h736f;
21199: douta=16'h730d;
21200: douta=16'h93ee;
21201: douta=16'hf6d6;
21202: douta=16'had15;
21203: douta=16'hacf5;
21204: douta=16'h94b6;
21205: douta=16'h8c74;
21206: douta=16'h8c95;
21207: douta=16'h7390;
21208: douta=16'h7390;
21209: douta=16'h7b90;
21210: douta=16'h6b0d;
21211: douta=16'h628b;
21212: douta=16'h62cc;
21213: douta=16'h5a6b;
21214: douta=16'hb4d3;
21215: douta=16'hacd3;
21216: douta=16'h428d;
21217: douta=16'h83d1;
21218: douta=16'h6b4f;
21219: douta=16'h6b2e;
21220: douta=16'h41c8;
21221: douta=16'h2988;
21222: douta=16'h39e8;
21223: douta=16'h420a;
21224: douta=16'h2968;
21225: douta=16'h732d;
21226: douta=16'hc574;
21227: douta=16'hbd13;
21228: douta=16'hacf5;
21229: douta=16'h6391;
21230: douta=16'h6370;
21231: douta=16'h8c74;
21232: douta=16'h6b70;
21233: douta=16'h6b2f;
21234: douta=16'h6b2e;
21235: douta=16'h6b0e;
21236: douta=16'h736f;
21237: douta=16'h6b4f;
21238: douta=16'ha470;
21239: douta=16'hd5f4;
21240: douta=16'heeb7;
21241: douta=16'he677;
21242: douta=16'hcdf7;
21243: douta=16'hb577;
21244: douta=16'hc5d7;
21245: douta=16'hc5b6;
21246: douta=16'hbd96;
21247: douta=16'hb556;
21248: douta=16'ha515;
21249: douta=16'h8c74;
21250: douta=16'h8453;
21251: douta=16'h9472;
21252: douta=16'h9473;
21253: douta=16'h8c73;
21254: douta=16'h8432;
21255: douta=16'h73b0;
21256: douta=16'h7c12;
21257: douta=16'h62ee;
21258: douta=16'h630d;
21259: douta=16'h730b;
21260: douta=16'ha46f;
21261: douta=16'hd5d3;
21262: douta=16'hde55;
21263: douta=16'he634;
21264: douta=16'he655;
21265: douta=16'hde15;
21266: douta=16'hde34;
21267: douta=16'hde15;
21268: douta=16'had14;
21269: douta=16'had14;
21270: douta=16'ha4f5;
21271: douta=16'h8cb5;
21272: douta=16'h7c34;
21273: douta=16'h7414;
21274: douta=16'h7c75;
21275: douta=16'h63f4;
21276: douta=16'h5351;
21277: douta=16'h42cf;
21278: douta=16'h42ae;
21279: douta=16'h29aa;
21280: douta=16'h0064;
21281: douta=16'h7c54;
21282: douta=16'h1927;
21283: douta=16'h1906;
21284: douta=16'h18e5;
21285: douta=16'h1927;
21286: douta=16'h8ac5;
21287: douta=16'h7aa5;
21288: douta=16'h8285;
21289: douta=16'h7a84;
21290: douta=16'h7a65;
21291: douta=16'h7a64;
21292: douta=16'h7224;
21293: douta=16'h7224;
21294: douta=16'h6a25;
21295: douta=16'h6a04;
21296: douta=16'h61c4;
21297: douta=16'h61a4;
21298: douta=16'h59a4;
21299: douta=16'h59e5;
21300: douta=16'h6a88;
21301: douta=16'h7b8c;
21302: douta=16'h8c51;
21303: douta=16'h9492;
21304: douta=16'ha534;
21305: douta=16'h9d13;
21306: douta=16'h94b1;
21307: douta=16'h83ee;
21308: douta=16'h7b8d;
21309: douta=16'h6aea;
21310: douta=16'h5a69;
21311: douta=16'h4a27;
21312: douta=16'hed6b;
21313: douta=16'he54a;
21314: douta=16'he52a;
21315: douta=16'hdd2a;
21316: douta=16'hcc44;
21317: douta=16'hcd11;
21318: douta=16'hddf4;
21319: douta=16'hd594;
21320: douta=16'hddb3;
21321: douta=16'hee76;
21322: douta=16'hde57;
21323: douta=16'hd5f6;
21324: douta=16'h73f2;
21325: douta=16'h7c75;
21326: douta=16'h8496;
21327: douta=16'h73d2;
21328: douta=16'h8cb6;
21329: douta=16'h8cd7;
21330: douta=16'h94f8;
21331: douta=16'h29eb;
21332: douta=16'h322d;
21333: douta=16'h322c;
21334: douta=16'h3aae;
21335: douta=16'h3a8e;
21336: douta=16'h3a8e;
21337: douta=16'h3a4e;
21338: douta=16'h324d;
21339: douta=16'h2a0b;
21340: douta=16'h2168;
21341: douta=16'h29ea;
21342: douta=16'h29ca;
21343: douta=16'h18e5;
21344: douta=16'h10c3;
21345: douta=16'h18e5;
21346: douta=16'h31c9;
21347: douta=16'h39ea;
21348: douta=16'h39e9;
21349: douta=16'h52ac;
21350: douta=16'h62cd;
21351: douta=16'h62ed;
21352: douta=16'h52ac;
21353: douta=16'h528c;
21354: douta=16'h4a8d;
21355: douta=16'h3a2c;
21356: douta=16'h31ea;
21357: douta=16'h29a9;
21358: douta=16'h1106;
21359: douta=16'h10c5;
21360: douta=16'h10e4;
21361: douta=16'h10a4;
21362: douta=16'h1946;
21363: douta=16'h3a8c;
21364: douta=16'h4aad;
21365: douta=16'h426b;
21366: douta=16'h4aac;
21367: douta=16'h5b2e;
21368: douta=16'h4acd;
21369: douta=16'h636f;
21370: douta=16'h6b90;
21371: douta=16'h638f;
21372: douta=16'h638f;
21373: douta=16'h6bd0;
21374: douta=16'h636f;
21375: douta=16'h6bb0;
21376: douta=16'h6bb0;
21377: douta=16'h6bb0;
21378: douta=16'h6b8f;
21379: douta=16'h638f;
21380: douta=16'h6baf;
21381: douta=16'h6baf;
21382: douta=16'h6b6e;
21383: douta=16'h73cf;
21384: douta=16'h9452;
21385: douta=16'ha4d4;
21386: douta=16'ha4d4;
21387: douta=16'h9473;
21388: douta=16'h7bf1;
21389: douta=16'h736e;
21390: douta=16'h6b2d;
21391: douta=16'hd593;
21392: douta=16'hcd72;
21393: douta=16'he655;
21394: douta=16'ha4f5;
21395: douta=16'had36;
21396: douta=16'h94b6;
21397: douta=16'h9496;
21398: douta=16'h8c74;
21399: douta=16'h7bf1;
21400: douta=16'h736f;
21401: douta=16'h738f;
21402: douta=16'h6b0e;
21403: douta=16'h6acc;
21404: douta=16'h524a;
21405: douta=16'h5a6b;
21406: douta=16'h9c73;
21407: douta=16'h9453;
21408: douta=16'h4a8c;
21409: douta=16'h83d0;
21410: douta=16'h62ed;
21411: douta=16'h62cc;
21412: douta=16'h5a6a;
21413: douta=16'h41c8;
21414: douta=16'h2147;
21415: douta=16'h2966;
21416: douta=16'h422a;
21417: douta=16'hb4f4;
21418: douta=16'h94b4;
21419: douta=16'had15;
21420: douta=16'ha4f5;
21421: douta=16'h7bf3;
21422: douta=16'h5b30;
21423: douta=16'h8412;
21424: douta=16'h6b2f;
21425: douta=16'h6b2e;
21426: douta=16'h6b0e;
21427: douta=16'h630e;
21428: douta=16'h5aee;
21429: douta=16'hacd2;
21430: douta=16'he697;
21431: douta=16'heed9;
21432: douta=16'he698;
21433: douta=16'hd616;
21434: douta=16'hc5f7;
21435: douta=16'hb577;
21436: douta=16'hb597;
21437: douta=16'hb577;
21438: douta=16'hb577;
21439: douta=16'hbdb7;
21440: douta=16'hb597;
21441: douta=16'h94d5;
21442: douta=16'h7bf3;
21443: douta=16'h7c33;
21444: douta=16'h8c52;
21445: douta=16'h8432;
21446: douta=16'h8432;
21447: douta=16'h7bf2;
21448: douta=16'h5acc;
21449: douta=16'ha46f;
21450: douta=16'hc511;
21451: douta=16'hcd93;
21452: douta=16'hd5d2;
21453: douta=16'he635;
21454: douta=16'hde35;
21455: douta=16'he676;
21456: douta=16'he676;
21457: douta=16'hde15;
21458: douta=16'hc594;
21459: douta=16'hc574;
21460: douta=16'ha4f5;
21461: douta=16'ha515;
21462: douta=16'ha516;
21463: douta=16'h8c95;
21464: douta=16'h7c34;
21465: douta=16'h7434;
21466: douta=16'h7c55;
21467: douta=16'h7414;
21468: douta=16'h63b3;
21469: douta=16'h5310;
21470: douta=16'h42cf;
21471: douta=16'h31ca;
21472: douta=16'h2988;
21473: douta=16'h5351;
21474: douta=16'h5b71;
21475: douta=16'h1906;
21476: douta=16'h1906;
21477: douta=16'h2167;
21478: douta=16'h7a66;
21479: douta=16'h8285;
21480: douta=16'h8285;
21481: douta=16'h7a64;
21482: douta=16'h7a44;
21483: douta=16'h7244;
21484: douta=16'h6a04;
21485: douta=16'h69e4;
21486: douta=16'h61c4;
21487: douta=16'h6205;
21488: douta=16'h6a66;
21489: douta=16'h72c8;
21490: douta=16'h8c0e;
21491: douta=16'h944f;
21492: douta=16'ha513;
21493: douta=16'had53;
21494: douta=16'ha513;
21495: douta=16'ha4d2;
21496: douta=16'h83ee;
21497: douta=16'h734b;
21498: douta=16'h62c9;
21499: douta=16'h5207;
21500: douta=16'h4985;
21501: douta=16'h4164;
21502: douta=16'h4124;
21503: douta=16'h3944;
21504: douta=16'he506;
21505: douta=16'hdd06;
21506: douta=16'he4e6;
21507: douta=16'hdce6;
21508: douta=16'hff7d;
21509: douta=16'hf6f8;
21510: douta=16'hff39;
21511: douta=16'he676;
21512: douta=16'heeb8;
21513: douta=16'hff7c;
21514: douta=16'hde36;
21515: douta=16'had15;
21516: douta=16'h73f3;
21517: douta=16'h8c76;
21518: douta=16'h73f2;
21519: douta=16'h5aee;
21520: douta=16'h9539;
21521: douta=16'h8cb7;
21522: douta=16'h84b6;
21523: douta=16'h29eb;
21524: douta=16'h322c;
21525: douta=16'h324d;
21526: douta=16'h326e;
21527: douta=16'h3a8e;
21528: douta=16'h3aaf;
21529: douta=16'h326d;
21530: douta=16'h3a6e;
21531: douta=16'h1927;
21532: douta=16'h1926;
21533: douta=16'h1947;
21534: douta=16'h2189;
21535: douta=16'h29a9;
21536: douta=16'h2168;
21537: douta=16'h31ca;
21538: douta=16'h31c9;
21539: douta=16'h31a8;
21540: douta=16'h29a8;
21541: douta=16'h3a0a;
21542: douta=16'h422a;
21543: douta=16'h424b;
21544: douta=16'h3a0a;
21545: douta=16'h3a0a;
21546: douta=16'h3a2b;
21547: douta=16'h424c;
21548: douta=16'h39eb;
21549: douta=16'h31eb;
21550: douta=16'h3a2b;
21551: douta=16'h3a2b;
21552: douta=16'h3a0a;
21553: douta=16'h18e5;
21554: douta=16'h1084;
21555: douta=16'h10a4;
21556: douta=16'h31c9;
21557: douta=16'h4aac;
21558: douta=16'h4aac;
21559: douta=16'h4acd;
21560: douta=16'h52ed;
21561: douta=16'h530d;
21562: douta=16'h5b2e;
21563: douta=16'h5b4e;
21564: douta=16'h5b2e;
21565: douta=16'h636f;
21566: douta=16'h5b4e;
21567: douta=16'h5b4e;
21568: douta=16'h636f;
21569: douta=16'h636f;
21570: douta=16'h6b90;
21571: douta=16'h6bb0;
21572: douta=16'h73d0;
21573: douta=16'h6baf;
21574: douta=16'h73af;
21575: douta=16'h73cf;
21576: douta=16'h6b8f;
21577: douta=16'h6b8f;
21578: douta=16'h6b8e;
21579: douta=16'h7baf;
21580: douta=16'h7bcf;
21581: douta=16'h6b4d;
21582: douta=16'h5aeb;
21583: douta=16'h9c92;
21584: douta=16'ha4b4;
21585: douta=16'ha4f5;
21586: douta=16'h9453;
21587: douta=16'h8412;
21588: douta=16'h83f1;
21589: douta=16'h7b8f;
21590: douta=16'h734e;
21591: douta=16'h7b6e;
21592: douta=16'h734d;
21593: douta=16'h732d;
21594: douta=16'h6acb;
21595: douta=16'ha451;
21596: douta=16'hbd13;
21597: douta=16'hacd3;
21598: douta=16'h8433;
21599: douta=16'h73b1;
21600: douta=16'h62ed;
21601: douta=16'h7bf1;
21602: douta=16'h62cc;
21603: douta=16'h62aa;
21604: douta=16'h628a;
21605: douta=16'h49c7;
21606: douta=16'h838e;
21607: douta=16'h6b71;
21608: douta=16'h8c74;
21609: douta=16'hacf5;
21610: douta=16'h9cd5;
21611: douta=16'h8412;
21612: douta=16'h7bf2;
21613: douta=16'h4aad;
21614: douta=16'h424c;
21615: douta=16'h3a4c;
21616: douta=16'h62ed;
21617: douta=16'h4a6b;
21618: douta=16'h5aad;
21619: douta=16'hb4b2;
21620: douta=16'hf6d8;
21621: douta=16'hcdb5;
21622: douta=16'hde56;
21623: douta=16'hcdf6;
21624: douta=16'hc5b6;
21625: douta=16'had36;
21626: douta=16'ha4f5;
21627: douta=16'h9cf5;
21628: douta=16'h9494;
21629: douta=16'h9cf5;
21630: douta=16'h9cd6;
21631: douta=16'h9cf6;
21632: douta=16'h94b5;
21633: douta=16'h8453;
21634: douta=16'h7bf2;
21635: douta=16'h6b90;
21636: douta=16'h6b90;
21637: douta=16'h62aa;
21638: douta=16'h836c;
21639: douta=16'ha44e;
21640: douta=16'hc551;
21641: douta=16'hb4d0;
21642: douta=16'h834c;
21643: douta=16'hac50;
21644: douta=16'hacf1;
21645: douta=16'hcd93;
21646: douta=16'hde34;
21647: douta=16'he655;
21648: douta=16'hb513;
21649: douta=16'h9cb3;
21650: douta=16'ha4f5;
21651: douta=16'ha515;
21652: douta=16'h8c94;
21653: douta=16'h8c95;
21654: douta=16'h8474;
21655: douta=16'h7c13;
21656: douta=16'h7c34;
21657: douta=16'h7413;
21658: douta=16'h6bb3;
21659: douta=16'h63b2;
21660: douta=16'h63b3;
21661: douta=16'h5331;
21662: douta=16'h4aaf;
21663: douta=16'h428d;
21664: douta=16'h320b;
21665: douta=16'h6c13;
21666: douta=16'h428d;
21667: douta=16'h1906;
21668: douta=16'h1906;
21669: douta=16'h2127;
21670: douta=16'h1927;
21671: douta=16'h9beb;
21672: douta=16'h9c0b;
21673: douta=16'hc572;
21674: douta=16'hce13;
21675: douta=16'hd612;
21676: douta=16'hc5b1;
21677: douta=16'hbd70;
21678: douta=16'ha4ad;
21679: douta=16'h8bab;
21680: douta=16'h7b09;
21681: douta=16'h72c8;
21682: douta=16'h59c5;
21683: douta=16'h51a4;
21684: douta=16'h59a5;
21685: douta=16'h51a5;
21686: douta=16'h59c5;
21687: douta=16'h51c5;
21688: douta=16'h51c5;
21689: douta=16'h51c5;
21690: douta=16'h4985;
21691: douta=16'h4985;
21692: douta=16'h4985;
21693: douta=16'h4985;
21694: douta=16'h4986;
21695: douta=16'h4985;
21696: douta=16'hdca3;
21697: douta=16'hd4a3;
21698: douta=16'hd484;
21699: douta=16'hcc20;
21700: douta=16'hf6f8;
21701: douta=16'hff3a;
21702: douta=16'hff3a;
21703: douta=16'heeb8;
21704: douta=16'hff3a;
21705: douta=16'hff9c;
21706: douta=16'hb555;
21707: douta=16'h8433;
21708: douta=16'h8455;
21709: douta=16'h8c95;
21710: douta=16'h6b2f;
21711: douta=16'h7b91;
21712: douta=16'h8c76;
21713: douta=16'h9518;
21714: douta=16'h5330;
21715: douta=16'h21a9;
21716: douta=16'h21ca;
21717: douta=16'h2a2c;
21718: douta=16'h324c;
21719: douta=16'h3a6d;
21720: douta=16'h322c;
21721: douta=16'h3a4d;
21722: douta=16'h42af;
21723: douta=16'h1127;
21724: douta=16'h1968;
21725: douta=16'h1947;
21726: douta=16'h2147;
21727: douta=16'h1926;
21728: douta=16'h1927;
21729: douta=16'h31c9;
21730: douta=16'h2988;
21731: douta=16'h31c9;
21732: douta=16'h39ea;
21733: douta=16'h424c;
21734: douta=16'h426c;
21735: douta=16'h424c;
21736: douta=16'h426c;
21737: douta=16'h4a8c;
21738: douta=16'h4a8d;
21739: douta=16'h3a2b;
21740: douta=16'h424c;
21741: douta=16'h3a2b;
21742: douta=16'h31ca;
21743: douta=16'h31c9;
21744: douta=16'h3189;
21745: douta=16'h422a;
21746: douta=16'h29a8;
21747: douta=16'h1084;
21748: douta=16'h1906;
21749: douta=16'h320a;
21750: douta=16'h3a2b;
21751: douta=16'h4acc;
21752: douta=16'h52cd;
21753: douta=16'h4acd;
21754: douta=16'h52ed;
21755: douta=16'h5b2e;
21756: douta=16'h5b2e;
21757: douta=16'h5b4e;
21758: douta=16'h5b2e;
21759: douta=16'h634f;
21760: douta=16'h5b4e;
21761: douta=16'h636f;
21762: douta=16'h6baf;
21763: douta=16'h6baf;
21764: douta=16'h73f0;
21765: douta=16'h73af;
21766: douta=16'h634d;
21767: douta=16'h634d;
21768: douta=16'h632d;
21769: douta=16'h634e;
21770: douta=16'h6b6e;
21771: douta=16'h6b8e;
21772: douta=16'h6b6e;
21773: douta=16'h7baf;
21774: douta=16'h7bae;
21775: douta=16'h736d;
21776: douta=16'h736d;
21777: douta=16'h83ef;
21778: douta=16'h8c0f;
21779: douta=16'h8bcf;
21780: douta=16'h8bf0;
21781: douta=16'h838f;
21782: douta=16'h736d;
21783: douta=16'h732c;
21784: douta=16'h730b;
21785: douta=16'h836d;
21786: douta=16'ha4b3;
21787: douta=16'h8412;
21788: douta=16'h8c32;
21789: douta=16'h7bf1;
21790: douta=16'h734d;
21791: douta=16'h732d;
21792: douta=16'h6b2c;
21793: douta=16'h6aab;
21794: douta=16'h6acb;
21795: douta=16'h62ab;
21796: douta=16'h730b;
21797: douta=16'hc574;
21798: douta=16'h8413;
21799: douta=16'h6b50;
21800: douta=16'h9495;
21801: douta=16'ha516;
21802: douta=16'h8453;
21803: douta=16'h7bf1;
21804: douta=16'h7bd1;
21805: douta=16'h7390;
21806: douta=16'h734f;
21807: douta=16'h62cd;
21808: douta=16'h422b;
21809: douta=16'hb535;
21810: douta=16'ha493;
21811: douta=16'hf6f8;
21812: douta=16'hd5f6;
21813: douta=16'hbd96;
21814: douta=16'ha515;
21815: douta=16'had56;
21816: douta=16'ha516;
21817: douta=16'h8c74;
21818: douta=16'h7bf1;
21819: douta=16'h7bd1;
21820: douta=16'h8c94;
21821: douta=16'h7bf2;
21822: douta=16'h8c94;
21823: douta=16'h7c33;
21824: douta=16'h7c12;
21825: douta=16'h8433;
21826: douta=16'h5aad;
21827: douta=16'h524a;
21828: douta=16'h5a69;
21829: douta=16'hcd92;
21830: douta=16'hddf4;
21831: douta=16'hde14;
21832: douta=16'he655;
21833: douta=16'hde35;
21834: douta=16'he675;
21835: douta=16'hd5f4;
21836: douta=16'hacd1;
21837: douta=16'hacb2;
21838: douta=16'hacd4;
21839: douta=16'hacb4;
21840: douta=16'hb514;
21841: douta=16'had14;
21842: douta=16'h9cb4;
21843: douta=16'h9cb4;
21844: douta=16'h8c54;
21845: douta=16'h8453;
21846: douta=16'h73f1;
21847: douta=16'h73d2;
21848: douta=16'h73b2;
21849: douta=16'h6bb1;
21850: douta=16'h6371;
21851: douta=16'h5b51;
21852: douta=16'h6371;
21853: douta=16'h3a4c;
21854: douta=16'h6b2d;
21855: douta=16'h94b4;
21856: douta=16'h5aed;
21857: douta=16'h52cc;
21858: douta=16'h3a4c;
21859: douta=16'h10a4;
21860: douta=16'h1926;
21861: douta=16'h1905;
21862: douta=16'h18c4;
21863: douta=16'h83cc;
21864: douta=16'hbced;
21865: douta=16'h936a;
21866: douta=16'h82c7;
21867: douta=16'h7265;
21868: douta=16'h69e4;
21869: douta=16'h61c4;
21870: douta=16'h69e4;
21871: douta=16'h61e5;
21872: douta=16'h61e5;
21873: douta=16'h61e5;
21874: douta=16'h59e4;
21875: douta=16'h59e5;
21876: douta=16'h59c5;
21877: douta=16'h51c5;
21878: douta=16'h51a5;
21879: douta=16'h59c5;
21880: douta=16'h51a5;
21881: douta=16'h4985;
21882: douta=16'h49a5;
21883: douta=16'h4985;
21884: douta=16'h49a5;
21885: douta=16'h4985;
21886: douta=16'h4986;
21887: douta=16'h4186;
21888: douta=16'hcc01;
21889: douta=16'hd443;
21890: douta=16'hd462;
21891: douta=16'hdccb;
21892: douta=16'hf6f9;
21893: douta=16'hff5b;
21894: douta=16'hff3a;
21895: douta=16'hf6b8;
21896: douta=16'hff7b;
21897: douta=16'hff7b;
21898: douta=16'h9493;
21899: douta=16'h7c13;
21900: douta=16'h8475;
21901: douta=16'h8cb6;
21902: douta=16'h6b2e;
21903: douta=16'h8412;
21904: douta=16'h8cb6;
21905: douta=16'h94d7;
21906: douta=16'h322b;
21907: douta=16'h2168;
21908: douta=16'h2189;
21909: douta=16'h2189;
21910: douta=16'h322c;
21911: douta=16'h3a8e;
21912: douta=16'h324d;
21913: douta=16'h3a4e;
21914: douta=16'h328e;
21915: douta=16'h1968;
21916: douta=16'h1947;
21917: douta=16'h2147;
21918: douta=16'h2147;
21919: douta=16'h1905;
21920: douta=16'h10a5;
21921: douta=16'h31ca;
21922: douta=16'h2987;
21923: douta=16'h39e9;
21924: douta=16'h424b;
21925: douta=16'h424c;
21926: douta=16'h426c;
21927: douta=16'h3a4c;
21928: douta=16'h3a2c;
21929: douta=16'h3a2c;
21930: douta=16'h426c;
21931: douta=16'h4ace;
21932: douta=16'h426c;
21933: douta=16'h426d;
21934: douta=16'h426c;
21935: douta=16'h3a0a;
21936: douta=16'h3188;
21937: douta=16'h39ea;
21938: douta=16'h422b;
21939: douta=16'h18e5;
21940: douta=16'h0883;
21941: douta=16'h31ca;
21942: douta=16'h3a2b;
21943: douta=16'h4acd;
21944: douta=16'h52ed;
21945: douta=16'h52ed;
21946: douta=16'h530d;
21947: douta=16'h530e;
21948: douta=16'h530d;
21949: douta=16'h5b2e;
21950: douta=16'h5b2e;
21951: douta=16'h5b4e;
21952: douta=16'h5b0d;
21953: douta=16'h5b4e;
21954: douta=16'h73d0;
21955: douta=16'h6b90;
21956: douta=16'h6b8f;
21957: douta=16'h6b4e;
21958: douta=16'h634d;
21959: douta=16'h634d;
21960: douta=16'h634e;
21961: douta=16'h73af;
21962: douta=16'h73cf;
21963: douta=16'h73cf;
21964: douta=16'h6b8e;
21965: douta=16'h738e;
21966: douta=16'h6b4d;
21967: douta=16'h7bae;
21968: douta=16'h7bae;
21969: douta=16'h736d;
21970: douta=16'h8c10;
21971: douta=16'h8bf0;
21972: douta=16'h83cf;
21973: douta=16'h8bef;
21974: douta=16'h8bcf;
21975: douta=16'h838e;
21976: douta=16'h7b6d;
21977: douta=16'h8bef;
21978: douta=16'ha4b4;
21979: douta=16'h7baf;
21980: douta=16'h838f;
21981: douta=16'h7b6e;
21982: douta=16'h6b0c;
21983: douta=16'h730c;
21984: douta=16'h6acc;
21985: douta=16'h6aaa;
21986: douta=16'h6aab;
21987: douta=16'h6a8a;
21988: douta=16'hcd71;
21989: douta=16'h8412;
21990: douta=16'h7bb0;
21991: douta=16'h62cd;
21992: douta=16'h7bb0;
21993: douta=16'h8411;
21994: douta=16'h83d1;
21995: douta=16'h7bf1;
21996: douta=16'h73b0;
21997: douta=16'h734f;
21998: douta=16'h6b2e;
21999: douta=16'h62ed;
22000: douta=16'h9c70;
22001: douta=16'h8c73;
22002: douta=16'hacb1;
22003: douta=16'hde36;
22004: douta=16'hcdd6;
22005: douta=16'hc596;
22006: douta=16'ha4f5;
22007: douta=16'h9cd5;
22008: douta=16'h9cd5;
22009: douta=16'h9494;
22010: douta=16'h7bf0;
22011: douta=16'h7bb0;
22012: douta=16'h8c53;
22013: douta=16'h8433;
22014: douta=16'h73d1;
22015: douta=16'h8453;
22016: douta=16'h7c12;
22017: douta=16'h6b4f;
22018: douta=16'h6aeb;
22019: douta=16'hbd73;
22020: douta=16'hc572;
22021: douta=16'he656;
22022: douta=16'he676;
22023: douta=16'hd5f4;
22024: douta=16'hcd93;
22025: douta=16'hd5d4;
22026: douta=16'hcd93;
22027: douta=16'hd5f4;
22028: douta=16'he655;
22029: douta=16'hbd32;
22030: douta=16'h9c72;
22031: douta=16'h9c93;
22032: douta=16'h83f1;
22033: douta=16'h9cb3;
22034: douta=16'h9c94;
22035: douta=16'h8c73;
22036: douta=16'h8453;
22037: douta=16'h8454;
22038: douta=16'h7c12;
22039: douta=16'h6350;
22040: douta=16'h6b91;
22041: douta=16'h6b91;
22042: douta=16'h6371;
22043: douta=16'h6330;
22044: douta=16'h41e7;
22045: douta=16'h9c4e;
22046: douta=16'hbd72;
22047: douta=16'h4aae;
22048: douta=16'h52cd;
22049: douta=16'h52cc;
22050: douta=16'h3a4c;
22051: douta=16'h10c4;
22052: douta=16'h0863;
22053: douta=16'h1083;
22054: douta=16'h1906;
22055: douta=16'h2127;
22056: douta=16'h7aa7;
22057: douta=16'h7224;
22058: douta=16'h7224;
22059: douta=16'h7225;
22060: douta=16'h7225;
22061: douta=16'h7225;
22062: douta=16'h6a25;
22063: douta=16'h6204;
22064: douta=16'h6205;
22065: douta=16'h61e5;
22066: douta=16'h61e5;
22067: douta=16'h59c5;
22068: douta=16'h59e5;
22069: douta=16'h59c5;
22070: douta=16'h51c5;
22071: douta=16'h51c5;
22072: douta=16'h51a5;
22073: douta=16'h51a5;
22074: douta=16'h49a5;
22075: douta=16'h4985;
22076: douta=16'h4985;
22077: douta=16'h4986;
22078: douta=16'h41a5;
22079: douta=16'h4165;
22080: douta=16'hf718;
22081: douta=16'h71a1;
22082: douta=16'h89e1;
22083: douta=16'hffbd;
22084: douta=16'hff3b;
22085: douta=16'hff3a;
22086: douta=16'hff3a;
22087: douta=16'hf6f8;
22088: douta=16'hff9c;
22089: douta=16'heeb7;
22090: douta=16'h9494;
22091: douta=16'h8c53;
22092: douta=16'h8cb5;
22093: douta=16'h8433;
22094: douta=16'h8c53;
22095: douta=16'h8c74;
22096: douta=16'h8cb5;
22097: douta=16'h8475;
22098: douta=16'h10e5;
22099: douta=16'h2189;
22100: douta=16'h21aa;
22101: douta=16'h21a9;
22102: douta=16'h1967;
22103: douta=16'h1126;
22104: douta=16'h1948;
22105: douta=16'h1947;
22106: douta=16'h1968;
22107: douta=16'h2168;
22108: douta=16'h1106;
22109: douta=16'h1948;
22110: douta=16'h2168;
22111: douta=16'h1967;
22112: douta=16'h29a9;
22113: douta=16'h18e6;
22114: douta=16'h2168;
22115: douta=16'h29a9;
22116: douta=16'h31c9;
22117: douta=16'h426d;
22118: douta=16'h31ea;
22119: douta=16'h31ea;
22120: douta=16'h4a6c;
22121: douta=16'h424c;
22122: douta=16'h424c;
22123: douta=16'h320b;
22124: douta=16'h3a0b;
22125: douta=16'h3a0b;
22126: douta=16'h3a2c;
22127: douta=16'h39ea;
22128: douta=16'h420a;
22129: douta=16'h424a;
22130: douta=16'h2968;
22131: douta=16'h39e9;
22132: douta=16'h2967;
22133: douta=16'h31ca;
22134: douta=16'h3a2b;
22135: douta=16'h4aad;
22136: douta=16'h4aed;
22137: douta=16'h4aad;
22138: douta=16'h4acd;
22139: douta=16'h530d;
22140: douta=16'h4aac;
22141: douta=16'h4aac;
22142: douta=16'h4aac;
22143: douta=16'h4aab;
22144: douta=16'h5b0d;
22145: douta=16'h632e;
22146: douta=16'h636e;
22147: douta=16'h6b8f;
22148: douta=16'h6b6f;
22149: douta=16'h6b8f;
22150: douta=16'h632e;
22151: douta=16'h634d;
22152: douta=16'h5acb;
22153: douta=16'h62cb;
22154: douta=16'h62cb;
22155: douta=16'h62cb;
22156: douta=16'h6b0c;
22157: douta=16'h62cb;
22158: douta=16'h630c;
22159: douta=16'h6aeb;
22160: douta=16'h62cb;
22161: douta=16'h6b0c;
22162: douta=16'h630c;
22163: douta=16'h6b0c;
22164: douta=16'h6b2c;
22165: douta=16'h6b0c;
22166: douta=16'h62cb;
22167: douta=16'h6b0b;
22168: douta=16'h734c;
22169: douta=16'h6b0b;
22170: douta=16'h732c;
22171: douta=16'h732d;
22172: douta=16'h83ef;
22173: douta=16'h9431;
22174: douta=16'h8bef;
22175: douta=16'h9430;
22176: douta=16'h9491;
22177: douta=16'h8c50;
22178: douta=16'hb597;
22179: douta=16'hb5b6;
22180: douta=16'h7baf;
22181: douta=16'h7b90;
22182: douta=16'h736f;
22183: douta=16'h632e;
22184: douta=16'h6b2e;
22185: douta=16'h7b8e;
22186: douta=16'h7baf;
22187: douta=16'h732e;
22188: douta=16'h732e;
22189: douta=16'hb4b0;
22190: douta=16'hc571;
22191: douta=16'he697;
22192: douta=16'h9cf5;
22193: douta=16'hbd55;
22194: douta=16'hd616;
22195: douta=16'had57;
22196: douta=16'h9d16;
22197: douta=16'h8c94;
22198: douta=16'h8454;
22199: douta=16'h73f2;
22200: douta=16'h8432;
22201: douta=16'h73b0;
22202: douta=16'h52cd;
22203: douta=16'h5aef;
22204: douta=16'h52ac;
22205: douta=16'h5aad;
22206: douta=16'h526a;
22207: douta=16'h730b;
22208: douta=16'h8bee;
22209: douta=16'hde13;
22210: douta=16'he697;
22211: douta=16'hbd54;
22212: douta=16'hbd34;
22213: douta=16'hddf5;
22214: douta=16'hcdb6;
22215: douta=16'hcdd4;
22216: douta=16'ha4b4;
22217: douta=16'h9473;
22218: douta=16'h9452;
22219: douta=16'h9432;
22220: douta=16'h7bd1;
22221: douta=16'h73b0;
22222: douta=16'h8411;
22223: douta=16'h8c53;
22224: douta=16'h8412;
22225: douta=16'h8c33;
22226: douta=16'h8c32;
22227: douta=16'h7bf1;
22228: douta=16'h7390;
22229: douta=16'h7390;
22230: douta=16'h6b4f;
22231: douta=16'h630e;
22232: douta=16'h526a;
22233: douta=16'h41c8;
22234: douta=16'h732b;
22235: douta=16'hac6f;
22236: douta=16'hcdd2;
22237: douta=16'hc573;
22238: douta=16'h9c52;
22239: douta=16'h6390;
22240: douta=16'h6b90;
22241: douta=16'h5b2f;
22242: douta=16'h29a9;
22243: douta=16'h18e5;
22244: douta=16'h1926;
22245: douta=16'h29a9;
22246: douta=16'h10e5;
22247: douta=16'h18e4;
22248: douta=16'h10e5;
22249: douta=16'h8286;
22250: douta=16'h7a65;
22251: douta=16'h7a65;
22252: douta=16'h7225;
22253: douta=16'h7245;
22254: douta=16'h6a04;
22255: douta=16'h61e5;
22256: douta=16'h6205;
22257: douta=16'h61e5;
22258: douta=16'h59c5;
22259: douta=16'h59e5;
22260: douta=16'h59c5;
22261: douta=16'h51c5;
22262: douta=16'h51a5;
22263: douta=16'h51c5;
22264: douta=16'h51a5;
22265: douta=16'h49a5;
22266: douta=16'h49a5;
22267: douta=16'h49a5;
22268: douta=16'h4185;
22269: douta=16'h4985;
22270: douta=16'h4185;
22271: douta=16'h4165;
22272: douta=16'he653;
22273: douta=16'hcd6c;
22274: douta=16'hf6b7;
22275: douta=16'hf6f8;
22276: douta=16'hff5b;
22277: douta=16'hff3a;
22278: douta=16'hf719;
22279: douta=16'hff5b;
22280: douta=16'hf718;
22281: douta=16'he697;
22282: douta=16'h8c53;
22283: douta=16'h8c94;
22284: douta=16'h94b6;
22285: douta=16'h7bf2;
22286: douta=16'h8c74;
22287: douta=16'h94b6;
22288: douta=16'h94f7;
22289: douta=16'h31e9;
22290: douta=16'h10c3;
22291: douta=16'h18e4;
22292: douta=16'h18e5;
22293: douta=16'h2168;
22294: douta=16'h1947;
22295: douta=16'h1926;
22296: douta=16'h1105;
22297: douta=16'h1927;
22298: douta=16'h1967;
22299: douta=16'h1947;
22300: douta=16'h1968;
22301: douta=16'h1148;
22302: douta=16'h1947;
22303: douta=16'h2168;
22304: douta=16'h1906;
22305: douta=16'h29ca;
22306: douta=16'h1926;
22307: douta=16'h18e5;
22308: douta=16'h1927;
22309: douta=16'h3a0b;
22310: douta=16'h2148;
22311: douta=16'h2188;
22312: douta=16'h6b2e;
22313: douta=16'h5b30;
22314: douta=16'h42f0;
22315: douta=16'h31c9;
22316: douta=16'h2988;
22317: douta=16'h29a9;
22318: douta=16'h3a0b;
22319: douta=16'h31a9;
22320: douta=16'h39a9;
22321: douta=16'h2967;
22322: douta=16'h31c9;
22323: douta=16'h31c9;
22324: douta=16'h2147;
22325: douta=16'h29ea;
22326: douta=16'h320a;
22327: douta=16'h428c;
22328: douta=16'h4aad;
22329: douta=16'h4acd;
22330: douta=16'h530d;
22331: douta=16'h52ed;
22332: douta=16'h530d;
22333: douta=16'h52cc;
22334: douta=16'h634e;
22335: douta=16'h5b2e;
22336: douta=16'h634e;
22337: douta=16'h5b2d;
22338: douta=16'h5b0d;
22339: douta=16'h5b2d;
22340: douta=16'h52ab;
22341: douta=16'h524a;
22342: douta=16'h5aec;
22343: douta=16'h528a;
22344: douta=16'h528b;
22345: douta=16'h632d;
22346: douta=16'h5acb;
22347: douta=16'h62ec;
22348: douta=16'h5acb;
22349: douta=16'h630c;
22350: douta=16'h62ec;
22351: douta=16'h62cb;
22352: douta=16'h62cb;
22353: douta=16'h6b0c;
22354: douta=16'h6b2c;
22355: douta=16'h734d;
22356: douta=16'h734d;
22357: douta=16'h7bcf;
22358: douta=16'h7baf;
22359: douta=16'h83ef;
22360: douta=16'h7b6d;
22361: douta=16'h83cf;
22362: douta=16'h736d;
22363: douta=16'h83d0;
22364: douta=16'h8431;
22365: douta=16'h83cf;
22366: douta=16'ha534;
22367: douta=16'hb533;
22368: douta=16'hb552;
22369: douta=16'hc4ad;
22370: douta=16'hccaa;
22371: douta=16'hd4aa;
22372: douta=16'hdcc4;
22373: douta=16'hc468;
22374: douta=16'ha42c;
22375: douta=16'h7b8f;
22376: douta=16'h7b6f;
22377: douta=16'h734f;
22378: douta=16'h736d;
22379: douta=16'h7b4d;
22380: douta=16'h93ef;
22381: douta=16'hde76;
22382: douta=16'he697;
22383: douta=16'hd637;
22384: douta=16'h7c33;
22385: douta=16'hbd96;
22386: douta=16'hc595;
22387: douta=16'h94d5;
22388: douta=16'h94d5;
22389: douta=16'h7bf1;
22390: douta=16'h7bd1;
22391: douta=16'h736f;
22392: douta=16'h6b70;
22393: douta=16'h6b4f;
22394: douta=16'h6b2e;
22395: douta=16'h630e;
22396: douta=16'h4a4a;
22397: douta=16'h8bee;
22398: douta=16'hac6e;
22399: douta=16'hde14;
22400: douta=16'he656;
22401: douta=16'he677;
22402: douta=16'he656;
22403: douta=16'hddf5;
22404: douta=16'hbd33;
22405: douta=16'hb555;
22406: douta=16'hbd95;
22407: douta=16'had55;
22408: douta=16'h8c53;
22409: douta=16'h8c74;
22410: douta=16'h7bd1;
22411: douta=16'h7bd0;
22412: douta=16'h7bd1;
22413: douta=16'h6b8f;
22414: douta=16'h7390;
22415: douta=16'h6b4f;
22416: douta=16'h734f;
22417: douta=16'h6b0d;
22418: douta=16'h5acc;
22419: douta=16'h5aed;
22420: douta=16'h524a;
22421: douta=16'h5a8a;
22422: douta=16'h730c;
22423: douta=16'h7b6c;
22424: douta=16'h942e;
22425: douta=16'h9c4f;
22426: douta=16'hb510;
22427: douta=16'hd5d3;
22428: douta=16'hde35;
22429: douta=16'hbd33;
22430: douta=16'hacf4;
22431: douta=16'h8c73;
22432: douta=16'h7c12;
22433: douta=16'h5b30;
22434: douta=16'h42ae;
22435: douta=16'h31eb;
22436: douta=16'h31ea;
22437: douta=16'h426d;
22438: douta=16'h1905;
22439: douta=16'h1906;
22440: douta=16'h2147;
22441: douta=16'h2105;
22442: douta=16'h8286;
22443: douta=16'h6a44;
22444: douta=16'h6a25;
22445: douta=16'h6a04;
22446: douta=16'h6a25;
22447: douta=16'h6205;
22448: douta=16'h61e4;
22449: douta=16'h61e5;
22450: douta=16'h59e5;
22451: douta=16'h59c5;
22452: douta=16'h51a5;
22453: douta=16'h59c5;
22454: douta=16'h51c5;
22455: douta=16'h51c5;
22456: douta=16'h51c5;
22457: douta=16'h51c5;
22458: douta=16'h49a6;
22459: douta=16'h4986;
22460: douta=16'h49a6;
22461: douta=16'h4986;
22462: douta=16'h4165;
22463: douta=16'h41a6;
22464: douta=16'hde32;
22465: douta=16'hd58e;
22466: douta=16'hff5b;
22467: douta=16'hf6f8;
22468: douta=16'hff3a;
22469: douta=16'hff3a;
22470: douta=16'hf719;
22471: douta=16'hff7c;
22472: douta=16'heeb7;
22473: douta=16'hde16;
22474: douta=16'h8c54;
22475: douta=16'h94b5;
22476: douta=16'h8c74;
22477: douta=16'h8412;
22478: douta=16'h8c74;
22479: douta=16'h94b6;
22480: douta=16'h9d17;
22481: douta=16'h1105;
22482: douta=16'h0842;
22483: douta=16'h0882;
22484: douta=16'h10c4;
22485: douta=16'h1905;
22486: douta=16'h1927;
22487: douta=16'h1905;
22488: douta=16'h10e5;
22489: douta=16'h1927;
22490: douta=16'h1948;
22491: douta=16'h1947;
22492: douta=16'h1968;
22493: douta=16'h2168;
22494: douta=16'h2168;
22495: douta=16'h2189;
22496: douta=16'h1927;
22497: douta=16'h2188;
22498: douta=16'h2988;
22499: douta=16'h2147;
22500: douta=16'h10e5;
22501: douta=16'h2988;
22502: douta=16'h31ca;
22503: douta=16'h31c9;
22504: douta=16'h9c31;
22505: douta=16'h73d2;
22506: douta=16'h4332;
22507: douta=16'h2988;
22508: douta=16'h31ca;
22509: douta=16'h2988;
22510: douta=16'h31ca;
22511: douta=16'h2988;
22512: douta=16'h39e9;
22513: douta=16'h2988;
22514: douta=16'h31c9;
22515: douta=16'h2988;
22516: douta=16'h29a9;
22517: douta=16'h3a2b;
22518: douta=16'h3a4b;
22519: douta=16'h4aad;
22520: douta=16'h4aad;
22521: douta=16'h4aac;
22522: douta=16'h52cd;
22523: douta=16'h52ed;
22524: douta=16'h52ed;
22525: douta=16'h52cc;
22526: douta=16'h52ed;
22527: douta=16'h5b0d;
22528: douta=16'h5b2d;
22529: douta=16'h5b2d;
22530: douta=16'h52cc;
22531: douta=16'h5b0d;
22532: douta=16'h62ed;
22533: douta=16'h528b;
22534: douta=16'h5aab;
22535: douta=16'h5acb;
22536: douta=16'h634d;
22537: douta=16'h73af;
22538: douta=16'h62ec;
22539: douta=16'h62eb;
22540: douta=16'h630c;
22541: douta=16'h62ec;
22542: douta=16'h62cb;
22543: douta=16'h732c;
22544: douta=16'h6b0c;
22545: douta=16'h6b0c;
22546: douta=16'h738d;
22547: douta=16'h736e;
22548: douta=16'h7b8e;
22549: douta=16'h8c31;
22550: douta=16'h8410;
22551: douta=16'h7bcf;
22552: douta=16'h83f0;
22553: douta=16'h7bef;
22554: douta=16'h8c51;
22555: douta=16'had55;
22556: douta=16'hc638;
22557: douta=16'hce38;
22558: douta=16'hcd0c;
22559: douta=16'hd4ea;
22560: douta=16'hd4a7;
22561: douta=16'hdc85;
22562: douta=16'hcc23;
22563: douta=16'hcc44;
22564: douta=16'hcc46;
22565: douta=16'hdc84;
22566: douta=16'hdc84;
22567: douta=16'hbc4b;
22568: douta=16'hb42a;
22569: douta=16'hb42c;
22570: douta=16'hcdd5;
22571: douta=16'hd5d4;
22572: douta=16'he677;
22573: douta=16'hde16;
22574: douta=16'hd5f6;
22575: douta=16'hc5d7;
22576: douta=16'h7c33;
22577: douta=16'hbd96;
22578: douta=16'hc5b6;
22579: douta=16'h9495;
22580: douta=16'h8c53;
22581: douta=16'h7bd1;
22582: douta=16'h7bb0;
22583: douta=16'h736f;
22584: douta=16'h7390;
22585: douta=16'h62cd;
22586: douta=16'h52ad;
22587: douta=16'h52ad;
22588: douta=16'hb4d1;
22589: douta=16'he634;
22590: douta=16'hd5f4;
22591: douta=16'he656;
22592: douta=16'he656;
22593: douta=16'he656;
22594: douta=16'hd5f6;
22595: douta=16'hd5d5;
22596: douta=16'hcdb4;
22597: douta=16'had14;
22598: douta=16'hb556;
22599: douta=16'hb556;
22600: douta=16'h8452;
22601: douta=16'h8433;
22602: douta=16'h8412;
22603: douta=16'h7bb0;
22604: douta=16'h7391;
22605: douta=16'h73b0;
22606: douta=16'h73b0;
22607: douta=16'h6b4f;
22608: douta=16'h5acd;
22609: douta=16'h736f;
22610: douta=16'h6b2e;
22611: douta=16'h6b2d;
22612: douta=16'h3965;
22613: douta=16'h5a47;
22614: douta=16'h9c4e;
22615: douta=16'hbd51;
22616: douta=16'hcdb2;
22617: douta=16'hd5b3;
22618: douta=16'hd5f3;
22619: douta=16'hde34;
22620: douta=16'hde15;
22621: douta=16'hb534;
22622: douta=16'hacf4;
22623: douta=16'h8c73;
22624: douta=16'h7c33;
22625: douta=16'h5b50;
22626: douta=16'h5310;
22627: douta=16'h3a4c;
22628: douta=16'h320b;
22629: douta=16'h2168;
22630: douta=16'h10c5;
22631: douta=16'h2127;
22632: douta=16'h1926;
22633: douta=16'h00a5;
22634: douta=16'h82a5;
22635: douta=16'h7244;
22636: douta=16'h7225;
22637: douta=16'h6a24;
22638: douta=16'h6a04;
22639: douta=16'h6205;
22640: douta=16'h61e4;
22641: douta=16'h6205;
22642: douta=16'h59e5;
22643: douta=16'h59c5;
22644: douta=16'h59c5;
22645: douta=16'h59c5;
22646: douta=16'h51c5;
22647: douta=16'h51c6;
22648: douta=16'h51c5;
22649: douta=16'h51c6;
22650: douta=16'h49a6;
22651: douta=16'h49a6;
22652: douta=16'h4986;
22653: douta=16'h49a5;
22654: douta=16'h4165;
22655: douta=16'h4165;
22656: douta=16'heeb6;
22657: douta=16'hf6d8;
22658: douta=16'hf719;
22659: douta=16'hfef9;
22660: douta=16'hff19;
22661: douta=16'hf719;
22662: douta=16'hf719;
22663: douta=16'hff9b;
22664: douta=16'hd5d6;
22665: douta=16'hb535;
22666: douta=16'h9cf6;
22667: douta=16'h9cd5;
22668: douta=16'h94d5;
22669: douta=16'h9c94;
22670: douta=16'h94d5;
22671: douta=16'h94d6;
22672: douta=16'h8c75;
22673: douta=16'h5b72;
22674: douta=16'h7415;
22675: douta=16'h84d8;
22676: douta=16'h8d3a;
22677: douta=16'h21a8;
22678: douta=16'h10a3;
22679: douta=16'h10e5;
22680: douta=16'h10e4;
22681: douta=16'h1127;
22682: douta=16'h1927;
22683: douta=16'h1947;
22684: douta=16'h2169;
22685: douta=16'h1968;
22686: douta=16'h2188;
22687: douta=16'h1947;
22688: douta=16'h1946;
22689: douta=16'h1947;
22690: douta=16'h2168;
22691: douta=16'h29a9;
22692: douta=16'h2189;
22693: douta=16'h29a9;
22694: douta=16'h29a9;
22695: douta=16'h2187;
22696: douta=16'h2126;
22697: douta=16'h1906;
22698: douta=16'h1906;
22699: douta=16'h2168;
22700: douta=16'h2167;
22701: douta=16'h2167;
22702: douta=16'h2126;
22703: douta=16'h2106;
22704: douta=16'h1082;
22705: douta=16'h31c9;
22706: douta=16'h31c9;
22707: douta=16'h2106;
22708: douta=16'h31ea;
22709: douta=16'h31e9;
22710: douta=16'h3a0a;
22711: douta=16'h424b;
22712: douta=16'h428c;
22713: douta=16'h4aad;
22714: douta=16'h424a;
22715: douta=16'h4aac;
22716: douta=16'h4a8c;
22717: douta=16'h4aac;
22718: douta=16'h52ac;
22719: douta=16'h4a8b;
22720: douta=16'h4249;
22721: douta=16'h4249;
22722: douta=16'h4a4a;
22723: douta=16'h5b0d;
22724: douta=16'h52cb;
22725: douta=16'h52cc;
22726: douta=16'h5269;
22727: douta=16'h5acb;
22728: douta=16'h5aaa;
22729: douta=16'h738f;
22730: douta=16'h6b8e;
22731: douta=16'h6b0c;
22732: douta=16'h736e;
22733: douta=16'h62ec;
22734: douta=16'h6b2d;
22735: douta=16'h7bf1;
22736: douta=16'h73b0;
22737: douta=16'h83cf;
22738: douta=16'hb553;
22739: douta=16'hd615;
22740: douta=16'he6b8;
22741: douta=16'he5d0;
22742: douta=16'he56d;
22743: douta=16'hcc24;
22744: douta=16'hc3c2;
22745: douta=16'hc3c2;
22746: douta=16'hc3c2;
22747: douta=16'hcc25;
22748: douta=16'hcc25;
22749: douta=16'hcc25;
22750: douta=16'hcc25;
22751: douta=16'hcc25;
22752: douta=16'hcc66;
22753: douta=16'hcc66;
22754: douta=16'hd466;
22755: douta=16'hcc45;
22756: douta=16'hcc66;
22757: douta=16'hcc66;
22758: douta=16'hcc66;
22759: douta=16'hd466;
22760: douta=16'hcc66;
22761: douta=16'hd466;
22762: douta=16'hd466;
22763: douta=16'hc447;
22764: douta=16'hb4b2;
22765: douta=16'ha4f4;
22766: douta=16'ha4d4;
22767: douta=16'ha4d5;
22768: douta=16'h8c53;
22769: douta=16'hb576;
22770: douta=16'hc5d7;
22771: douta=16'h8453;
22772: douta=16'h7bd1;
22773: douta=16'h7bb1;
22774: douta=16'h7bb0;
22775: douta=16'h736f;
22776: douta=16'h52ac;
22777: douta=16'h9410;
22778: douta=16'hd5d4;
22779: douta=16'h8bee;
22780: douta=16'hde15;
22781: douta=16'hddf5;
22782: douta=16'hde15;
22783: douta=16'hd5f5;
22784: douta=16'hcdb4;
22785: douta=16'hbd56;
22786: douta=16'ha4d6;
22787: douta=16'h9c95;
22788: douta=16'h9cd5;
22789: douta=16'ha4d5;
22790: douta=16'hacf5;
22791: douta=16'h9494;
22792: douta=16'h8432;
22793: douta=16'h6b70;
22794: douta=16'h62ed;
22795: douta=16'h6b6f;
22796: douta=16'h6b4f;
22797: douta=16'h7bf1;
22798: douta=16'h5b0e;
22799: douta=16'h630d;
22800: douta=16'h41e8;
22801: douta=16'h3985;
22802: douta=16'h62c9;
22803: douta=16'h732a;
22804: douta=16'h942d;
22805: douta=16'ha4af;
22806: douta=16'ha4ef;
22807: douta=16'h9c2e;
22808: douta=16'hbd4f;
22809: douta=16'hcdb2;
22810: douta=16'hde15;
22811: douta=16'hd614;
22812: douta=16'hc554;
22813: douta=16'had15;
22814: douta=16'ha4f5;
22815: douta=16'h94d5;
22816: douta=16'h7c34;
22817: douta=16'h6bf2;
22818: douta=16'h5b50;
22819: douta=16'h4aae;
22820: douta=16'h428e;
22821: douta=16'h3a4d;
22822: douta=16'h532f;
22823: douta=16'h2147;
22824: douta=16'h1905;
22825: douta=16'h18e5;
22826: douta=16'h00a5;
22827: douta=16'h8286;
22828: douta=16'h7225;
22829: douta=16'h7225;
22830: douta=16'h6a04;
22831: douta=16'h6205;
22832: douta=16'h61e5;
22833: douta=16'h61e5;
22834: douta=16'h59e5;
22835: douta=16'h59c5;
22836: douta=16'h59c5;
22837: douta=16'h59e6;
22838: douta=16'h51e5;
22839: douta=16'h51c6;
22840: douta=16'h51c6;
22841: douta=16'h49c6;
22842: douta=16'h49a6;
22843: douta=16'h49a6;
22844: douta=16'h4985;
22845: douta=16'h4186;
22846: douta=16'h4185;
22847: douta=16'h4165;
22848: douta=16'hf6d7;
22849: douta=16'hff1a;
22850: douta=16'hf6f9;
22851: douta=16'hf73a;
22852: douta=16'hff19;
22853: douta=16'hf6f9;
22854: douta=16'hff3a;
22855: douta=16'hf6d8;
22856: douta=16'hc5b6;
22857: douta=16'had16;
22858: douta=16'h9cf6;
22859: douta=16'h94b5;
22860: douta=16'h9cb5;
22861: douta=16'h9c94;
22862: douta=16'ha517;
22863: douta=16'h9cf6;
22864: douta=16'h6c14;
22865: douta=16'h7435;
22866: douta=16'h7456;
22867: douta=16'h7c77;
22868: douta=16'h8497;
22869: douta=16'h84b8;
22870: douta=16'h0001;
22871: douta=16'h1105;
22872: douta=16'h10e5;
22873: douta=16'h1947;
22874: douta=16'h1947;
22875: douta=16'h1127;
22876: douta=16'h1967;
22877: douta=16'h1927;
22878: douta=16'h1926;
22879: douta=16'h1948;
22880: douta=16'h1926;
22881: douta=16'h2167;
22882: douta=16'h18e5;
22883: douta=16'h1082;
22884: douta=16'h2188;
22885: douta=16'h2168;
22886: douta=16'h2168;
22887: douta=16'h2146;
22888: douta=16'h2126;
22889: douta=16'h18e4;
22890: douta=16'h29c9;
22891: douta=16'h3a2b;
22892: douta=16'h18a1;
22893: douta=16'h3144;
22894: douta=16'h0800;
22895: douta=16'h0821;
22896: douta=16'h0820;
22897: douta=16'h2126;
22898: douta=16'h1905;
22899: douta=16'h29c8;
22900: douta=16'h31e9;
22901: douta=16'h3a0a;
22902: douta=16'h3a2b;
22903: douta=16'h31e9;
22904: douta=16'h31e9;
22905: douta=16'h31c9;
22906: douta=16'h39e9;
22907: douta=16'h39c8;
22908: douta=16'h4229;
22909: douta=16'h4229;
22910: douta=16'h3a09;
22911: douta=16'h4a8b;
22912: douta=16'h4a4a;
22913: douta=16'h4a4a;
22914: douta=16'h526b;
22915: douta=16'h5acc;
22916: douta=16'h638e;
22917: douta=16'h6baf;
22918: douta=16'h73f1;
22919: douta=16'h8473;
22920: douta=16'h73f1;
22921: douta=16'h5aed;
22922: douta=16'h6b8f;
22923: douta=16'h7b6d;
22924: douta=16'hac4e;
22925: douta=16'hcd70;
22926: douta=16'hc50e;
22927: douta=16'hcc24;
22928: douta=16'hcbe3;
22929: douta=16'hc403;
22930: douta=16'hbba3;
22931: douta=16'hc3e2;
22932: douta=16'hc3e2;
22933: douta=16'hcc25;
22934: douta=16'hcc25;
22935: douta=16'hcc25;
22936: douta=16'hcc25;
22937: douta=16'hcc45;
22938: douta=16'hcc45;
22939: douta=16'hcc45;
22940: douta=16'hcc45;
22941: douta=16'hcc45;
22942: douta=16'hcc45;
22943: douta=16'hcc46;
22944: douta=16'hcc45;
22945: douta=16'hcc45;
22946: douta=16'hcc46;
22947: douta=16'hcc45;
22948: douta=16'hd465;
22949: douta=16'hd466;
22950: douta=16'hcc66;
22951: douta=16'hd466;
22952: douta=16'hd466;
22953: douta=16'hcc66;
22954: douta=16'hcc66;
22955: douta=16'hd486;
22956: douta=16'hd444;
22957: douta=16'h9c53;
22958: douta=16'h9c51;
22959: douta=16'h9c72;
22960: douta=16'h9452;
22961: douta=16'ha4f5;
22962: douta=16'ha516;
22963: douta=16'h8412;
22964: douta=16'h73d0;
22965: douta=16'h736f;
22966: douta=16'h4a6b;
22967: douta=16'h732e;
22968: douta=16'hb4b0;
22969: douta=16'hde36;
22970: douta=16'hbd52;
22971: douta=16'hde96;
22972: douta=16'hd5b4;
22973: douta=16'hde15;
22974: douta=16'hde15;
22975: douta=16'hbd34;
22976: douta=16'hb535;
22977: douta=16'h9c94;
22978: douta=16'h9494;
22979: douta=16'h8412;
22980: douta=16'h83f1;
22981: douta=16'h8453;
22982: douta=16'h9494;
22983: douta=16'ha4f6;
22984: douta=16'h73d1;
22985: douta=16'h630e;
22986: douta=16'h5aee;
22987: douta=16'h632f;
22988: douta=16'h632f;
22989: douta=16'h524a;
22990: douta=16'h3985;
22991: douta=16'h5228;
22992: douta=16'h93ed;
22993: douta=16'hc551;
22994: douta=16'hc550;
22995: douta=16'hd5b1;
22996: douta=16'hde35;
22997: douta=16'he676;
22998: douta=16'he656;
22999: douta=16'he696;
23000: douta=16'he656;
23001: douta=16'hde35;
23002: douta=16'he655;
23003: douta=16'hcdb5;
23004: douta=16'had16;
23005: douta=16'h9cf5;
23006: douta=16'h94d5;
23007: douta=16'h94d6;
23008: douta=16'h7c34;
23009: douta=16'h6bf3;
23010: douta=16'h7414;
23011: douta=16'h5330;
23012: douta=16'h4b10;
23013: douta=16'h5331;
23014: douta=16'h52ef;
23015: douta=16'h1106;
23016: douta=16'h2168;
23017: douta=16'h2127;
23018: douta=16'h10c6;
23019: douta=16'h8a85;
23020: douta=16'h6a24;
23021: douta=16'h6a24;
23022: douta=16'h6a05;
23023: douta=16'h61e5;
23024: douta=16'h6205;
23025: douta=16'h61e5;
23026: douta=16'h59c5;
23027: douta=16'h59c5;
23028: douta=16'h59c5;
23029: douta=16'h59c6;
23030: douta=16'h51c6;
23031: douta=16'h51c6;
23032: douta=16'h49c6;
23033: douta=16'h49c6;
23034: douta=16'h49a5;
23035: douta=16'h49a6;
23036: douta=16'h4985;
23037: douta=16'h4185;
23038: douta=16'h4185;
23039: douta=16'h4165;
23040: douta=16'heed7;
23041: douta=16'hf71a;
23042: douta=16'hf6f9;
23043: douta=16'hf73a;
23044: douta=16'hf6f9;
23045: douta=16'hff19;
23046: douta=16'hff3a;
23047: douta=16'hee97;
23048: douta=16'hbd96;
23049: douta=16'had16;
23050: douta=16'ha516;
23051: douta=16'h94d5;
23052: douta=16'h9c94;
23053: douta=16'h9cb4;
23054: douta=16'h9cd6;
23055: douta=16'ha516;
23056: douta=16'h7455;
23057: douta=16'h7c97;
23058: douta=16'h7cb7;
23059: douta=16'h7c76;
23060: douta=16'h7c96;
23061: douta=16'h7c76;
23062: douta=16'h3a6c;
23063: douta=16'h0042;
23064: douta=16'h1083;
23065: douta=16'h1947;
23066: douta=16'h1927;
23067: douta=16'h1927;
23068: douta=16'h1906;
23069: douta=16'h1105;
23070: douta=16'h1105;
23071: douta=16'h1947;
23072: douta=16'h2189;
23073: douta=16'h21a9;
23074: douta=16'h2168;
23075: douta=16'h1927;
23076: douta=16'h10e4;
23077: douta=16'h2189;
23078: douta=16'h2188;
23079: douta=16'h2168;
23080: douta=16'h2146;
23081: douta=16'h10c5;
23082: douta=16'h29a8;
23083: douta=16'h29ca;
23084: douta=16'h1061;
23085: douta=16'h18a2;
23086: douta=16'h0000;
23087: douta=16'h2924;
23088: douta=16'h1882;
23089: douta=16'h2967;
23090: douta=16'h31c9;
23091: douta=16'h29c9;
23092: douta=16'h3a2b;
23093: douta=16'h31c9;
23094: douta=16'h3a0a;
23095: douta=16'h39c9;
23096: douta=16'h31a8;
23097: douta=16'h39e9;
23098: douta=16'h39e8;
23099: douta=16'h39c9;
23100: douta=16'h39e9;
23101: douta=16'h424a;
23102: douta=16'h4a6b;
23103: douta=16'h52ac;
23104: douta=16'h4aab;
23105: douta=16'h52ab;
23106: douta=16'h528b;
23107: douta=16'h634e;
23108: douta=16'h636f;
23109: douta=16'h6b90;
23110: douta=16'h6b4e;
23111: douta=16'h738f;
23112: douta=16'h834b;
23113: douta=16'h8b27;
23114: douta=16'h9b47;
23115: douta=16'hb3a5;
23116: douta=16'hc3e5;
23117: douta=16'hc3e3;
23118: douta=16'hbb83;
23119: douta=16'hbbe4;
23120: douta=16'hbbe5;
23121: douta=16'hc3e5;
23122: douta=16'hc403;
23123: douta=16'hc406;
23124: douta=16'hcc25;
23125: douta=16'hc425;
23126: douta=16'hcc25;
23127: douta=16'hcc25;
23128: douta=16'hc425;
23129: douta=16'hc425;
23130: douta=16'hcc45;
23131: douta=16'hcc45;
23132: douta=16'hcc45;
23133: douta=16'hcc25;
23134: douta=16'hcc45;
23135: douta=16'hcc66;
23136: douta=16'hcc45;
23137: douta=16'hd445;
23138: douta=16'hcc66;
23139: douta=16'hcc66;
23140: douta=16'hcc66;
23141: douta=16'hd465;
23142: douta=16'hcc66;
23143: douta=16'hd466;
23144: douta=16'hcc66;
23145: douta=16'hd466;
23146: douta=16'hcc65;
23147: douta=16'hcc66;
23148: douta=16'hd466;
23149: douta=16'ha42d;
23150: douta=16'h9410;
23151: douta=16'h9430;
23152: douta=16'h9430;
23153: douta=16'h9cb3;
23154: douta=16'h9453;
23155: douta=16'h83d0;
23156: douta=16'h7bb0;
23157: douta=16'h632f;
23158: douta=16'hacb0;
23159: douta=16'he675;
23160: douta=16'h93cd;
23161: douta=16'hb555;
23162: douta=16'hc574;
23163: douta=16'he677;
23164: douta=16'hc554;
23165: douta=16'hd5d6;
23166: douta=16'hc595;
23167: douta=16'hbd34;
23168: douta=16'hb515;
23169: douta=16'h9cb4;
23170: douta=16'h8c73;
23171: douta=16'h7bf2;
23172: douta=16'h73b1;
23173: douta=16'h7bf1;
23174: douta=16'h8432;
23175: douta=16'h8c73;
23176: douta=16'h7390;
23177: douta=16'h7370;
23178: douta=16'h6b50;
23179: douta=16'h632f;
23180: douta=16'h41e7;
23181: douta=16'h4a08;
23182: douta=16'h734b;
23183: douta=16'h83ac;
23184: douta=16'h93ed;
23185: douta=16'hcd72;
23186: douta=16'hde34;
23187: douta=16'hde14;
23188: douta=16'he656;
23189: douta=16'hde55;
23190: douta=16'he656;
23191: douta=16'hd5f4;
23192: douta=16'hd5f4;
23193: douta=16'hd5f4;
23194: douta=16'hcd93;
23195: douta=16'hb535;
23196: douta=16'ha516;
23197: douta=16'h94d5;
23198: douta=16'h94d5;
23199: douta=16'h8cb5;
23200: douta=16'h7c54;
23201: douta=16'h7413;
23202: douta=16'h7413;
23203: douta=16'h5330;
23204: douta=16'h5330;
23205: douta=16'h5b72;
23206: douta=16'h324b;
23207: douta=16'h4a8c;
23208: douta=16'h2968;
23209: douta=16'h2127;
23210: douta=16'h1927;
23211: douta=16'h7a65;
23212: douta=16'h7245;
23213: douta=16'h6a25;
23214: douta=16'h6a25;
23215: douta=16'h6205;
23216: douta=16'h61e5;
23217: douta=16'h61e5;
23218: douta=16'h59c5;
23219: douta=16'h59e5;
23220: douta=16'h59e5;
23221: douta=16'h51c5;
23222: douta=16'h51c6;
23223: douta=16'h51c5;
23224: douta=16'h49c6;
23225: douta=16'h49a5;
23226: douta=16'h49a6;
23227: douta=16'h49a6;
23228: douta=16'h49a6;
23229: douta=16'h4185;
23230: douta=16'h4185;
23231: douta=16'h4186;
23232: douta=16'hf6f8;
23233: douta=16'hf6f8;
23234: douta=16'hf719;
23235: douta=16'hff19;
23236: douta=16'hff19;
23237: douta=16'hff19;
23238: douta=16'hff7b;
23239: douta=16'hd5d5;
23240: douta=16'had16;
23241: douta=16'h9cb4;
23242: douta=16'h9cd5;
23243: douta=16'ha516;
23244: douta=16'h9cb4;
23245: douta=16'h9cf5;
23246: douta=16'ha516;
23247: douta=16'ha516;
23248: douta=16'h6bf3;
23249: douta=16'h7414;
23250: douta=16'h73f4;
23251: douta=16'h7c76;
23252: douta=16'h8497;
23253: douta=16'h7c76;
23254: douta=16'h8476;
23255: douta=16'h7c76;
23256: douta=16'h8497;
23257: douta=16'h0884;
23258: douta=16'h10c5;
23259: douta=16'h10c5;
23260: douta=16'h1105;
23261: douta=16'h1105;
23262: douta=16'h08c5;
23263: douta=16'h10e5;
23264: douta=16'h1906;
23265: douta=16'h1926;
23266: douta=16'h1926;
23267: douta=16'h1927;
23268: douta=16'h2147;
23269: douta=16'h18e5;
23270: douta=16'h10c4;
23271: douta=16'h18c4;
23272: douta=16'h2126;
23273: douta=16'h10c5;
23274: douta=16'h2126;
23275: douta=16'h2146;
23276: douta=16'h2147;
23277: douta=16'h20e5;
23278: douta=16'h1083;
23279: douta=16'h2145;
23280: douta=16'h320b;
23281: douta=16'h3a2c;
23282: douta=16'h3a2c;
23283: douta=16'h320a;
23284: douta=16'h3a2b;
23285: douta=16'h4aad;
23286: douta=16'h4ace;
23287: douta=16'h4ace;
23288: douta=16'h426c;
23289: douta=16'h3a2a;
23290: douta=16'h3a2b;
23291: douta=16'h4a8c;
23292: douta=16'h4aac;
23293: douta=16'h62cb;
23294: douta=16'h6aea;
23295: douta=16'h6267;
23296: douta=16'h8263;
23297: douta=16'h8283;
23298: douta=16'h8aa2;
23299: douta=16'h9ac2;
23300: douta=16'ha325;
23301: douta=16'ha345;
23302: douta=16'hab84;
23303: douta=16'hab64;
23304: douta=16'hb365;
23305: douta=16'hb3a5;
23306: douta=16'hb3a5;
23307: douta=16'hb3c5;
23308: douta=16'hb3c4;
23309: douta=16'hbbe5;
23310: douta=16'hbbc6;
23311: douta=16'hbbe5;
23312: douta=16'hc3e5;
23313: douta=16'hc405;
23314: douta=16'hc425;
23315: douta=16'hcc05;
23316: douta=16'hc406;
23317: douta=16'hcc25;
23318: douta=16'hcc46;
23319: douta=16'hcc47;
23320: douta=16'hcc46;
23321: douta=16'hcc66;
23322: douta=16'hcc25;
23323: douta=16'hcc25;
23324: douta=16'hcc46;
23325: douta=16'hcc45;
23326: douta=16'hcc45;
23327: douta=16'hcc46;
23328: douta=16'hcc44;
23329: douta=16'hcc45;
23330: douta=16'hcc24;
23331: douta=16'hcc02;
23332: douta=16'hcc00;
23333: douta=16'hcc44;
23334: douta=16'hcc87;
23335: douta=16'hd56e;
23336: douta=16'he5d0;
23337: douta=16'he694;
23338: douta=16'hf77a;
23339: douta=16'hffbc;
23340: douta=16'hf7dc;
23341: douta=16'hf6f6;
23342: douta=16'he693;
23343: douta=16'hf650;
23344: douta=16'hbc29;
23345: douta=16'ha3ca;
23346: douta=16'hac6f;
23347: douta=16'hd5d4;
23348: douta=16'hde14;
23349: douta=16'he656;
23350: douta=16'hde36;
23351: douta=16'hd5f5;
23352: douta=16'heeb7;
23353: douta=16'hbd76;
23354: douta=16'hc5d7;
23355: douta=16'hcdd7;
23356: douta=16'h8c96;
23357: douta=16'h8454;
23358: douta=16'h94b5;
23359: douta=16'h8453;
23360: douta=16'h8c53;
23361: douta=16'h8412;
23362: douta=16'h8412;
23363: douta=16'h6b6f;
23364: douta=16'h6b6f;
23365: douta=16'h6b2f;
23366: douta=16'h73b0;
23367: douta=16'h6b70;
23368: douta=16'h524a;
23369: douta=16'h41c6;
23370: douta=16'h5228;
23371: douta=16'h9c4e;
23372: douta=16'hc530;
23373: douta=16'hcd91;
23374: douta=16'hd5f4;
23375: douta=16'he655;
23376: douta=16'hc533;
23377: douta=16'hcd93;
23378: douta=16'hd5b3;
23379: douta=16'hd5d4;
23380: douta=16'hd5b3;
23381: douta=16'hd5b4;
23382: douta=16'hbd34;
23383: douta=16'hbd75;
23384: douta=16'h9cb3;
23385: douta=16'h9cb3;
23386: douta=16'h9cd5;
23387: douta=16'h9cf5;
23388: douta=16'h9d16;
23389: douta=16'h8cb5;
23390: douta=16'h8cd5;
23391: douta=16'h8c95;
23392: douta=16'h7c54;
23393: douta=16'h7434;
23394: douta=16'h7434;
23395: douta=16'h7c75;
23396: douta=16'h7414;
23397: douta=16'h63b2;
23398: douta=16'h52ef;
23399: douta=16'h31a7;
23400: douta=16'h7b90;
23401: douta=16'h2127;
23402: douta=16'h1926;
23403: douta=16'h08c5;
23404: douta=16'h7245;
23405: douta=16'h6a25;
23406: douta=16'h6a25;
23407: douta=16'h61e5;
23408: douta=16'h59e5;
23409: douta=16'h61e5;
23410: douta=16'h59e5;
23411: douta=16'h59e5;
23412: douta=16'h59c5;
23413: douta=16'h51c5;
23414: douta=16'h51c5;
23415: douta=16'h51c5;
23416: douta=16'h51c5;
23417: douta=16'h49a5;
23418: douta=16'h49a6;
23419: douta=16'h4986;
23420: douta=16'h49a6;
23421: douta=16'h4185;
23422: douta=16'h4186;
23423: douta=16'h3966;
23424: douta=16'hff19;
23425: douta=16'hf6d8;
23426: douta=16'hff19;
23427: douta=16'hff19;
23428: douta=16'hf719;
23429: douta=16'hff19;
23430: douta=16'hff9b;
23431: douta=16'hcdb6;
23432: douta=16'ha4d5;
23433: douta=16'h9473;
23434: douta=16'ha516;
23435: douta=16'ha4f5;
23436: douta=16'ha4d4;
23437: douta=16'h9cf5;
23438: douta=16'h9cd5;
23439: douta=16'h8c95;
23440: douta=16'h7414;
23441: douta=16'h7434;
23442: douta=16'h7c55;
23443: douta=16'h7c35;
23444: douta=16'h7c76;
23445: douta=16'h84d7;
23446: douta=16'h7c76;
23447: douta=16'h73f3;
23448: douta=16'h6bf4;
23449: douta=16'h0883;
23450: douta=16'h10c5;
23451: douta=16'h08a5;
23452: douta=16'h10e5;
23453: douta=16'h10e5;
23454: douta=16'h10c5;
23455: douta=16'h10e5;
23456: douta=16'h10e5;
23457: douta=16'h10c5;
23458: douta=16'h1105;
23459: douta=16'h1906;
23460: douta=16'h1905;
23461: douta=16'h18e5;
23462: douta=16'h18e5;
23463: douta=16'h2125;
23464: douta=16'h2106;
23465: douta=16'h10e4;
23466: douta=16'h18e5;
23467: douta=16'h18e5;
23468: douta=16'h2125;
23469: douta=16'h2167;
23470: douta=16'h18e4;
23471: douta=16'h31ea;
23472: douta=16'h324c;
23473: douta=16'h3a6c;
23474: douta=16'h3a2c;
23475: douta=16'h3a6c;
23476: douta=16'h3a4c;
23477: douta=16'h42ce;
23478: douta=16'h42ad;
23479: douta=16'h51a5;
23480: douta=16'h51a5;
23481: douta=16'h59e4;
23482: douta=16'h61a3;
23483: douta=16'h69e3;
23484: douta=16'h7203;
23485: douta=16'h7a44;
23486: douta=16'h8aa4;
23487: douta=16'h8ac4;
23488: douta=16'h92e4;
23489: douta=16'h92e4;
23490: douta=16'h9b04;
23491: douta=16'h9b04;
23492: douta=16'ha345;
23493: douta=16'ha344;
23494: douta=16'hab64;
23495: douta=16'hab85;
23496: douta=16'hb385;
23497: douta=16'hab84;
23498: douta=16'hb384;
23499: douta=16'hb3a5;
23500: douta=16'hbbc5;
23501: douta=16'hbbc5;
23502: douta=16'hbbc6;
23503: douta=16'hc3e5;
23504: douta=16'hc3e5;
23505: douta=16'hc405;
23506: douta=16'hc426;
23507: douta=16'hc426;
23508: douta=16'hcc46;
23509: douta=16'hcc46;
23510: douta=16'hcc25;
23511: douta=16'hcc25;
23512: douta=16'hcc25;
23513: douta=16'hcc25;
23514: douta=16'hcc25;
23515: douta=16'hcc04;
23516: douta=16'hc3e2;
23517: douta=16'hc3e1;
23518: douta=16'hcc66;
23519: douta=16'hcca8;
23520: douta=16'hdd6e;
23521: douta=16'he633;
23522: douta=16'heed7;
23523: douta=16'hef39;
23524: douta=16'hffdc;
23525: douta=16'hf7bb;
23526: douta=16'hf738;
23527: douta=16'he611;
23528: douta=16'hddaf;
23529: douta=16'hd50a;
23530: douta=16'hcc65;
23531: douta=16'hcc22;
23532: douta=16'hcc02;
23533: douta=16'hcc45;
23534: douta=16'hd466;
23535: douta=16'hd467;
23536: douta=16'hd486;
23537: douta=16'hd466;
23538: douta=16'hd443;
23539: douta=16'hd5d6;
23540: douta=16'hd5d5;
23541: douta=16'hd5f5;
23542: douta=16'hde56;
23543: douta=16'hde35;
23544: douta=16'hbd97;
23545: douta=16'had77;
23546: douta=16'hbd98;
23547: douta=16'hb598;
23548: douta=16'h8453;
23549: douta=16'h7bf2;
23550: douta=16'h73b1;
23551: douta=16'h73d0;
23552: douta=16'h7b90;
23553: douta=16'h6b6f;
23554: douta=16'h734e;
23555: douta=16'h630e;
23556: douta=16'h632e;
23557: douta=16'h630e;
23558: douta=16'h4a49;
23559: douta=16'h49c6;
23560: douta=16'h7bad;
23561: douta=16'hc571;
23562: douta=16'hc571;
23563: douta=16'hde14;
23564: douta=16'hde56;
23565: douta=16'he656;
23566: douta=16'hde36;
23567: douta=16'hde55;
23568: douta=16'hcdd4;
23569: douta=16'hde36;
23570: douta=16'hde56;
23571: douta=16'hcdd4;
23572: douta=16'hb514;
23573: douta=16'hbd14;
23574: douta=16'h9493;
23575: douta=16'h9c94;
23576: douta=16'h8c93;
23577: douta=16'h94b4;
23578: douta=16'h9493;
23579: douta=16'h7c32;
23580: douta=16'h7c33;
23581: douta=16'h7c33;
23582: douta=16'h7c33;
23583: douta=16'h8454;
23584: douta=16'h73f2;
23585: douta=16'h6bf2;
23586: douta=16'h6bf2;
23587: douta=16'h6bf2;
23588: douta=16'h6b91;
23589: douta=16'h3165;
23590: douta=16'h52cd;
23591: douta=16'h428d;
23592: douta=16'h29a9;
23593: douta=16'h10c5;
23594: douta=16'h10e5;
23595: douta=16'h18e5;
23596: douta=16'h8a85;
23597: douta=16'h7245;
23598: douta=16'h6225;
23599: douta=16'h6a05;
23600: douta=16'h6205;
23601: douta=16'h6205;
23602: douta=16'h59e5;
23603: douta=16'h5a05;
23604: douta=16'h59c5;
23605: douta=16'h51c5;
23606: douta=16'h51c6;
23607: douta=16'h51c6;
23608: douta=16'h49a6;
23609: douta=16'h49a6;
23610: douta=16'h49a6;
23611: douta=16'h49a6;
23612: douta=16'h4185;
23613: douta=16'h41a6;
23614: douta=16'h4166;
23615: douta=16'h4166;
23616: douta=16'hf719;
23617: douta=16'hf6d8;
23618: douta=16'hff19;
23619: douta=16'hf6f8;
23620: douta=16'hf73a;
23621: douta=16'hf719;
23622: douta=16'hef18;
23623: douta=16'hc575;
23624: douta=16'h9c94;
23625: douta=16'h9c93;
23626: douta=16'ha4f5;
23627: douta=16'ha4d5;
23628: douta=16'ha4f5;
23629: douta=16'h9cf5;
23630: douta=16'h9cd5;
23631: douta=16'h7c54;
23632: douta=16'h7c34;
23633: douta=16'h7414;
23634: douta=16'h7c35;
23635: douta=16'h8496;
23636: douta=16'h7c35;
23637: douta=16'h8cd7;
23638: douta=16'h7c75;
23639: douta=16'h7c55;
23640: douta=16'h8476;
23641: douta=16'h10c4;
23642: douta=16'h10e5;
23643: douta=16'h10c4;
23644: douta=16'h10c5;
23645: douta=16'h1106;
23646: douta=16'h1106;
23647: douta=16'h1106;
23648: douta=16'h10e5;
23649: douta=16'h10c5;
23650: douta=16'h1906;
23651: douta=16'h10a4;
23652: douta=16'h10e4;
23653: douta=16'h1905;
23654: douta=16'h18c4;
23655: douta=16'h1905;
23656: douta=16'h1906;
23657: douta=16'h18e5;
23658: douta=16'h1906;
23659: douta=16'h2167;
23660: douta=16'h1926;
23661: douta=16'h2988;
23662: douta=16'h1905;
23663: douta=16'h322b;
23664: douta=16'h3a6c;
23665: douta=16'h3a8e;
23666: douta=16'h430f;
23667: douta=16'h3a4c;
23668: douta=16'h4a4b;
23669: douta=16'h4a07;
23670: douta=16'h51e6;
23671: douta=16'h61e3;
23672: douta=16'h61e3;
23673: douta=16'h59a2;
23674: douta=16'h69e3;
23675: douta=16'h7a44;
23676: douta=16'h7a64;
23677: douta=16'h8284;
23678: douta=16'h8aa4;
23679: douta=16'h8aa3;
23680: douta=16'h92e4;
23681: douta=16'h92e4;
23682: douta=16'h9b04;
23683: douta=16'h9b05;
23684: douta=16'ha345;
23685: douta=16'ha345;
23686: douta=16'hab64;
23687: douta=16'hab64;
23688: douta=16'hb385;
23689: douta=16'hb3a4;
23690: douta=16'hb385;
23691: douta=16'hb3c5;
23692: douta=16'hbbc5;
23693: douta=16'hbbc4;
23694: douta=16'hbbe5;
23695: douta=16'hbbe5;
23696: douta=16'hc3e5;
23697: douta=16'hc3e6;
23698: douta=16'hc405;
23699: douta=16'hc405;
23700: douta=16'hc405;
23701: douta=16'hcc06;
23702: douta=16'hcc25;
23703: douta=16'hc404;
23704: douta=16'hc3c2;
23705: douta=16'hc3c2;
23706: douta=16'hc3c2;
23707: douta=16'hcc67;
23708: douta=16'hd4eb;
23709: douta=16'hd52d;
23710: douta=16'he6b5;
23711: douta=16'heef8;
23712: douta=16'hf79b;
23713: douta=16'hffbc;
23714: douta=16'hf759;
23715: douta=16'hf717;
23716: douta=16'hde11;
23717: douta=16'hdd6d;
23718: douta=16'hd4c9;
23719: douta=16'hcc22;
23720: douta=16'hcc02;
23721: douta=16'hcc04;
23722: douta=16'hd446;
23723: douta=16'hd467;
23724: douta=16'hd467;
23725: douta=16'hd466;
23726: douta=16'hd467;
23727: douta=16'hd467;
23728: douta=16'hcc86;
23729: douta=16'hd487;
23730: douta=16'hd466;
23731: douta=16'hb514;
23732: douta=16'hc595;
23733: douta=16'hcdd7;
23734: douta=16'hd5d7;
23735: douta=16'hcdd6;
23736: douta=16'hb577;
23737: douta=16'had77;
23738: douta=16'hbd97;
23739: douta=16'h94d6;
23740: douta=16'h8412;
23741: douta=16'h7bf2;
23742: douta=16'h6b70;
23743: douta=16'h7390;
23744: douta=16'h7390;
23745: douta=16'h6b4f;
23746: douta=16'h6b4e;
23747: douta=16'h6b2f;
23748: douta=16'h6b2f;
23749: douta=16'h41e7;
23750: douta=16'h5248;
23751: douta=16'h6b0c;
23752: douta=16'hbd31;
23753: douta=16'hd5d3;
23754: douta=16'hcd72;
23755: douta=16'hde56;
23756: douta=16'hde55;
23757: douta=16'he656;
23758: douta=16'he635;
23759: douta=16'hde35;
23760: douta=16'hd5d4;
23761: douta=16'ha4d3;
23762: douta=16'he616;
23763: douta=16'hc574;
23764: douta=16'hb514;
23765: douta=16'hacd4;
23766: douta=16'h9494;
23767: douta=16'h8c73;
23768: douta=16'h8c52;
23769: douta=16'h8c73;
23770: douta=16'h8432;
23771: douta=16'h7bf2;
23772: douta=16'h73d1;
23773: douta=16'h73b1;
23774: douta=16'h73d2;
23775: douta=16'h73f2;
23776: douta=16'h6bb1;
23777: douta=16'h6bb1;
23778: douta=16'h6bb2;
23779: douta=16'h39a6;
23780: douta=16'h49e8;
23781: douta=16'h5228;
23782: douta=16'h52ce;
23783: douta=16'h4aad;
23784: douta=16'h320b;
23785: douta=16'h31c9;
23786: douta=16'h1906;
23787: douta=16'h18e5;
23788: douta=16'h2925;
23789: douta=16'h59e4;
23790: douta=16'h6a25;
23791: douta=16'h6a26;
23792: douta=16'h6205;
23793: douta=16'h6205;
23794: douta=16'h59e6;
23795: douta=16'h5a06;
23796: douta=16'h51a5;
23797: douta=16'h51c5;
23798: douta=16'h51a5;
23799: douta=16'h51c6;
23800: douta=16'h51a6;
23801: douta=16'h49a5;
23802: douta=16'h49a6;
23803: douta=16'h49a6;
23804: douta=16'h4186;
23805: douta=16'h41a6;
23806: douta=16'h4166;
23807: douta=16'h3966;
23808: douta=16'hf6f8;
23809: douta=16'hf6f9;
23810: douta=16'hff5b;
23811: douta=16'hff3a;
23812: douta=16'hf6f8;
23813: douta=16'hff5a;
23814: douta=16'hcd73;
23815: douta=16'hacf5;
23816: douta=16'h9473;
23817: douta=16'had36;
23818: douta=16'ha4f5;
23819: douta=16'hb556;
23820: douta=16'hb535;
23821: douta=16'h9cd6;
23822: douta=16'h8474;
23823: douta=16'h7413;
23824: douta=16'h7c55;
23825: douta=16'h7c35;
23826: douta=16'h7c55;
23827: douta=16'h8496;
23828: douta=16'h8496;
23829: douta=16'h7c54;
23830: douta=16'h7c34;
23831: douta=16'h9518;
23832: douta=16'h4b0f;
23833: douta=16'h10e5;
23834: douta=16'h1906;
23835: douta=16'h10a5;
23836: douta=16'h08e5;
23837: douta=16'h10e6;
23838: douta=16'h10e6;
23839: douta=16'h10e5;
23840: douta=16'h08a4;
23841: douta=16'h10e5;
23842: douta=16'h10e5;
23843: douta=16'h10c4;
23844: douta=16'h10c4;
23845: douta=16'h2127;
23846: douta=16'h1906;
23847: douta=16'h2126;
23848: douta=16'h10a3;
23849: douta=16'h29ca;
23850: douta=16'h320a;
23851: douta=16'h3166;
23852: douta=16'h30e3;
23853: douta=16'h3103;
23854: douta=16'h4143;
23855: douta=16'h28c2;
23856: douta=16'h4100;
23857: douta=16'h4964;
23858: douta=16'h4984;
23859: douta=16'h51a4;
23860: douta=16'h61e4;
23861: douta=16'h6a04;
23862: douta=16'h6a24;
23863: douta=16'h6a24;
23864: douta=16'h6a04;
23865: douta=16'h7204;
23866: douta=16'h7244;
23867: douta=16'h7a44;
23868: douta=16'h7a44;
23869: douta=16'h82a4;
23870: douta=16'h8aa4;
23871: douta=16'h8ac5;
23872: douta=16'h92e4;
23873: douta=16'h9305;
23874: douta=16'h9b05;
23875: douta=16'h9b25;
23876: douta=16'ha344;
23877: douta=16'ha345;
23878: douta=16'hab65;
23879: douta=16'hb385;
23880: douta=16'hb385;
23881: douta=16'hb3c4;
23882: douta=16'hbbc4;
23883: douta=16'hb3c4;
23884: douta=16'hb3a4;
23885: douta=16'hbb83;
23886: douta=16'hb363;
23887: douta=16'hbbe4;
23888: douta=16'hc405;
23889: douta=16'hc489;
23890: douta=16'hd590;
23891: douta=16'he654;
23892: douta=16'heeb6;
23893: douta=16'hf79b;
23894: douta=16'hf79a;
23895: douta=16'hef59;
23896: douta=16'he673;
23897: douta=16'hde31;
23898: douta=16'hdd8d;
23899: douta=16'hd487;
23900: douta=16'hcc24;
23901: douta=16'hcbe3;
23902: douta=16'hcc04;
23903: douta=16'hcc25;
23904: douta=16'hcc25;
23905: douta=16'hcc46;
23906: douta=16'hd446;
23907: douta=16'hd466;
23908: douta=16'hd467;
23909: douta=16'hcc66;
23910: douta=16'hd467;
23911: douta=16'hd467;
23912: douta=16'hd466;
23913: douta=16'hcc66;
23914: douta=16'hcc66;
23915: douta=16'hd466;
23916: douta=16'hd466;
23917: douta=16'hd467;
23918: douta=16'hd466;
23919: douta=16'hd466;
23920: douta=16'hd467;
23921: douta=16'hcc66;
23922: douta=16'hd467;
23923: douta=16'hcc66;
23924: douta=16'h9c52;
23925: douta=16'ha4f5;
23926: douta=16'h9cd5;
23927: douta=16'h9cd5;
23928: douta=16'h9cb5;
23929: douta=16'h9cd5;
23930: douta=16'h9cd4;
23931: douta=16'h8432;
23932: douta=16'h9494;
23933: douta=16'h8432;
23934: douta=16'h7390;
23935: douta=16'h6b2f;
23936: douta=16'h6b2f;
23937: douta=16'h630e;
23938: douta=16'h49e7;
23939: douta=16'h6b0c;
23940: douta=16'h7b8d;
23941: douta=16'hb511;
23942: douta=16'hacd1;
23943: douta=16'hde15;
23944: douta=16'hde55;
23945: douta=16'hde35;
23946: douta=16'hcd92;
23947: douta=16'hde56;
23948: douta=16'hd5d5;
23949: douta=16'hd5f5;
23950: douta=16'hbd55;
23951: douta=16'had14;
23952: douta=16'hacf5;
23953: douta=16'h8c73;
23954: douta=16'h8412;
23955: douta=16'h8433;
23956: douta=16'h8c73;
23957: douta=16'h8412;
23958: douta=16'h7bd1;
23959: douta=16'h6b90;
23960: douta=16'h7bf1;
23961: douta=16'h73b0;
23962: douta=16'h632e;
23963: douta=16'h632e;
23964: douta=16'h632f;
23965: douta=16'h62cd;
23966: douta=16'h5acd;
23967: douta=16'h49e8;
23968: douta=16'h62a8;
23969: douta=16'h6b0b;
23970: douta=16'h732b;
23971: douta=16'hacb0;
23972: douta=16'hb4f0;
23973: douta=16'h62ed;
23974: douta=16'h3a2b;
23975: douta=16'h422a;
23976: douta=16'h422b;
23977: douta=16'h52ae;
23978: douta=16'h29ca;
23979: douta=16'h29c9;
23980: douta=16'h2147;
23981: douta=16'h08a4;
23982: douta=16'h7245;
23983: douta=16'h6a26;
23984: douta=16'h6226;
23985: douta=16'h6206;
23986: douta=16'h59c5;
23987: douta=16'h59e6;
23988: douta=16'h59c6;
23989: douta=16'h51c5;
23990: douta=16'h49a5;
23991: douta=16'h51c5;
23992: douta=16'h51a6;
23993: douta=16'h4986;
23994: douta=16'h49a6;
23995: douta=16'h4185;
23996: douta=16'h41a6;
23997: douta=16'h4186;
23998: douta=16'h4186;
23999: douta=16'h3966;
24000: douta=16'hf6f9;
24001: douta=16'hff5b;
24002: douta=16'hff7b;
24003: douta=16'hff7b;
24004: douta=16'hff5a;
24005: douta=16'heeb9;
24006: douta=16'hddf5;
24007: douta=16'hacf5;
24008: douta=16'ha4d5;
24009: douta=16'hb577;
24010: douta=16'hb555;
24011: douta=16'hb514;
24012: douta=16'hb535;
24013: douta=16'h9cd6;
24014: douta=16'h73f3;
24015: douta=16'h7413;
24016: douta=16'h7c55;
24017: douta=16'h7c55;
24018: douta=16'h7c55;
24019: douta=16'h8cb6;
24020: douta=16'h8476;
24021: douta=16'h7413;
24022: douta=16'h8496;
24023: douta=16'h322a;
24024: douta=16'h0001;
24025: douta=16'h0863;
24026: douta=16'h0883;
24027: douta=16'h08a4;
24028: douta=16'h10a4;
24029: douta=16'h10a5;
24030: douta=16'h10e5;
24031: douta=16'h2168;
24032: douta=16'h2188;
24033: douta=16'h2168;
24034: douta=16'h29ca;
24035: douta=16'h29ca;
24036: douta=16'h29cb;
24037: douta=16'h2105;
24038: douta=16'h20e4;
24039: douta=16'h2126;
24040: douta=16'h18c4;
24041: douta=16'h28a1;
24042: douta=16'h30e2;
24043: douta=16'h3902;
24044: douta=16'h4143;
24045: douta=16'h4143;
24046: douta=16'h5184;
24047: douta=16'h3102;
24048: douta=16'h59c4;
24049: douta=16'h61c4;
24050: douta=16'h59c4;
24051: douta=16'h59e3;
24052: douta=16'h6204;
24053: douta=16'h61e4;
24054: douta=16'h6a04;
24055: douta=16'h6a24;
24056: douta=16'h7224;
24057: douta=16'h7224;
24058: douta=16'h7a44;
24059: douta=16'h7a64;
24060: douta=16'h7a64;
24061: douta=16'h8284;
24062: douta=16'h8aa4;
24063: douta=16'h8ac4;
24064: douta=16'h9304;
24065: douta=16'h9b05;
24066: douta=16'h9b05;
24067: douta=16'h9b25;
24068: douta=16'ha345;
24069: douta=16'ha324;
24070: douta=16'ha323;
24071: douta=16'hab22;
24072: douta=16'hab43;
24073: douta=16'hbc07;
24074: douta=16'hbc48;
24075: douta=16'hcd2e;
24076: douta=16'he675;
24077: douta=16'hef18;
24078: douta=16'hef59;
24079: douta=16'hef58;
24080: douta=16'hef17;
24081: douta=16'he672;
24082: douta=16'hd56d;
24083: douta=16'hcce9;
24084: douta=16'hcc87;
24085: douta=16'hc3e2;
24086: douta=16'hc3e2;
24087: douta=16'hc3e2;
24088: douta=16'hcc05;
24089: douta=16'hcc25;
24090: douta=16'hcc45;
24091: douta=16'hcc47;
24092: douta=16'hcc66;
24093: douta=16'hcc45;
24094: douta=16'hcc46;
24095: douta=16'hcc45;
24096: douta=16'hcc46;
24097: douta=16'hcc66;
24098: douta=16'hcc66;
24099: douta=16'hcc66;
24100: douta=16'hcc46;
24101: douta=16'hd466;
24102: douta=16'hd466;
24103: douta=16'hd467;
24104: douta=16'hd466;
24105: douta=16'hd466;
24106: douta=16'hd487;
24107: douta=16'hd466;
24108: douta=16'hd466;
24109: douta=16'hd467;
24110: douta=16'hd467;
24111: douta=16'hd466;
24112: douta=16'hd467;
24113: douta=16'hd467;
24114: douta=16'hcc86;
24115: douta=16'hd486;
24116: douta=16'hd465;
24117: douta=16'h8c10;
24118: douta=16'h9cd4;
24119: douta=16'h9453;
24120: douta=16'h8c11;
24121: douta=16'h9453;
24122: douta=16'h83f1;
24123: douta=16'h8412;
24124: douta=16'h7bd1;
24125: douta=16'h7391;
24126: douta=16'h7390;
24127: douta=16'h41c8;
24128: douta=16'h49e7;
24129: douta=16'hacd0;
24130: douta=16'ha46e;
24131: douta=16'hc592;
24132: douta=16'hd5f4;
24133: douta=16'hb532;
24134: douta=16'he6b7;
24135: douta=16'he656;
24136: douta=16'hde55;
24137: douta=16'he656;
24138: douta=16'hcdb4;
24139: douta=16'hd5f6;
24140: douta=16'hcd95;
24141: douta=16'hbd75;
24142: douta=16'ha4f6;
24143: douta=16'h9cd5;
24144: douta=16'h8c74;
24145: douta=16'h94b4;
24146: douta=16'h8c53;
24147: douta=16'h8c74;
24148: douta=16'h8452;
24149: douta=16'h7bf1;
24150: douta=16'h73d1;
24151: douta=16'h6b4f;
24152: douta=16'h8411;
24153: douta=16'h6b6f;
24154: douta=16'h630d;
24155: douta=16'h630c;
24156: douta=16'h5229;
24157: douta=16'h93ed;
24158: douta=16'h940d;
24159: douta=16'h940e;
24160: douta=16'h8bcd;
24161: douta=16'ha46e;
24162: douta=16'ha48f;
24163: douta=16'hb4f1;
24164: douta=16'hb4d1;
24165: douta=16'h5acd;
24166: douta=16'h4209;
24167: douta=16'h31a8;
24168: douta=16'h3188;
24169: douta=16'h31ea;
24170: douta=16'h10e6;
24171: douta=16'h10e4;
24172: douta=16'h18e5;
24173: douta=16'h18e5;
24174: douta=16'h3966;
24175: douta=16'h6206;
24176: douta=16'h6205;
24177: douta=16'h59e5;
24178: douta=16'h59e6;
24179: douta=16'h59e6;
24180: douta=16'h51c5;
24181: douta=16'h51a5;
24182: douta=16'h49a5;
24183: douta=16'h49a5;
24184: douta=16'h49a6;
24185: douta=16'h49a6;
24186: douta=16'h4165;
24187: douta=16'h41a6;
24188: douta=16'h4185;
24189: douta=16'h4186;
24190: douta=16'h4166;
24191: douta=16'h4166;
24192: douta=16'hf6d8;
24193: douta=16'hff7b;
24194: douta=16'hff9c;
24195: douta=16'hffbd;
24196: douta=16'hff3a;
24197: douta=16'hde57;
24198: douta=16'hde16;
24199: douta=16'h9c94;
24200: douta=16'hb536;
24201: douta=16'hb577;
24202: douta=16'hbd75;
24203: douta=16'hb535;
24204: douta=16'had15;
24205: douta=16'h9cb5;
24206: douta=16'h73f3;
24207: douta=16'h7c34;
24208: douta=16'h7c54;
24209: douta=16'h8475;
24210: douta=16'h8496;
24211: douta=16'h8496;
24212: douta=16'h7c75;
24213: douta=16'h7c33;
24214: douta=16'h94f7;
24215: douta=16'h0084;
24216: douta=16'h1063;
24217: douta=16'h1967;
24218: douta=16'h10e5;
24219: douta=16'h10e5;
24220: douta=16'h10e6;
24221: douta=16'h1928;
24222: douta=16'h29ca;
24223: douta=16'h220c;
24224: douta=16'h21aa;
24225: douta=16'h21ca;
24226: douta=16'h2167;
24227: douta=16'h2105;
24228: douta=16'h20e4;
24229: douta=16'h2081;
24230: douta=16'h2081;
24231: douta=16'h20e3;
24232: douta=16'h20c3;
24233: douta=16'h3103;
24234: douta=16'h3923;
24235: douta=16'h4144;
24236: douta=16'h4163;
24237: douta=16'h4964;
24238: douta=16'h4984;
24239: douta=16'h3923;
24240: douta=16'h61c4;
24241: douta=16'h59c4;
24242: douta=16'h61c4;
24243: douta=16'h59e4;
24244: douta=16'h61e4;
24245: douta=16'h61e4;
24246: douta=16'h6a04;
24247: douta=16'h7204;
24248: douta=16'h7224;
24249: douta=16'h7224;
24250: douta=16'h7a44;
24251: douta=16'h7a64;
24252: douta=16'h7a64;
24253: douta=16'h82a4;
24254: douta=16'h8aa4;
24255: douta=16'h8ac4;
24256: douta=16'h92c4;
24257: douta=16'h92c4;
24258: douta=16'h92c4;
24259: douta=16'h92a2;
24260: douta=16'h9ae3;
24261: douta=16'ha324;
24262: douta=16'hb408;
24263: douta=16'hbcac;
24264: douta=16'hd5d1;
24265: douta=16'he6d6;
24266: douta=16'hef18;
24267: douta=16'hf77a;
24268: douta=16'hef16;
24269: douta=16'he652;
24270: douta=16'hde11;
24271: douta=16'hcce9;
24272: douta=16'hc486;
24273: douta=16'hc423;
24274: douta=16'hc3a3;
24275: douta=16'hc3c3;
24276: douta=16'hc3c3;
24277: douta=16'hc405;
24278: douta=16'hcc26;
24279: douta=16'hcc25;
24280: douta=16'hc445;
24281: douta=16'hcc45;
24282: douta=16'hcc45;
24283: douta=16'hcc45;
24284: douta=16'hcc45;
24285: douta=16'hd466;
24286: douta=16'hcc46;
24287: douta=16'hcc46;
24288: douta=16'hd446;
24289: douta=16'hcc46;
24290: douta=16'hd466;
24291: douta=16'hcc66;
24292: douta=16'hcc66;
24293: douta=16'hd466;
24294: douta=16'hd467;
24295: douta=16'hd466;
24296: douta=16'hcc66;
24297: douta=16'hd466;
24298: douta=16'hcc66;
24299: douta=16'hd466;
24300: douta=16'hd466;
24301: douta=16'hd467;
24302: douta=16'hd466;
24303: douta=16'hd466;
24304: douta=16'hd487;
24305: douta=16'hd467;
24306: douta=16'hd485;
24307: douta=16'hd466;
24308: douta=16'hdc65;
24309: douta=16'hb44c;
24310: douta=16'h9473;
24311: douta=16'h9c93;
24312: douta=16'h8bf2;
24313: douta=16'h83d1;
24314: douta=16'h7bb0;
24315: douta=16'h83d1;
24316: douta=16'h73b1;
24317: douta=16'h6b6f;
24318: douta=16'h5269;
24319: douta=16'h5a49;
24320: douta=16'hacf1;
24321: douta=16'h836c;
24322: douta=16'hc5b2;
24323: douta=16'hd614;
24324: douta=16'hde35;
24325: douta=16'hb512;
24326: douta=16'he696;
24327: douta=16'he656;
24328: douta=16'hde35;
24329: douta=16'he675;
24330: douta=16'hd5f4;
24331: douta=16'hc595;
24332: douta=16'hbd54;
24333: douta=16'hb515;
24334: douta=16'h9cb5;
24335: douta=16'h9cd5;
24336: douta=16'h8c74;
24337: douta=16'h8412;
24338: douta=16'h8453;
24339: douta=16'h8c73;
24340: douta=16'h8432;
24341: douta=16'h73d1;
24342: douta=16'h7390;
24343: douta=16'h632f;
24344: douta=16'h8c32;
24345: douta=16'h8c12;
24346: douta=16'h4a28;
24347: douta=16'h3103;
24348: douta=16'h41a5;
24349: douta=16'h93ec;
24350: douta=16'hb4ef;
24351: douta=16'hc572;
24352: douta=16'ha4b0;
24353: douta=16'ha46f;
24354: douta=16'ha48f;
24355: douta=16'hb4d1;
24356: douta=16'hacd1;
24357: douta=16'h630d;
24358: douta=16'h3a09;
24359: douta=16'h39e8;
24360: douta=16'h31a9;
24361: douta=16'h1906;
24362: douta=16'h18e4;
24363: douta=16'h18e5;
24364: douta=16'h1926;
24365: douta=16'h1926;
24366: douta=16'h18e5;
24367: douta=16'h6226;
24368: douta=16'h59e5;
24369: douta=16'h6206;
24370: douta=16'h59c5;
24371: douta=16'h59e6;
24372: douta=16'h51c6;
24373: douta=16'h51a5;
24374: douta=16'h49a5;
24375: douta=16'h49a5;
24376: douta=16'h49a6;
24377: douta=16'h4986;
24378: douta=16'h4186;
24379: douta=16'h41a6;
24380: douta=16'h41a6;
24381: douta=16'h4186;
24382: douta=16'h4186;
24383: douta=16'h4166;
24384: douta=16'hff3a;
24385: douta=16'hff9d;
24386: douta=16'hffbc;
24387: douta=16'hff9c;
24388: douta=16'hde35;
24389: douta=16'hd5f5;
24390: douta=16'hd617;
24391: douta=16'h9c93;
24392: douta=16'hb556;
24393: douta=16'hb576;
24394: douta=16'hb534;
24395: douta=16'hbd75;
24396: douta=16'had15;
24397: douta=16'h8c75;
24398: douta=16'h7c34;
24399: douta=16'h8455;
24400: douta=16'h8475;
24401: douta=16'h8455;
24402: douta=16'h8476;
24403: douta=16'h8455;
24404: douta=16'h8475;
24405: douta=16'h7c13;
24406: douta=16'h1082;
24407: douta=16'h2126;
24408: douta=16'h21c9;
24409: douta=16'h2189;
24410: douta=16'h2168;
24411: douta=16'h18e5;
24412: douta=16'h1882;
24413: douta=16'h1861;
24414: douta=16'h1882;
24415: douta=16'h1882;
24416: douta=16'h2082;
24417: douta=16'h20a2;
24418: douta=16'h20a2;
24419: douta=16'h20a2;
24420: douta=16'h20c2;
24421: douta=16'h28e2;
24422: douta=16'h2903;
24423: douta=16'h2946;
24424: douta=16'h3103;
24425: douta=16'h4143;
24426: douta=16'h4144;
24427: douta=16'h4143;
24428: douta=16'h4964;
24429: douta=16'h4963;
24430: douta=16'h4984;
24431: douta=16'h59c4;
24432: douta=16'h3923;
24433: douta=16'h59c4;
24434: douta=16'h59c4;
24435: douta=16'h61e4;
24436: douta=16'h61e4;
24437: douta=16'h6a04;
24438: douta=16'h6a24;
24439: douta=16'h69e3;
24440: douta=16'h61a3;
24441: douta=16'h61a3;
24442: douta=16'h7244;
24443: douta=16'h8307;
24444: douta=16'h9369;
24445: douta=16'hb4ae;
24446: douta=16'hc5b1;
24447: douta=16'hde74;
24448: douta=16'he6b5;
24449: douta=16'hde94;
24450: douta=16'hd612;
24451: douta=16'hc4ec;
24452: douta=16'hb429;
24453: douta=16'hb3e8;
24454: douta=16'hab64;
24455: douta=16'hab43;
24456: douta=16'hb343;
24457: douta=16'hb364;
24458: douta=16'hbbc4;
24459: douta=16'hbbe5;
24460: douta=16'hc405;
24461: douta=16'hc405;
24462: douta=16'hc406;
24463: douta=16'hc426;
24464: douta=16'hc426;
24465: douta=16'hc425;
24466: douta=16'hc425;
24467: douta=16'hc425;
24468: douta=16'hcc25;
24469: douta=16'hc425;
24470: douta=16'hcc25;
24471: douta=16'hcc26;
24472: douta=16'hcc46;
24473: douta=16'hcc46;
24474: douta=16'hcc46;
24475: douta=16'hcc45;
24476: douta=16'hcc46;
24477: douta=16'hcc66;
24478: douta=16'hcc66;
24479: douta=16'hcc47;
24480: douta=16'hcc66;
24481: douta=16'hcc66;
24482: douta=16'hcc66;
24483: douta=16'hd466;
24484: douta=16'hcc66;
24485: douta=16'hd466;
24486: douta=16'hd466;
24487: douta=16'hd466;
24488: douta=16'hd466;
24489: douta=16'hd466;
24490: douta=16'hd466;
24491: douta=16'hcc66;
24492: douta=16'hd466;
24493: douta=16'hd467;
24494: douta=16'hd466;
24495: douta=16'hd467;
24496: douta=16'hd467;
24497: douta=16'hd466;
24498: douta=16'hd466;
24499: douta=16'hd466;
24500: douta=16'hd468;
24501: douta=16'hd466;
24502: douta=16'hdc84;
24503: douta=16'hcc69;
24504: douta=16'h7c12;
24505: douta=16'h83b0;
24506: douta=16'h62ab;
24507: douta=16'h5249;
24508: douta=16'hacd0;
24509: douta=16'ha4b0;
24510: douta=16'h9c4e;
24511: douta=16'hde35;
24512: douta=16'h83ac;
24513: douta=16'hf6f8;
24514: douta=16'hde36;
24515: douta=16'hd615;
24516: douta=16'hde35;
24517: douta=16'hacd3;
24518: douta=16'hc575;
24519: douta=16'hb575;
24520: douta=16'hacf5;
24521: douta=16'h9495;
24522: douta=16'h8c94;
24523: douta=16'h94b4;
24524: douta=16'h8c74;
24525: douta=16'h8453;
24526: douta=16'h7bd1;
24527: douta=16'h7bf1;
24528: douta=16'h73d0;
24529: douta=16'h7c12;
24530: douta=16'h5b2f;
24531: douta=16'h52cd;
24532: douta=16'h7bf1;
24533: douta=16'h6b2c;
24534: douta=16'h3965;
24535: douta=16'h6ac9;
24536: douta=16'h62c9;
24537: douta=16'h5269;
24538: douta=16'h49c6;
24539: douta=16'hacb0;
24540: douta=16'hcd93;
24541: douta=16'hacaf;
24542: douta=16'ha46e;
24543: douta=16'h5aa9;
24544: douta=16'h838c;
24545: douta=16'hbd31;
24546: douta=16'hcdd3;
24547: douta=16'hb511;
24548: douta=16'hac91;
24549: douta=16'h83cf;
24550: douta=16'h6b4e;
24551: douta=16'h31c8;
24552: douta=16'h2126;
24553: douta=16'h2126;
24554: douta=16'h2126;
24555: douta=16'h10e5;
24556: douta=16'h29a8;
24557: douta=16'h29a9;
24558: douta=16'h1926;
24559: douta=16'h6226;
24560: douta=16'h6206;
24561: douta=16'h59e5;
24562: douta=16'h59e6;
24563: douta=16'h59e6;
24564: douta=16'h51c5;
24565: douta=16'h51a5;
24566: douta=16'h4985;
24567: douta=16'h4985;
24568: douta=16'h49a6;
24569: douta=16'h4986;
24570: douta=16'h49a6;
24571: douta=16'h49a6;
24572: douta=16'h4186;
24573: douta=16'h4166;
24574: douta=16'h3966;
24575: douta=16'h4166;
24576: douta=16'hf73a;
24577: douta=16'hff9c;
24578: douta=16'hffbc;
24579: douta=16'hffbd;
24580: douta=16'hd593;
24581: douta=16'hd5b3;
24582: douta=16'hb555;
24583: douta=16'hb556;
24584: douta=16'hb556;
24585: douta=16'hb556;
24586: douta=16'hbd75;
24587: douta=16'hb555;
24588: douta=16'ha516;
24589: douta=16'h8c95;
24590: douta=16'h8454;
24591: douta=16'h8455;
24592: douta=16'h8c96;
24593: douta=16'h7c34;
24594: douta=16'h8496;
24595: douta=16'h7c34;
24596: douta=16'h8454;
24597: douta=16'h94d6;
24598: douta=16'h1882;
24599: douta=16'h18c3;
24600: douta=16'h20a3;
24601: douta=16'h1061;
24602: douta=16'h1861;
24603: douta=16'h1882;
24604: douta=16'h1862;
24605: douta=16'h1883;
24606: douta=16'h18a2;
24607: douta=16'h18a2;
24608: douta=16'h20a2;
24609: douta=16'h20a2;
24610: douta=16'h20a2;
24611: douta=16'h28c3;
24612: douta=16'h20c2;
24613: douta=16'h28e3;
24614: douta=16'h2904;
24615: douta=16'h2947;
24616: douta=16'h3903;
24617: douta=16'h3903;
24618: douta=16'h4124;
24619: douta=16'h4163;
24620: douta=16'h4964;
24621: douta=16'h4984;
24622: douta=16'h49a4;
24623: douta=16'h5984;
24624: douta=16'h30e2;
24625: douta=16'h5162;
24626: douta=16'h5983;
24627: douta=16'h59c3;
24628: douta=16'h72a7;
24629: douta=16'h8329;
24630: douta=16'h8b8a;
24631: douta=16'hbd50;
24632: douta=16'hbd91;
24633: douta=16'hc5d2;
24634: douta=16'hc591;
24635: douta=16'hb4ee;
24636: douta=16'hac6c;
24637: douta=16'h9bc9;
24638: douta=16'h9306;
24639: douta=16'h8ac3;
24640: douta=16'h92a2;
24641: douta=16'h9282;
24642: douta=16'h9b04;
24643: douta=16'ha345;
24644: douta=16'hab85;
24645: douta=16'ha364;
24646: douta=16'hab65;
24647: douta=16'hb3a5;
24648: douta=16'hb3a5;
24649: douta=16'hbbc4;
24650: douta=16'hc405;
24651: douta=16'hbbe5;
24652: douta=16'hc405;
24653: douta=16'hc405;
24654: douta=16'hc406;
24655: douta=16'hc425;
24656: douta=16'hc425;
24657: douta=16'hc425;
24658: douta=16'hc425;
24659: douta=16'hc425;
24660: douta=16'hc425;
24661: douta=16'hc425;
24662: douta=16'hcc25;
24663: douta=16'hcc25;
24664: douta=16'hcc46;
24665: douta=16'hcc26;
24666: douta=16'hcc45;
24667: douta=16'hcc45;
24668: douta=16'hcc46;
24669: douta=16'hcc45;
24670: douta=16'hcc66;
24671: douta=16'hcc46;
24672: douta=16'hcc47;
24673: douta=16'hcc66;
24674: douta=16'hcc66;
24675: douta=16'hcc66;
24676: douta=16'hcc66;
24677: douta=16'hcc66;
24678: douta=16'hd467;
24679: douta=16'hd466;
24680: douta=16'hcc66;
24681: douta=16'hd466;
24682: douta=16'hd467;
24683: douta=16'hd467;
24684: douta=16'hd466;
24685: douta=16'hd466;
24686: douta=16'hd466;
24687: douta=16'hd466;
24688: douta=16'hd466;
24689: douta=16'hd467;
24690: douta=16'hd466;
24691: douta=16'hd466;
24692: douta=16'hd467;
24693: douta=16'hd467;
24694: douta=16'hcc86;
24695: douta=16'hd487;
24696: douta=16'hcc89;
24697: douta=16'h940d;
24698: douta=16'h9c4e;
24699: douta=16'hacb0;
24700: douta=16'hbd51;
24701: douta=16'hc573;
24702: douta=16'he676;
24703: douta=16'h9c0f;
24704: douta=16'hde16;
24705: douta=16'hd5f5;
24706: douta=16'hd615;
24707: douta=16'hcdd5;
24708: douta=16'hcdd6;
24709: douta=16'ha4b3;
24710: douta=16'ha4d3;
24711: douta=16'ha4f5;
24712: douta=16'h8c94;
24713: douta=16'h9494;
24714: douta=16'h8433;
24715: douta=16'h8c74;
24716: douta=16'h7bf2;
24717: douta=16'h7bd1;
24718: douta=16'h73b1;
24719: douta=16'h73d1;
24720: douta=16'h634e;
24721: douta=16'h6b6f;
24722: douta=16'h4a28;
24723: douta=16'h41a8;
24724: douta=16'h5247;
24725: douta=16'h83cd;
24726: douta=16'h942e;
24727: douta=16'h7b8b;
24728: douta=16'hb4f1;
24729: douta=16'hc551;
24730: douta=16'hacd0;
24731: douta=16'h83ac;
24732: douta=16'h730b;
24733: douta=16'hcd93;
24734: douta=16'hd5d4;
24735: douta=16'hde36;
24736: douta=16'hbd31;
24737: douta=16'h9c6f;
24738: douta=16'hac6f;
24739: douta=16'hc532;
24740: douta=16'hacd2;
24741: douta=16'h8431;
24742: douta=16'h6b4f;
24743: douta=16'h4ace;
24744: douta=16'h4a8d;
24745: douta=16'h3a0a;
24746: douta=16'h18e5;
24747: douta=16'h52ee;
24748: douta=16'h1906;
24749: douta=16'h1926;
24750: douta=16'h1927;
24751: douta=16'h6226;
24752: douta=16'h59e6;
24753: douta=16'h6206;
24754: douta=16'h59e6;
24755: douta=16'h51c5;
24756: douta=16'h51c6;
24757: douta=16'h51a5;
24758: douta=16'h49a5;
24759: douta=16'h49a5;
24760: douta=16'h49a5;
24761: douta=16'h4986;
24762: douta=16'h4185;
24763: douta=16'h4185;
24764: douta=16'h4186;
24765: douta=16'h4186;
24766: douta=16'h4166;
24767: douta=16'h3986;
24768: douta=16'hff5a;
24769: douta=16'hff9c;
24770: douta=16'hff9c;
24771: douta=16'hff7b;
24772: douta=16'hcd94;
24773: douta=16'hee78;
24774: douta=16'had35;
24775: douta=16'hb576;
24776: douta=16'hbd97;
24777: douta=16'hbd77;
24778: douta=16'hbd95;
24779: douta=16'hb555;
24780: douta=16'h9cf6;
24781: douta=16'h8c74;
24782: douta=16'h8475;
24783: douta=16'h8454;
24784: douta=16'h8496;
24785: douta=16'h7c54;
24786: douta=16'h8475;
24787: douta=16'h8454;
24788: douta=16'h8433;
24789: douta=16'h8454;
24790: douta=16'h20c3;
24791: douta=16'h18a2;
24792: douta=16'h18a3;
24793: douta=16'h1882;
24794: douta=16'h1082;
24795: douta=16'h1882;
24796: douta=16'h18a2;
24797: douta=16'h1882;
24798: douta=16'h1882;
24799: douta=16'h2082;
24800: douta=16'h20a2;
24801: douta=16'h20a2;
24802: douta=16'h20c2;
24803: douta=16'h20c2;
24804: douta=16'h28e2;
24805: douta=16'h30e2;
24806: douta=16'h2924;
24807: douta=16'h2967;
24808: douta=16'h3923;
24809: douta=16'h3923;
24810: douta=16'h4143;
24811: douta=16'h4123;
24812: douta=16'h4122;
24813: douta=16'h4122;
24814: douta=16'h4922;
24815: douta=16'h5184;
24816: douta=16'h3924;
24817: douta=16'h8329;
24818: douta=16'h8bab;
24819: douta=16'h944d;
24820: douta=16'hb531;
24821: douta=16'hbd72;
24822: douta=16'hbd71;
24823: douta=16'hac8e;
24824: douta=16'h9c2c;
24825: douta=16'h8b69;
24826: douta=16'h82c6;
24827: douta=16'h7a63;
24828: douta=16'h7a43;
24829: douta=16'h8244;
24830: douta=16'h8284;
24831: douta=16'h8ac5;
24832: douta=16'h9b05;
24833: douta=16'h9b05;
24834: douta=16'ha325;
24835: douta=16'ha345;
24836: douta=16'hab65;
24837: douta=16'hab65;
24838: douta=16'hab85;
24839: douta=16'hb3a5;
24840: douta=16'hb3a5;
24841: douta=16'hbc05;
24842: douta=16'hc406;
24843: douta=16'hc406;
24844: douta=16'hc406;
24845: douta=16'hc405;
24846: douta=16'hc405;
24847: douta=16'hcc66;
24848: douta=16'hc446;
24849: douta=16'hcc46;
24850: douta=16'hc405;
24851: douta=16'hc405;
24852: douta=16'hc405;
24853: douta=16'hcc25;
24854: douta=16'hcc46;
24855: douta=16'hcc25;
24856: douta=16'hcc25;
24857: douta=16'hcc26;
24858: douta=16'hcc45;
24859: douta=16'hcc45;
24860: douta=16'hcc46;
24861: douta=16'hcc45;
24862: douta=16'hcc46;
24863: douta=16'hcc66;
24864: douta=16'hd467;
24865: douta=16'hcc47;
24866: douta=16'hcc47;
24867: douta=16'hd466;
24868: douta=16'hcc66;
24869: douta=16'hcc66;
24870: douta=16'hd467;
24871: douta=16'hcc66;
24872: douta=16'hcc66;
24873: douta=16'hd466;
24874: douta=16'hd467;
24875: douta=16'hd467;
24876: douta=16'hd467;
24877: douta=16'hd467;
24878: douta=16'hd466;
24879: douta=16'hd487;
24880: douta=16'hd467;
24881: douta=16'hd467;
24882: douta=16'hd467;
24883: douta=16'hd467;
24884: douta=16'hd467;
24885: douta=16'hd487;
24886: douta=16'hd468;
24887: douta=16'hd467;
24888: douta=16'hd466;
24889: douta=16'hac8f;
24890: douta=16'hbd11;
24891: douta=16'hbd11;
24892: douta=16'hc592;
24893: douta=16'hd5f4;
24894: douta=16'he697;
24895: douta=16'hbd31;
24896: douta=16'heeb7;
24897: douta=16'hd5f6;
24898: douta=16'hd5d5;
24899: douta=16'hcdb5;
24900: douta=16'hc596;
24901: douta=16'h9c93;
24902: douta=16'h9c73;
24903: douta=16'h9494;
24904: douta=16'h8c53;
24905: douta=16'h8433;
24906: douta=16'h8412;
24907: douta=16'h7bf2;
24908: douta=16'h8433;
24909: douta=16'h7390;
24910: douta=16'h6b90;
24911: douta=16'h73b1;
24912: douta=16'h6b90;
24913: douta=16'h5228;
24914: douta=16'h3143;
24915: douta=16'h49c5;
24916: douta=16'h732c;
24917: douta=16'h7b6c;
24918: douta=16'hb510;
24919: douta=16'h9c2e;
24920: douta=16'h9c4f;
24921: douta=16'hb4d0;
24922: douta=16'hcdd3;
24923: douta=16'hcdb3;
24924: douta=16'ha46f;
24925: douta=16'ha46e;
24926: douta=16'hc551;
24927: douta=16'hd5f4;
24928: douta=16'he615;
24929: douta=16'hd5d4;
24930: douta=16'hcd73;
24931: douta=16'hacd2;
24932: douta=16'hacb1;
24933: douta=16'h8c73;
24934: douta=16'h6b6f;
24935: douta=16'h52ce;
24936: douta=16'h4a8d;
24937: douta=16'h3a2b;
24938: douta=16'h2167;
24939: douta=16'h3a0a;
24940: douta=16'h1926;
24941: douta=16'h2126;
24942: douta=16'h2188;
24943: douta=16'h6a46;
24944: douta=16'h6206;
24945: douta=16'h5a06;
24946: douta=16'h59c6;
24947: douta=16'h51e5;
24948: douta=16'h51c6;
24949: douta=16'h49a5;
24950: douta=16'h4985;
24951: douta=16'h49a5;
24952: douta=16'h49a5;
24953: douta=16'h49a6;
24954: douta=16'h4185;
24955: douta=16'h41a6;
24956: douta=16'h4186;
24957: douta=16'h4186;
24958: douta=16'h3986;
24959: douta=16'h3986;
24960: douta=16'hff7b;
24961: douta=16'hffbd;
24962: douta=16'hffbc;
24963: douta=16'hff7c;
24964: douta=16'hee98;
24965: douta=16'hd616;
24966: douta=16'h9c93;
24967: douta=16'hb596;
24968: douta=16'hb576;
24969: douta=16'hb555;
24970: douta=16'hbd75;
24971: douta=16'had36;
24972: douta=16'h8474;
24973: douta=16'h8454;
24974: douta=16'h8455;
24975: douta=16'h8475;
24976: douta=16'h8475;
24977: douta=16'h8496;
24978: douta=16'h7c54;
24979: douta=16'h8c96;
24980: douta=16'h8c96;
24981: douta=16'h1020;
24982: douta=16'h20c3;
24983: douta=16'h18a2;
24984: douta=16'h18c3;
24985: douta=16'h1882;
24986: douta=16'h1882;
24987: douta=16'h1882;
24988: douta=16'h1882;
24989: douta=16'h1882;
24990: douta=16'h1882;
24991: douta=16'h2082;
24992: douta=16'h20a2;
24993: douta=16'h2082;
24994: douta=16'h2081;
24995: douta=16'h2081;
24996: douta=16'h28c2;
24997: douta=16'h3124;
24998: douta=16'h2967;
24999: douta=16'h2967;
25000: douta=16'h7bae;
25001: douta=16'h7bae;
25002: douta=16'h840f;
25003: douta=16'h83cd;
25004: douta=16'h734a;
25005: douta=16'h6ae9;
25006: douta=16'h6245;
25007: douta=16'h6aa8;
25008: douta=16'h83cc;
25009: douta=16'h5983;
25010: douta=16'h5983;
25011: douta=16'h61a3;
25012: douta=16'h61e4;
25013: douta=16'h6a04;
25014: douta=16'h6a24;
25015: douta=16'h7223;
25016: douta=16'h7223;
25017: douta=16'h7244;
25018: douta=16'h7a64;
25019: douta=16'h7a63;
25020: douta=16'h8284;
25021: douta=16'h8aa4;
25022: douta=16'h8ac4;
25023: douta=16'h92e5;
25024: douta=16'h9b05;
25025: douta=16'h9b26;
25026: douta=16'h9b25;
25027: douta=16'ha345;
25028: douta=16'hab64;
25029: douta=16'hab65;
25030: douta=16'hb385;
25031: douta=16'hb385;
25032: douta=16'hbbc6;
25033: douta=16'hbc05;
25034: douta=16'hbbe5;
25035: douta=16'hbbe5;
25036: douta=16'hc406;
25037: douta=16'hc406;
25038: douta=16'hc406;
25039: douta=16'hc425;
25040: douta=16'hc445;
25041: douta=16'hc425;
25042: douta=16'hc405;
25043: douta=16'hc425;
25044: douta=16'hcc25;
25045: douta=16'hc425;
25046: douta=16'hc425;
25047: douta=16'hcc26;
25048: douta=16'hcc25;
25049: douta=16'hcc26;
25050: douta=16'hcc46;
25051: douta=16'hcc46;
25052: douta=16'hcc47;
25053: douta=16'hcc46;
25054: douta=16'hcc46;
25055: douta=16'hcc47;
25056: douta=16'hcc66;
25057: douta=16'hcc46;
25058: douta=16'hcc47;
25059: douta=16'hd467;
25060: douta=16'hcc66;
25061: douta=16'hcc47;
25062: douta=16'hd467;
25063: douta=16'hd467;
25064: douta=16'hd467;
25065: douta=16'hd466;
25066: douta=16'hd466;
25067: douta=16'hd467;
25068: douta=16'hd467;
25069: douta=16'hd467;
25070: douta=16'hd467;
25071: douta=16'hd467;
25072: douta=16'hd467;
25073: douta=16'hd467;
25074: douta=16'hd467;
25075: douta=16'hd466;
25076: douta=16'hd467;
25077: douta=16'hd467;
25078: douta=16'hd467;
25079: douta=16'hd467;
25080: douta=16'hd487;
25081: douta=16'hac4d;
25082: douta=16'hac91;
25083: douta=16'ha491;
25084: douta=16'hc573;
25085: douta=16'hc594;
25086: douta=16'hd616;
25087: douta=16'hc5b6;
25088: douta=16'had16;
25089: douta=16'had36;
25090: douta=16'ha516;
25091: douta=16'h9cd6;
25092: douta=16'h9495;
25093: douta=16'h73f2;
25094: douta=16'h6b91;
25095: douta=16'h8c52;
25096: douta=16'h7c11;
25097: douta=16'h73b1;
25098: douta=16'h73b0;
25099: douta=16'h6b70;
25100: douta=16'h630d;
25101: douta=16'h41e7;
25102: douta=16'h5aa9;
25103: douta=16'h62ca;
25104: douta=16'h8bcd;
25105: douta=16'h8c0e;
25106: douta=16'h9c6f;
25107: douta=16'h942e;
25108: douta=16'hc572;
25109: douta=16'hbd31;
25110: douta=16'h836c;
25111: douta=16'hcdd4;
25112: douta=16'hcdd3;
25113: douta=16'hcdd4;
25114: douta=16'hc572;
25115: douta=16'hcdb4;
25116: douta=16'hd615;
25117: douta=16'hde35;
25118: douta=16'he656;
25119: douta=16'hd614;
25120: douta=16'hcd93;
25121: douta=16'hc533;
25122: douta=16'hbcf3;
25123: douta=16'h8c93;
25124: douta=16'h8c74;
25125: douta=16'h9494;
25126: douta=16'h73b1;
25127: douta=16'h6350;
25128: douta=16'h634f;
25129: douta=16'h5b0f;
25130: douta=16'h4aae;
25131: douta=16'h21a8;
25132: douta=16'h08a5;
25133: douta=16'h10e4;
25134: douta=16'h10e4;
25135: douta=16'h3965;
25136: douta=16'h59e5;
25137: douta=16'h5a26;
25138: douta=16'h51c6;
25139: douta=16'h59c6;
25140: douta=16'h51c5;
25141: douta=16'h49a5;
25142: douta=16'h49a6;
25143: douta=16'h49a6;
25144: douta=16'h49a6;
25145: douta=16'h49a6;
25146: douta=16'h4185;
25147: douta=16'h4186;
25148: douta=16'h4166;
25149: douta=16'h4186;
25150: douta=16'h3966;
25151: douta=16'h3986;
25152: douta=16'hff7c;
25153: douta=16'hffdd;
25154: douta=16'hfffe;
25155: douta=16'hde15;
25156: douta=16'he657;
25157: douta=16'hb555;
25158: douta=16'h9453;
25159: douta=16'hb576;
25160: douta=16'hbd75;
25161: douta=16'hc596;
25162: douta=16'hbd76;
25163: douta=16'ha516;
25164: douta=16'h9495;
25165: douta=16'h8475;
25166: douta=16'h8c75;
25167: douta=16'h8474;
25168: douta=16'h8455;
25169: douta=16'h8475;
25170: douta=16'h7c33;
25171: douta=16'h8495;
25172: douta=16'h324b;
25173: douta=16'h29c8;
25174: douta=16'h1861;
25175: douta=16'h18a2;
25176: douta=16'h1882;
25177: douta=16'h1061;
25178: douta=16'h1040;
25179: douta=16'h1061;
25180: douta=16'h1861;
25181: douta=16'h20c3;
25182: douta=16'h20c3;
25183: douta=16'h3145;
25184: douta=16'h39a6;
25185: douta=16'h39c7;
25186: douta=16'h5269;
25187: douta=16'h5269;
25188: douta=16'h5248;
25189: douta=16'h4a27;
25190: douta=16'h2967;
25191: douta=16'h2967;
25192: douta=16'h4123;
25193: douta=16'h3902;
25194: douta=16'h3902;
25195: douta=16'h4142;
25196: douta=16'h4963;
25197: douta=16'h4964;
25198: douta=16'h51a4;
25199: douta=16'h6aea;
25200: douta=16'h834a;
25201: douta=16'h6a04;
25202: douta=16'h61e4;
25203: douta=16'h61e4;
25204: douta=16'h6a24;
25205: douta=16'h7224;
25206: douta=16'h6a24;
25207: douta=16'h7224;
25208: douta=16'h7244;
25209: douta=16'h7224;
25210: douta=16'h8284;
25211: douta=16'h7a63;
25212: douta=16'h8284;
25213: douta=16'h8aa4;
25214: douta=16'h8ac5;
25215: douta=16'h92e5;
25216: douta=16'h9b05;
25217: douta=16'h9b05;
25218: douta=16'ha325;
25219: douta=16'hab65;
25220: douta=16'hab65;
25221: douta=16'hab65;
25222: douta=16'hb385;
25223: douta=16'hb3a5;
25224: douta=16'hb3a5;
25225: douta=16'hbbc4;
25226: douta=16'hbbc5;
25227: douta=16'hbbc6;
25228: douta=16'hbbc5;
25229: douta=16'hc405;
25230: douta=16'hc405;
25231: douta=16'hc405;
25232: douta=16'hc405;
25233: douta=16'hc426;
25234: douta=16'hc405;
25235: douta=16'hc405;
25236: douta=16'hc405;
25237: douta=16'hcc26;
25238: douta=16'hc425;
25239: douta=16'hcc25;
25240: douta=16'hcc26;
25241: douta=16'hcc26;
25242: douta=16'hcc46;
25243: douta=16'hcc46;
25244: douta=16'hcc46;
25245: douta=16'hcc46;
25246: douta=16'hcc66;
25247: douta=16'hcc46;
25248: douta=16'hcc66;
25249: douta=16'hcc47;
25250: douta=16'hd467;
25251: douta=16'hd467;
25252: douta=16'hd467;
25253: douta=16'hd466;
25254: douta=16'hcc47;
25255: douta=16'hd466;
25256: douta=16'hd466;
25257: douta=16'hd466;
25258: douta=16'hcc66;
25259: douta=16'hd466;
25260: douta=16'hcc66;
25261: douta=16'hd467;
25262: douta=16'hd467;
25263: douta=16'hd467;
25264: douta=16'hd467;
25265: douta=16'hd467;
25266: douta=16'hd467;
25267: douta=16'hd467;
25268: douta=16'hd467;
25269: douta=16'hd467;
25270: douta=16'hd487;
25271: douta=16'hd487;
25272: douta=16'hd467;
25273: douta=16'hd486;
25274: douta=16'h942f;
25275: douta=16'ha4b1;
25276: douta=16'ha493;
25277: douta=16'ha4d3;
25278: douta=16'hc596;
25279: douta=16'had16;
25280: douta=16'h94b5;
25281: douta=16'h9cd5;
25282: douta=16'h83f2;
25283: douta=16'h7bf2;
25284: douta=16'h7bf1;
25285: douta=16'h73d1;
25286: douta=16'h6bb1;
25287: douta=16'h6b70;
25288: douta=16'h6b70;
25289: douta=16'h5acb;
25290: douta=16'h526a;
25291: douta=16'h41e7;
25292: douta=16'h5a8a;
25293: douta=16'h940e;
25294: douta=16'h9c2e;
25295: douta=16'hb4d0;
25296: douta=16'h9c4e;
25297: douta=16'hc550;
25298: douta=16'hbd10;
25299: douta=16'hc551;
25300: douta=16'hc552;
25301: douta=16'hbd52;
25302: douta=16'hd5f4;
25303: douta=16'hbd30;
25304: douta=16'hd635;
25305: douta=16'hde35;
25306: douta=16'hde35;
25307: douta=16'hde35;
25308: douta=16'hd615;
25309: douta=16'hcd94;
25310: douta=16'hc573;
25311: douta=16'hbd53;
25312: douta=16'hb4f4;
25313: douta=16'h9cb4;
25314: douta=16'h9cb4;
25315: douta=16'h8c73;
25316: douta=16'h8c93;
25317: douta=16'h8c74;
25318: douta=16'h7bf3;
25319: douta=16'h6b6f;
25320: douta=16'h5b2e;
25321: douta=16'h4aad;
25322: douta=16'h424b;
25323: douta=16'h39ea;
25324: douta=16'h83f1;
25325: douta=16'h3189;
25326: douta=16'h1905;
25327: douta=16'h1905;
25328: douta=16'h1905;
25329: douta=16'h51c5;
25330: douta=16'h51c6;
25331: douta=16'h51c5;
25332: douta=16'h51c6;
25333: douta=16'h51e6;
25334: douta=16'h49a6;
25335: douta=16'h49a6;
25336: douta=16'h49a6;
25337: douta=16'h49a6;
25338: douta=16'h4165;
25339: douta=16'h4186;
25340: douta=16'h4166;
25341: douta=16'h4166;
25342: douta=16'h4166;
25343: douta=16'h3986;
25344: douta=16'hff7c;
25345: douta=16'hffbd;
25346: douta=16'hffff;
25347: douta=16'hd5d5;
25348: douta=16'hd617;
25349: douta=16'had15;
25350: douta=16'h9c73;
25351: douta=16'hbd96;
25352: douta=16'hbd75;
25353: douta=16'hc5b6;
25354: douta=16'hb556;
25355: douta=16'h9cb5;
25356: douta=16'h94b5;
25357: douta=16'h8c75;
25358: douta=16'h8475;
25359: douta=16'h8454;
25360: douta=16'h8475;
25361: douta=16'h7c54;
25362: douta=16'h7c33;
25363: douta=16'h4a8b;
25364: douta=16'h1062;
25365: douta=16'h3a6a;
25366: douta=16'h2126;
25367: douta=16'h1882;
25368: douta=16'h1841;
25369: douta=16'h18a3;
25370: douta=16'h18c3;
25371: douta=16'h2124;
25372: douta=16'h2965;
25373: douta=16'h29a6;
25374: douta=16'h31a7;
25375: douta=16'h39e8;
25376: douta=16'h39c7;
25377: douta=16'h39a6;
25378: douta=16'h3965;
25379: douta=16'h3144;
25380: douta=16'h3103;
25381: douta=16'h30e2;
25382: douta=16'h31a7;
25383: douta=16'h2967;
25384: douta=16'h3903;
25385: douta=16'h4123;
25386: douta=16'h4143;
25387: douta=16'h4963;
25388: douta=16'h5184;
25389: douta=16'h49a4;
25390: douta=16'h51a3;
25391: douta=16'h734c;
25392: douta=16'h7b08;
25393: douta=16'h6a03;
25394: douta=16'h61e4;
25395: douta=16'h69e4;
25396: douta=16'h6a04;
25397: douta=16'h7224;
25398: douta=16'h7224;
25399: douta=16'h7224;
25400: douta=16'h7224;
25401: douta=16'h7244;
25402: douta=16'h7a64;
25403: douta=16'h82a4;
25404: douta=16'h8284;
25405: douta=16'h8aa4;
25406: douta=16'h8ac4;
25407: douta=16'h92e4;
25408: douta=16'h9b26;
25409: douta=16'h9b25;
25410: douta=16'h9b25;
25411: douta=16'ha365;
25412: douta=16'hab65;
25413: douta=16'hab65;
25414: douta=16'hb385;
25415: douta=16'hb385;
25416: douta=16'hb3c5;
25417: douta=16'hbbc5;
25418: douta=16'hb3c5;
25419: douta=16'hbbc6;
25420: douta=16'hbbe5;
25421: douta=16'hbbe5;
25422: douta=16'hbbe5;
25423: douta=16'hc405;
25424: douta=16'hc405;
25425: douta=16'hc426;
25426: douta=16'hc425;
25427: douta=16'hc425;
25428: douta=16'hc425;
25429: douta=16'hc425;
25430: douta=16'hc425;
25431: douta=16'hcc25;
25432: douta=16'hcc46;
25433: douta=16'hcc46;
25434: douta=16'hcc46;
25435: douta=16'hcc46;
25436: douta=16'hcc46;
25437: douta=16'hcc47;
25438: douta=16'hcc66;
25439: douta=16'hcc46;
25440: douta=16'hcc66;
25441: douta=16'hcc47;
25442: douta=16'hcc46;
25443: douta=16'hcc47;
25444: douta=16'hd467;
25445: douta=16'hcc66;
25446: douta=16'hd467;
25447: douta=16'hcc66;
25448: douta=16'hd466;
25449: douta=16'hd467;
25450: douta=16'hd466;
25451: douta=16'hd466;
25452: douta=16'hcc66;
25453: douta=16'hd467;
25454: douta=16'hd487;
25455: douta=16'hd467;
25456: douta=16'hd467;
25457: douta=16'hd467;
25458: douta=16'hd467;
25459: douta=16'hd467;
25460: douta=16'hd467;
25461: douta=16'hd467;
25462: douta=16'hd487;
25463: douta=16'hd466;
25464: douta=16'hd487;
25465: douta=16'hd487;
25466: douta=16'h9c0d;
25467: douta=16'h9430;
25468: douta=16'h9c72;
25469: douta=16'h9c72;
25470: douta=16'hb536;
25471: douta=16'ha4d5;
25472: douta=16'h9495;
25473: douta=16'h8c74;
25474: douta=16'h7390;
25475: douta=16'h73d1;
25476: douta=16'h73d0;
25477: douta=16'h73b0;
25478: douta=16'h6b90;
25479: douta=16'h6b90;
25480: douta=16'h634e;
25481: douta=16'h1881;
25482: douta=16'h3124;
25483: douta=16'h7b6e;
25484: douta=16'h942f;
25485: douta=16'ha46e;
25486: douta=16'hb531;
25487: douta=16'hc571;
25488: douta=16'hb4ef;
25489: douta=16'hcd92;
25490: douta=16'hc531;
25491: douta=16'hd5b3;
25492: douta=16'hc573;
25493: douta=16'hc573;
25494: douta=16'hde36;
25495: douta=16'hcdd4;
25496: douta=16'hd616;
25497: douta=16'hcdb4;
25498: douta=16'hde15;
25499: douta=16'hcdd4;
25500: douta=16'hde35;
25501: douta=16'hd5b4;
25502: douta=16'hc554;
25503: douta=16'hb514;
25504: douta=16'ha4d5;
25505: douta=16'h9494;
25506: douta=16'h9c94;
25507: douta=16'h9494;
25508: douta=16'h8c93;
25509: douta=16'h8c74;
25510: douta=16'h7bf3;
25511: douta=16'h6b91;
25512: douta=16'h634f;
25513: douta=16'h424c;
25514: douta=16'h31a8;
25515: douta=16'h39ea;
25516: douta=16'h9c92;
25517: douta=16'h424b;
25518: douta=16'h2189;
25519: douta=16'h1905;
25520: douta=16'h1926;
25521: douta=16'h41a6;
25522: douta=16'h51c6;
25523: douta=16'h51c6;
25524: douta=16'h51c6;
25525: douta=16'h51c5;
25526: douta=16'h49a6;
25527: douta=16'h49a6;
25528: douta=16'h49a6;
25529: douta=16'h4185;
25530: douta=16'h4185;
25531: douta=16'h4166;
25532: douta=16'h4186;
25533: douta=16'h3945;
25534: douta=16'h4166;
25535: douta=16'h4186;
25536: douta=16'hff9c;
25537: douta=16'hffbd;
25538: douta=16'hf71a;
25539: douta=16'he698;
25540: douta=16'hbd96;
25541: douta=16'ha4b4;
25542: douta=16'hb535;
25543: douta=16'hb514;
25544: douta=16'hcdb5;
25545: douta=16'hc5b6;
25546: douta=16'h94b4;
25547: douta=16'h8433;
25548: douta=16'h8c74;
25549: douta=16'h8474;
25550: douta=16'h8454;
25551: douta=16'h8474;
25552: douta=16'h7413;
25553: douta=16'h7c13;
25554: douta=16'h9d17;
25555: douta=16'h18a2;
25556: douta=16'h20a2;
25557: douta=16'h18c3;
25558: douta=16'h1882;
25559: douta=16'h18a3;
25560: douta=16'h1883;
25561: douta=16'h1861;
25562: douta=16'h1882;
25563: douta=16'h1881;
25564: douta=16'h1881;
25565: douta=16'h2082;
25566: douta=16'h2082;
25567: douta=16'h20a2;
25568: douta=16'h20a2;
25569: douta=16'h20a2;
25570: douta=16'h28c2;
25571: douta=16'h28c2;
25572: douta=16'h28e2;
25573: douta=16'h2903;
25574: douta=16'h2988;
25575: douta=16'h1905;
25576: douta=16'h4143;
25577: douta=16'h4143;
25578: douta=16'h4143;
25579: douta=16'h4964;
25580: douta=16'h5184;
25581: douta=16'h51a4;
25582: douta=16'h5163;
25583: douta=16'h8c91;
25584: douta=16'h61c4;
25585: douta=16'h51a4;
25586: douta=16'h6a04;
25587: douta=16'h69e4;
25588: douta=16'h6a04;
25589: douta=16'h7224;
25590: douta=16'h7244;
25591: douta=16'h7224;
25592: douta=16'h7224;
25593: douta=16'h7a44;
25594: douta=16'h7a64;
25595: douta=16'h8285;
25596: douta=16'h82a4;
25597: douta=16'h8ac5;
25598: douta=16'h8ae4;
25599: douta=16'h9304;
25600: douta=16'h9b05;
25601: douta=16'h9b25;
25602: douta=16'ha345;
25603: douta=16'hab45;
25604: douta=16'hab65;
25605: douta=16'hab65;
25606: douta=16'hb385;
25607: douta=16'hb3a5;
25608: douta=16'hb3a5;
25609: douta=16'hbbc5;
25610: douta=16'hbbc5;
25611: douta=16'hbbc6;
25612: douta=16'hbbe5;
25613: douta=16'hbc06;
25614: douta=16'hbc06;
25615: douta=16'hc405;
25616: douta=16'hc406;
25617: douta=16'hc426;
25618: douta=16'hc405;
25619: douta=16'hc425;
25620: douta=16'hc425;
25621: douta=16'hcc26;
25622: douta=16'hcc26;
25623: douta=16'hcc25;
25624: douta=16'hcc46;
25625: douta=16'hcc46;
25626: douta=16'hcc46;
25627: douta=16'hcc47;
25628: douta=16'hcc46;
25629: douta=16'hcc46;
25630: douta=16'hcc46;
25631: douta=16'hcc46;
25632: douta=16'hcc47;
25633: douta=16'hd467;
25634: douta=16'hcc47;
25635: douta=16'hd467;
25636: douta=16'hcc66;
25637: douta=16'hd467;
25638: douta=16'hd467;
25639: douta=16'hcc47;
25640: douta=16'hd466;
25641: douta=16'hcc66;
25642: douta=16'hd467;
25643: douta=16'hd467;
25644: douta=16'hd467;
25645: douta=16'hd467;
25646: douta=16'hd467;
25647: douta=16'hd467;
25648: douta=16'hd487;
25649: douta=16'hd467;
25650: douta=16'hd467;
25651: douta=16'hd467;
25652: douta=16'hd467;
25653: douta=16'hd467;
25654: douta=16'hd487;
25655: douta=16'hd468;
25656: douta=16'hd488;
25657: douta=16'hd468;
25658: douta=16'hbd0e;
25659: douta=16'hc614;
25660: douta=16'h9430;
25661: douta=16'h9451;
25662: douta=16'h9452;
25663: douta=16'h7bb0;
25664: douta=16'h7bd0;
25665: douta=16'h736f;
25666: douta=16'h6b4e;
25667: douta=16'h630e;
25668: douta=16'h632e;
25669: douta=16'h41a6;
25670: douta=16'h3124;
25671: douta=16'h940e;
25672: douta=16'h732a;
25673: douta=16'h9c4f;
25674: douta=16'hacaf;
25675: douta=16'hbd72;
25676: douta=16'hb531;
25677: douta=16'hc593;
25678: douta=16'hd5f4;
25679: douta=16'hcdd3;
25680: douta=16'hd5f3;
25681: douta=16'hd5f4;
25682: douta=16'hde15;
25683: douta=16'hde36;
25684: douta=16'hb513;
25685: douta=16'hc5b4;
25686: douta=16'he657;
25687: douta=16'hbd34;
25688: douta=16'hb534;
25689: douta=16'hc575;
25690: douta=16'hc574;
25691: douta=16'hb534;
25692: douta=16'hbd54;
25693: douta=16'hacf4;
25694: douta=16'ha4d4;
25695: douta=16'h9cb4;
25696: douta=16'h9494;
25697: douta=16'h8c73;
25698: douta=16'h8c53;
25699: douta=16'h7bf2;
25700: douta=16'h73b1;
25701: douta=16'h73b1;
25702: douta=16'h62cc;
25703: douta=16'h41c6;
25704: douta=16'h3144;
25705: douta=16'h3985;
25706: douta=16'h8369;
25707: douta=16'h4208;
25708: douta=16'h426c;
25709: douta=16'h734e;
25710: douta=16'h18e5;
25711: douta=16'h2189;
25712: douta=16'h18e5;
25713: douta=16'h1907;
25714: douta=16'h51e5;
25715: douta=16'h59e6;
25716: douta=16'h51c5;
25717: douta=16'h49c6;
25718: douta=16'h49a6;
25719: douta=16'h49a6;
25720: douta=16'h4185;
25721: douta=16'h49a6;
25722: douta=16'h4185;
25723: douta=16'h4166;
25724: douta=16'h4166;
25725: douta=16'h4166;
25726: douta=16'h3966;
25727: douta=16'h3966;
25728: douta=16'hffbd;
25729: douta=16'hffdd;
25730: douta=16'hde77;
25731: douta=16'he677;
25732: douta=16'had14;
25733: douta=16'ha4b4;
25734: douta=16'hb554;
25735: douta=16'hc595;
25736: douta=16'hc595;
25737: douta=16'hbd76;
25738: douta=16'h8453;
25739: douta=16'h8c74;
25740: douta=16'h8c94;
25741: douta=16'h8474;
25742: douta=16'h8454;
25743: douta=16'h8474;
25744: douta=16'h7c13;
25745: douta=16'h8454;
25746: douta=16'h8cb6;
25747: douta=16'h20e3;
25748: douta=16'h18c3;
25749: douta=16'h18c3;
25750: douta=16'h20c3;
25751: douta=16'h1082;
25752: douta=16'h1882;
25753: douta=16'h1882;
25754: douta=16'h1882;
25755: douta=16'h1881;
25756: douta=16'h20a2;
25757: douta=16'h20a2;
25758: douta=16'h20a2;
25759: douta=16'h2082;
25760: douta=16'h20a2;
25761: douta=16'h20c2;
25762: douta=16'h28e3;
25763: douta=16'h28e2;
25764: douta=16'h30e3;
25765: douta=16'h3125;
25766: douta=16'h2988;
25767: douta=16'h18e5;
25768: douta=16'h4143;
25769: douta=16'h4143;
25770: douta=16'h4963;
25771: douta=16'h4963;
25772: douta=16'h51a4;
25773: douta=16'h51a4;
25774: douta=16'h5183;
25775: douta=16'h9d13;
25776: douta=16'h5983;
25777: douta=16'h4964;
25778: douta=16'h7224;
25779: douta=16'h7204;
25780: douta=16'h7224;
25781: douta=16'h7244;
25782: douta=16'h7244;
25783: douta=16'h7224;
25784: douta=16'h7224;
25785: douta=16'h7244;
25786: douta=16'h8284;
25787: douta=16'h8284;
25788: douta=16'h8283;
25789: douta=16'h8ac5;
25790: douta=16'h92c4;
25791: douta=16'h9305;
25792: douta=16'h9b05;
25793: douta=16'ha325;
25794: douta=16'ha325;
25795: douta=16'hab45;
25796: douta=16'hab85;
25797: douta=16'hab65;
25798: douta=16'hb385;
25799: douta=16'hb385;
25800: douta=16'hb3c5;
25801: douta=16'hbbe6;
25802: douta=16'hbbe5;
25803: douta=16'hbbe5;
25804: douta=16'hbbe5;
25805: douta=16'hbc06;
25806: douta=16'hbbe5;
25807: douta=16'hc405;
25808: douta=16'hc426;
25809: douta=16'hc426;
25810: douta=16'hc406;
25811: douta=16'hc425;
25812: douta=16'hc425;
25813: douta=16'hc425;
25814: douta=16'hc425;
25815: douta=16'hcc26;
25816: douta=16'hcc46;
25817: douta=16'hcc46;
25818: douta=16'hcc46;
25819: douta=16'hcc46;
25820: douta=16'hcc47;
25821: douta=16'hcc46;
25822: douta=16'hcc66;
25823: douta=16'hd466;
25824: douta=16'hcc46;
25825: douta=16'hd467;
25826: douta=16'hd467;
25827: douta=16'hd467;
25828: douta=16'hcc66;
25829: douta=16'hd467;
25830: douta=16'hd467;
25831: douta=16'hd467;
25832: douta=16'hd466;
25833: douta=16'hd467;
25834: douta=16'hd467;
25835: douta=16'hd467;
25836: douta=16'hd467;
25837: douta=16'hd467;
25838: douta=16'hd467;
25839: douta=16'hd467;
25840: douta=16'hd467;
25841: douta=16'hd467;
25842: douta=16'hd467;
25843: douta=16'hd468;
25844: douta=16'hd467;
25845: douta=16'hd467;
25846: douta=16'hd467;
25847: douta=16'hd487;
25848: douta=16'hd467;
25849: douta=16'hd468;
25850: douta=16'hbccd;
25851: douta=16'hce56;
25852: douta=16'h9430;
25853: douta=16'h9410;
25854: douta=16'h8bd0;
25855: douta=16'h734e;
25856: douta=16'h734e;
25857: douta=16'h6b4e;
25858: douta=16'h62cc;
25859: douta=16'h49e6;
25860: douta=16'h41a5;
25861: douta=16'h8c0e;
25862: douta=16'hd614;
25863: douta=16'h734b;
25864: douta=16'hacaf;
25865: douta=16'hbd30;
25866: douta=16'hc571;
25867: douta=16'hcdb3;
25868: douta=16'hbd52;
25869: douta=16'he676;
25870: douta=16'hd614;
25871: douta=16'he676;
25872: douta=16'hde15;
25873: douta=16'hde15;
25874: douta=16'hde35;
25875: douta=16'hd5f4;
25876: douta=16'hb513;
25877: douta=16'ha4d3;
25878: douta=16'hc596;
25879: douta=16'h9c93;
25880: douta=16'hb534;
25881: douta=16'hacf4;
25882: douta=16'hb515;
25883: douta=16'hb514;
25884: douta=16'ha4f4;
25885: douta=16'h8c74;
25886: douta=16'h8432;
25887: douta=16'h7bd1;
25888: douta=16'h7bd1;
25889: douta=16'h73b1;
25890: douta=16'h7bd1;
25891: douta=16'h6b0c;
25892: douta=16'h5a69;
25893: douta=16'h2903;
25894: douta=16'h41a6;
25895: douta=16'h62ca;
25896: douta=16'h5a68;
25897: douta=16'h528b;
25898: douta=16'h5b50;
25899: douta=16'h4aef;
25900: douta=16'h29a9;
25901: douta=16'h736f;
25902: douta=16'h31eb;
25903: douta=16'h18e5;
25904: douta=16'h2126;
25905: douta=16'h1905;
25906: douta=16'h59e6;
25907: douta=16'h51e6;
25908: douta=16'h51c6;
25909: douta=16'h49c6;
25910: douta=16'h49a6;
25911: douta=16'h49a5;
25912: douta=16'h49a6;
25913: douta=16'h4186;
25914: douta=16'h4185;
25915: douta=16'h4186;
25916: douta=16'h3966;
25917: douta=16'h3966;
25918: douta=16'h3965;
25919: douta=16'h4166;
25920: douta=16'hffbc;
25921: douta=16'hfffd;
25922: douta=16'hde16;
25923: douta=16'hee77;
25924: douta=16'ha4f5;
25925: douta=16'ha493;
25926: douta=16'hbd55;
25927: douta=16'hcdd6;
25928: douta=16'hbd75;
25929: douta=16'hbd55;
25930: douta=16'h8c53;
25931: douta=16'h9494;
25932: douta=16'h8c94;
25933: douta=16'h8474;
25934: douta=16'h8434;
25935: douta=16'h8454;
25936: douta=16'h8475;
25937: douta=16'h8c74;
25938: douta=16'h6bb1;
25939: douta=16'h18c3;
25940: douta=16'h18a2;
25941: douta=16'h18a3;
25942: douta=16'h20c3;
25943: douta=16'h1082;
25944: douta=16'h1882;
25945: douta=16'h1882;
25946: douta=16'h1882;
25947: douta=16'h1881;
25948: douta=16'h18a2;
25949: douta=16'h2082;
25950: douta=16'h20a2;
25951: douta=16'h20a2;
25952: douta=16'h28c2;
25953: douta=16'h20c2;
25954: douta=16'h28c2;
25955: douta=16'h28e2;
25956: douta=16'h28e2;
25957: douta=16'h3146;
25958: douta=16'h2967;
25959: douta=16'h18a5;
25960: douta=16'h4143;
25961: douta=16'h4143;
25962: douta=16'h4964;
25963: douta=16'h4984;
25964: douta=16'h5184;
25965: douta=16'h51a4;
25966: douta=16'h5183;
25967: douta=16'h9d13;
25968: douta=16'h5983;
25969: douta=16'h4964;
25970: douta=16'h7224;
25971: douta=16'h6a04;
25972: douta=16'h7224;
25973: douta=16'h7224;
25974: douta=16'h7244;
25975: douta=16'h7224;
25976: douta=16'h7224;
25977: douta=16'h7a44;
25978: douta=16'h8285;
25979: douta=16'h8284;
25980: douta=16'h8aa4;
25981: douta=16'h8ac4;
25982: douta=16'h92e4;
25983: douta=16'h9304;
25984: douta=16'h9b05;
25985: douta=16'h9b25;
25986: douta=16'ha325;
25987: douta=16'hab64;
25988: douta=16'hab65;
25989: douta=16'hab85;
25990: douta=16'hb385;
25991: douta=16'hb3a5;
25992: douta=16'hb3c5;
25993: douta=16'hbbe6;
25994: douta=16'hbbe5;
25995: douta=16'hbbe5;
25996: douta=16'hbbe5;
25997: douta=16'hbc06;
25998: douta=16'hbbe5;
25999: douta=16'hc405;
26000: douta=16'hc426;
26001: douta=16'hc426;
26002: douta=16'hc426;
26003: douta=16'hc425;
26004: douta=16'hc425;
26005: douta=16'hc405;
26006: douta=16'hc425;
26007: douta=16'hcc26;
26008: douta=16'hcc26;
26009: douta=16'hcc26;
26010: douta=16'hcc46;
26011: douta=16'hcc46;
26012: douta=16'hcc46;
26013: douta=16'hcc46;
26014: douta=16'hcc46;
26015: douta=16'hcc46;
26016: douta=16'hd467;
26017: douta=16'hd467;
26018: douta=16'hd467;
26019: douta=16'hd467;
26020: douta=16'hd466;
26021: douta=16'hcc47;
26022: douta=16'hd467;
26023: douta=16'hcc66;
26024: douta=16'hd466;
26025: douta=16'hd467;
26026: douta=16'hd467;
26027: douta=16'hd467;
26028: douta=16'hd468;
26029: douta=16'hd467;
26030: douta=16'hd467;
26031: douta=16'hd467;
26032: douta=16'hd467;
26033: douta=16'hd467;
26034: douta=16'hd467;
26035: douta=16'hd467;
26036: douta=16'hd467;
26037: douta=16'hd467;
26038: douta=16'hd467;
26039: douta=16'hd467;
26040: douta=16'hd467;
26041: douta=16'hd468;
26042: douta=16'hb4ad;
26043: douta=16'hce56;
26044: douta=16'h8c31;
26045: douta=16'h8bef;
26046: douta=16'h838f;
26047: douta=16'h6b4e;
26048: douta=16'h734e;
26049: douta=16'h6b4d;
26050: douta=16'h41c6;
26051: douta=16'h5248;
26052: douta=16'h6b2c;
26053: douta=16'hd615;
26054: douta=16'hde14;
26055: douta=16'h8bac;
26056: douta=16'hbd11;
26057: douta=16'hcd71;
26058: douta=16'hcdb2;
26059: douta=16'hc5b3;
26060: douta=16'hcdd4;
26061: douta=16'he697;
26062: douta=16'hcdb3;
26063: douta=16'he676;
26064: douta=16'hde15;
26065: douta=16'hde15;
26066: douta=16'hd5d4;
26067: douta=16'hbd74;
26068: douta=16'hc574;
26069: douta=16'ha4b3;
26070: douta=16'hbd75;
26071: douta=16'h94b3;
26072: douta=16'ha4b4;
26073: douta=16'h9cb4;
26074: douta=16'ha4d5;
26075: douta=16'ha4d5;
26076: douta=16'h9cb4;
26077: douta=16'h8c52;
26078: douta=16'h8412;
26079: douta=16'h73b0;
26080: douta=16'h6b6f;
26081: douta=16'h732e;
26082: douta=16'h6b2d;
26083: douta=16'h2903;
26084: douta=16'h2103;
26085: douta=16'h49e6;
26086: douta=16'h62ea;
26087: douta=16'h736c;
26088: douta=16'h83ad;
26089: douta=16'h6b6f;
26090: douta=16'h5b30;
26091: douta=16'h52ef;
26092: douta=16'h2989;
26093: douta=16'h6b2e;
26094: douta=16'h530f;
26095: douta=16'h10a3;
26096: douta=16'h1925;
26097: douta=16'h1906;
26098: douta=16'h51e6;
26099: douta=16'h51c6;
26100: douta=16'h51c5;
26101: douta=16'h49c6;
26102: douta=16'h49a6;
26103: douta=16'h49a5;
26104: douta=16'h49a6;
26105: douta=16'h4185;
26106: douta=16'h4185;
26107: douta=16'h4165;
26108: douta=16'h4186;
26109: douta=16'h4165;
26110: douta=16'h4165;
26111: douta=16'h3966;
26112: douta=16'hffbd;
26113: douta=16'hff7c;
26114: douta=16'hde36;
26115: douta=16'he677;
26116: douta=16'ha4b4;
26117: douta=16'h9c93;
26118: douta=16'had35;
26119: douta=16'hc5b5;
26120: douta=16'hbd55;
26121: douta=16'hbd75;
26122: douta=16'h94b5;
26123: douta=16'h94b5;
26124: douta=16'h8c94;
26125: douta=16'h8454;
26126: douta=16'h8454;
26127: douta=16'h7c13;
26128: douta=16'h8474;
26129: douta=16'h9d58;
26130: douta=16'h0800;
26131: douta=16'h20c3;
26132: douta=16'h18a3;
26133: douta=16'h18c3;
26134: douta=16'h20e3;
26135: douta=16'h1861;
26136: douta=16'h1882;
26137: douta=16'h1882;
26138: douta=16'h1881;
26139: douta=16'h18a2;
26140: douta=16'h2082;
26141: douta=16'h1881;
26142: douta=16'h2082;
26143: douta=16'h20a2;
26144: douta=16'h20a2;
26145: douta=16'h28c2;
26146: douta=16'h30e2;
26147: douta=16'h30e3;
26148: douta=16'h30e2;
26149: douta=16'h39e9;
26150: douta=16'h2126;
26151: douta=16'h18c4;
26152: douta=16'h4143;
26153: douta=16'h4963;
26154: douta=16'h4963;
26155: douta=16'h5184;
26156: douta=16'h51a4;
26157: douta=16'h51a4;
26158: douta=16'h6267;
26159: douta=16'h9c6f;
26160: douta=16'h69e4;
26161: douta=16'h4984;
26162: douta=16'h61c4;
26163: douta=16'h7224;
26164: douta=16'h7224;
26165: douta=16'h7a44;
26166: douta=16'h7244;
26167: douta=16'h7a44;
26168: douta=16'h7244;
26169: douta=16'h7a64;
26170: douta=16'h8284;
26171: douta=16'h82a4;
26172: douta=16'h8aa4;
26173: douta=16'h8ac5;
26174: douta=16'h92e4;
26175: douta=16'h9305;
26176: douta=16'h9b05;
26177: douta=16'h9b25;
26178: douta=16'ha345;
26179: douta=16'hab64;
26180: douta=16'hab85;
26181: douta=16'hb385;
26182: douta=16'hb385;
26183: douta=16'hb3a5;
26184: douta=16'hbbc6;
26185: douta=16'hbbe6;
26186: douta=16'hbbe6;
26187: douta=16'hbbe5;
26188: douta=16'hbbe5;
26189: douta=16'hbc06;
26190: douta=16'hc406;
26191: douta=16'hc406;
26192: douta=16'hc426;
26193: douta=16'hc426;
26194: douta=16'hcc26;
26195: douta=16'hc426;
26196: douta=16'hcc26;
26197: douta=16'hcc26;
26198: douta=16'hcc26;
26199: douta=16'hcc46;
26200: douta=16'hcc46;
26201: douta=16'hcc26;
26202: douta=16'hcc46;
26203: douta=16'hcc46;
26204: douta=16'hcc46;
26205: douta=16'hcc46;
26206: douta=16'hcc46;
26207: douta=16'hcc47;
26208: douta=16'hd467;
26209: douta=16'hd467;
26210: douta=16'hd467;
26211: douta=16'hd467;
26212: douta=16'hcc66;
26213: douta=16'hd467;
26214: douta=16'hcc47;
26215: douta=16'hd467;
26216: douta=16'hcc67;
26217: douta=16'hd466;
26218: douta=16'hd467;
26219: douta=16'hd487;
26220: douta=16'hd467;
26221: douta=16'hd488;
26222: douta=16'hd467;
26223: douta=16'hd467;
26224: douta=16'hd467;
26225: douta=16'hd467;
26226: douta=16'hcc67;
26227: douta=16'hd487;
26228: douta=16'hd487;
26229: douta=16'hd487;
26230: douta=16'hd467;
26231: douta=16'hd468;
26232: douta=16'hd488;
26233: douta=16'hd468;
26234: douta=16'hbccd;
26235: douta=16'hce56;
26236: douta=16'hdc86;
26237: douta=16'hcc89;
26238: douta=16'h6b2d;
26239: douta=16'h6aeb;
26240: douta=16'h7b8d;
26241: douta=16'hb4f2;
26242: douta=16'h8c2e;
26243: douta=16'hacd2;
26244: douta=16'hacf2;
26245: douta=16'ha490;
26246: douta=16'ha48f;
26247: douta=16'hde15;
26248: douta=16'hd5f5;
26249: douta=16'hd614;
26250: douta=16'hde15;
26251: douta=16'hd5f4;
26252: douta=16'hde36;
26253: douta=16'hde16;
26254: douta=16'hbd33;
26255: douta=16'hacf3;
26256: douta=16'hc594;
26257: douta=16'hb535;
26258: douta=16'ha4f5;
26259: douta=16'h9cb4;
26260: douta=16'h9cb4;
26261: douta=16'h9cb4;
26262: douta=16'h94b4;
26263: douta=16'h7c12;
26264: douta=16'h8433;
26265: douta=16'h8452;
26266: douta=16'h8432;
26267: douta=16'h8412;
26268: douta=16'h7bf1;
26269: douta=16'h7baf;
26270: douta=16'h5aaa;
26271: douta=16'h41a5;
26272: douta=16'h0000;
26273: douta=16'h5aa8;
26274: douta=16'h5aa8;
26275: douta=16'h6aeb;
26276: douta=16'h6acb;
26277: douta=16'h732b;
26278: douta=16'h838d;
26279: douta=16'h8bce;
26280: douta=16'h9c90;
26281: douta=16'h2127;
26282: douta=16'h18e5;
26283: douta=16'h10c4;
26284: douta=16'h10a4;
26285: douta=16'h39a6;
26286: douta=16'h08a3;
26287: douta=16'h2167;
26288: douta=16'h2167;
26289: douta=16'h08a4;
26290: douta=16'h51e6;
26291: douta=16'h51c6;
26292: douta=16'h49c6;
26293: douta=16'h49c6;
26294: douta=16'h49a6;
26295: douta=16'h49a6;
26296: douta=16'h4186;
26297: douta=16'h49a6;
26298: douta=16'h4185;
26299: douta=16'h4185;
26300: douta=16'h4185;
26301: douta=16'h4186;
26302: douta=16'h4186;
26303: douta=16'h4186;
26304: douta=16'hffbd;
26305: douta=16'hde16;
26306: douta=16'he698;
26307: douta=16'hd5f6;
26308: douta=16'h9c93;
26309: douta=16'had15;
26310: douta=16'hb515;
26311: douta=16'hc595;
26312: douta=16'hbd55;
26313: douta=16'hb576;
26314: douta=16'h94b5;
26315: douta=16'h9494;
26316: douta=16'h8c74;
26317: douta=16'h8454;
26318: douta=16'h8434;
26319: douta=16'h8454;
26320: douta=16'h8c74;
26321: douta=16'h73f2;
26322: douta=16'h20a2;
26323: douta=16'h20a3;
26324: douta=16'h20c3;
26325: douta=16'h18a3;
26326: douta=16'h18c3;
26327: douta=16'h1882;
26328: douta=16'h1882;
26329: douta=16'h1882;
26330: douta=16'h18a2;
26331: douta=16'h2082;
26332: douta=16'h20a2;
26333: douta=16'h20a2;
26334: douta=16'h20a2;
26335: douta=16'h20a2;
26336: douta=16'h20c2;
26337: douta=16'h28e2;
26338: douta=16'h28e2;
26339: douta=16'h28e2;
26340: douta=16'h3103;
26341: douta=16'h31c9;
26342: douta=16'h18e5;
26343: douta=16'h28e3;
26344: douta=16'h4163;
26345: douta=16'h4963;
26346: douta=16'h4984;
26347: douta=16'h5184;
26348: douta=16'h59a4;
26349: douta=16'h51a4;
26350: douta=16'h6aeb;
26351: douta=16'h8bec;
26352: douta=16'h6a04;
26353: douta=16'h4984;
26354: douta=16'h59a4;
26355: douta=16'h7224;
26356: douta=16'h7244;
26357: douta=16'h7a64;
26358: douta=16'h7a64;
26359: douta=16'h7244;
26360: douta=16'h7a44;
26361: douta=16'h7a64;
26362: douta=16'h8285;
26363: douta=16'h82a5;
26364: douta=16'h8aa4;
26365: douta=16'h8ae4;
26366: douta=16'h9304;
26367: douta=16'h9b05;
26368: douta=16'h9b25;
26369: douta=16'ha325;
26370: douta=16'ha345;
26371: douta=16'hab65;
26372: douta=16'hab85;
26373: douta=16'hab85;
26374: douta=16'hb3a5;
26375: douta=16'hb3a6;
26376: douta=16'hb3a6;
26377: douta=16'hbbe6;
26378: douta=16'hbbe6;
26379: douta=16'hbbe5;
26380: douta=16'hc406;
26381: douta=16'hbc06;
26382: douta=16'hbc06;
26383: douta=16'hc405;
26384: douta=16'hc406;
26385: douta=16'hc426;
26386: douta=16'hc426;
26387: douta=16'hcc47;
26388: douta=16'hcc46;
26389: douta=16'hc426;
26390: douta=16'hcc46;
26391: douta=16'hcc46;
26392: douta=16'hcc47;
26393: douta=16'hcc47;
26394: douta=16'hcc46;
26395: douta=16'hcc46;
26396: douta=16'hcc46;
26397: douta=16'hcc46;
26398: douta=16'hcc47;
26399: douta=16'hcc46;
26400: douta=16'hcc47;
26401: douta=16'hd467;
26402: douta=16'hd467;
26403: douta=16'hd467;
26404: douta=16'hd467;
26405: douta=16'hcc67;
26406: douta=16'hd467;
26407: douta=16'hd467;
26408: douta=16'hd467;
26409: douta=16'hcc67;
26410: douta=16'hcc67;
26411: douta=16'hd467;
26412: douta=16'hd467;
26413: douta=16'hd467;
26414: douta=16'hd467;
26415: douta=16'hd487;
26416: douta=16'hd487;
26417: douta=16'hd487;
26418: douta=16'hd487;
26419: douta=16'hd467;
26420: douta=16'hd467;
26421: douta=16'hd488;
26422: douta=16'hd467;
26423: douta=16'hd487;
26424: douta=16'hd468;
26425: douta=16'hd468;
26426: douta=16'hbcce;
26427: douta=16'hce77;
26428: douta=16'hcc87;
26429: douta=16'hd486;
26430: douta=16'h9430;
26431: douta=16'h7b6c;
26432: douta=16'h9c2e;
26433: douta=16'h734a;
26434: douta=16'hbd52;
26435: douta=16'hbd73;
26436: douta=16'hcdf5;
26437: douta=16'h9c8f;
26438: douta=16'hcdd6;
26439: douta=16'hd615;
26440: douta=16'hd5d4;
26441: douta=16'hd5f4;
26442: douta=16'hd5f4;
26443: douta=16'hcdd3;
26444: douta=16'hbd33;
26445: douta=16'hb514;
26446: douta=16'hb533;
26447: douta=16'hb513;
26448: douta=16'ha4d3;
26449: douta=16'h9cd4;
26450: douta=16'h9cb4;
26451: douta=16'h8c53;
26452: douta=16'h8c73;
26453: douta=16'h8c73;
26454: douta=16'h8412;
26455: douta=16'h8c53;
26456: douta=16'h7bb0;
26457: douta=16'h83d1;
26458: douta=16'h736d;
26459: douta=16'h51e6;
26460: douta=16'h49c4;
26461: douta=16'h41a5;
26462: douta=16'h5226;
26463: douta=16'h5a89;
26464: douta=16'h734b;
26465: douta=16'h62c9;
26466: douta=16'h6b0b;
26467: douta=16'h83cd;
26468: douta=16'h83cd;
26469: douta=16'h8bee;
26470: douta=16'h944f;
26471: douta=16'h9c4f;
26472: douta=16'hacf2;
26473: douta=16'h5acc;
26474: douta=16'h2967;
26475: douta=16'h1104;
26476: douta=16'h10c3;
26477: douta=16'h0883;
26478: douta=16'h39a7;
26479: douta=16'h1084;
26480: douta=16'h2126;
26481: douta=16'h2947;
26482: douta=16'h51a5;
26483: douta=16'h51c6;
26484: douta=16'h49a6;
26485: douta=16'h49a6;
26486: douta=16'h4986;
26487: douta=16'h4986;
26488: douta=16'h49a6;
26489: douta=16'h4185;
26490: douta=16'h4185;
26491: douta=16'h4185;
26492: douta=16'h4186;
26493: douta=16'h4166;
26494: douta=16'h4165;
26495: douta=16'h4186;
26496: douta=16'hffbd;
26497: douta=16'hd5b5;
26498: douta=16'he678;
26499: douta=16'hc5b6;
26500: douta=16'ha4b3;
26501: douta=16'hb535;
26502: douta=16'hb535;
26503: douta=16'hbd75;
26504: douta=16'hbd55;
26505: douta=16'had56;
26506: douta=16'h94b5;
26507: douta=16'h8c74;
26508: douta=16'h8c95;
26509: douta=16'h8474;
26510: douta=16'h8454;
26511: douta=16'h8474;
26512: douta=16'h8c75;
26513: douta=16'h4acd;
26514: douta=16'h20a3;
26515: douta=16'h20c3;
26516: douta=16'h20a3;
26517: douta=16'h20c2;
26518: douta=16'h18a2;
26519: douta=16'h1882;
26520: douta=16'h1882;
26521: douta=16'h1882;
26522: douta=16'h1881;
26523: douta=16'h2082;
26524: douta=16'h20a2;
26525: douta=16'h20a2;
26526: douta=16'h2082;
26527: douta=16'h20a2;
26528: douta=16'h28c2;
26529: douta=16'h28e2;
26530: douta=16'h30e3;
26531: douta=16'h28e2;
26532: douta=16'h30e2;
26533: douta=16'h31c9;
26534: douta=16'h18c5;
26535: douta=16'h28e3;
26536: douta=16'h4963;
26537: douta=16'h4963;
26538: douta=16'h4964;
26539: douta=16'h51a4;
26540: douta=16'h51a4;
26541: douta=16'h59c4;
26542: douta=16'h734d;
26543: douta=16'h836a;
26544: douta=16'h6a04;
26545: douta=16'h4984;
26546: douta=16'h59c4;
26547: douta=16'h7224;
26548: douta=16'h7224;
26549: douta=16'h7244;
26550: douta=16'h7244;
26551: douta=16'h7a44;
26552: douta=16'h7a44;
26553: douta=16'h7a64;
26554: douta=16'h8284;
26555: douta=16'h82a5;
26556: douta=16'h8aa4;
26557: douta=16'h8ac5;
26558: douta=16'h9305;
26559: douta=16'h9b05;
26560: douta=16'h9b45;
26561: douta=16'h9b25;
26562: douta=16'ha365;
26563: douta=16'hab65;
26564: douta=16'hab85;
26565: douta=16'haba5;
26566: douta=16'hb385;
26567: douta=16'hb3a5;
26568: douta=16'hbbc6;
26569: douta=16'hbbe6;
26570: douta=16'hbbe6;
26571: douta=16'hbbe6;
26572: douta=16'hbbe5;
26573: douta=16'hc406;
26574: douta=16'hc406;
26575: douta=16'hc426;
26576: douta=16'hc406;
26577: douta=16'hc426;
26578: douta=16'hc426;
26579: douta=16'hcc26;
26580: douta=16'hc426;
26581: douta=16'hcc26;
26582: douta=16'hcc26;
26583: douta=16'hcc46;
26584: douta=16'hcc47;
26585: douta=16'hcc47;
26586: douta=16'hcc46;
26587: douta=16'hcc46;
26588: douta=16'hcc46;
26589: douta=16'hcc47;
26590: douta=16'hcc47;
26591: douta=16'hcc47;
26592: douta=16'hcc46;
26593: douta=16'hcc47;
26594: douta=16'hcc47;
26595: douta=16'hcc67;
26596: douta=16'hd467;
26597: douta=16'hcc47;
26598: douta=16'hd467;
26599: douta=16'hd467;
26600: douta=16'hd467;
26601: douta=16'hcc67;
26602: douta=16'hd467;
26603: douta=16'hd467;
26604: douta=16'hd468;
26605: douta=16'hd487;
26606: douta=16'hd487;
26607: douta=16'hd467;
26608: douta=16'hd467;
26609: douta=16'hd487;
26610: douta=16'hd487;
26611: douta=16'hd467;
26612: douta=16'hd467;
26613: douta=16'hd488;
26614: douta=16'hd467;
26615: douta=16'hd487;
26616: douta=16'hd488;
26617: douta=16'hd468;
26618: douta=16'hbcce;
26619: douta=16'hce77;
26620: douta=16'hd487;
26621: douta=16'hd489;
26622: douta=16'hac2b;
26623: douta=16'h836d;
26624: douta=16'hbd53;
26625: douta=16'h838d;
26626: douta=16'hbd72;
26627: douta=16'hcdb4;
26628: douta=16'hde36;
26629: douta=16'had11;
26630: douta=16'he636;
26631: douta=16'hd5f5;
26632: douta=16'hd5d5;
26633: douta=16'hcd73;
26634: douta=16'hd5d4;
26635: douta=16'hc533;
26636: douta=16'hacf3;
26637: douta=16'hacd3;
26638: douta=16'hacd3;
26639: douta=16'hacf3;
26640: douta=16'ha4d3;
26641: douta=16'h8c74;
26642: douta=16'h8c73;
26643: douta=16'h7c12;
26644: douta=16'h83f2;
26645: douta=16'h8412;
26646: douta=16'h8412;
26647: douta=16'h8411;
26648: douta=16'h6aeb;
26649: douta=16'h6b0c;
26650: douta=16'h3984;
26651: douta=16'h28e2;
26652: douta=16'h5a87;
26653: douta=16'h62a9;
26654: douta=16'h628a;
26655: douta=16'h62ca;
26656: douta=16'h7b8c;
26657: douta=16'h736c;
26658: douta=16'h7b8c;
26659: douta=16'h940e;
26660: douta=16'h9c4e;
26661: douta=16'h942f;
26662: douta=16'ha490;
26663: douta=16'ha490;
26664: douta=16'hacd1;
26665: douta=16'h6b2e;
26666: douta=16'h4a8b;
26667: douta=16'h2127;
26668: douta=16'h1905;
26669: douta=16'h10e3;
26670: douta=16'h18c4;
26671: douta=16'h18c4;
26672: douta=16'h0882;
26673: douta=16'h18e5;
26674: douta=16'h4965;
26675: douta=16'h51c6;
26676: douta=16'h49a6;
26677: douta=16'h49a5;
26678: douta=16'h49a6;
26679: douta=16'h49a6;
26680: douta=16'h49a6;
26681: douta=16'h4186;
26682: douta=16'h4186;
26683: douta=16'h4165;
26684: douta=16'h4165;
26685: douta=16'h4145;
26686: douta=16'h3903;
26687: douta=16'h30e3;
26688: douta=16'hffdd;
26689: douta=16'hd5f6;
26690: douta=16'he677;
26691: douta=16'h9cb3;
26692: douta=16'hb535;
26693: douta=16'had15;
26694: douta=16'hcdf6;
26695: douta=16'hb555;
26696: douta=16'had35;
26697: douta=16'h9494;
26698: douta=16'h8c94;
26699: douta=16'h94b5;
26700: douta=16'h8c95;
26701: douta=16'h8454;
26702: douta=16'h8c74;
26703: douta=16'h8c74;
26704: douta=16'h9517;
26705: douta=16'h1040;
26706: douta=16'h20c3;
26707: douta=16'h20a3;
26708: douta=16'h20a3;
26709: douta=16'h18c3;
26710: douta=16'h1882;
26711: douta=16'h1882;
26712: douta=16'h18a2;
26713: douta=16'h1882;
26714: douta=16'h1882;
26715: douta=16'h20a2;
26716: douta=16'h20a2;
26717: douta=16'h20a2;
26718: douta=16'h20a2;
26719: douta=16'h20a2;
26720: douta=16'h28e3;
26721: douta=16'h28e2;
26722: douta=16'h30e2;
26723: douta=16'h30e3;
26724: douta=16'h30e2;
26725: douta=16'h31a8;
26726: douta=16'h18a4;
26727: douta=16'h4123;
26728: douta=16'h4963;
26729: douta=16'h4984;
26730: douta=16'h4963;
26731: douta=16'h59a4;
26732: douta=16'h59c4;
26733: douta=16'h59c4;
26734: douta=16'h94b2;
26735: douta=16'h6a44;
26736: douta=16'h6a04;
26737: douta=16'h4143;
26738: douta=16'h61c4;
26739: douta=16'h7224;
26740: douta=16'h7a44;
26741: douta=16'h7a64;
26742: douta=16'h7a84;
26743: douta=16'h7a64;
26744: douta=16'h7a44;
26745: douta=16'h7a64;
26746: douta=16'h82a4;
26747: douta=16'h82a4;
26748: douta=16'h8aa4;
26749: douta=16'h92e5;
26750: douta=16'h9304;
26751: douta=16'h9b05;
26752: douta=16'h9b45;
26753: douta=16'ha345;
26754: douta=16'ha365;
26755: douta=16'hab85;
26756: douta=16'hb385;
26757: douta=16'hb385;
26758: douta=16'hb3a5;
26759: douta=16'hbbc6;
26760: douta=16'hbbc6;
26761: douta=16'hbbe6;
26762: douta=16'hbbc6;
26763: douta=16'hbbe6;
26764: douta=16'hbc06;
26765: douta=16'hc406;
26766: douta=16'hc406;
26767: douta=16'hc426;
26768: douta=16'hc426;
26769: douta=16'hc426;
26770: douta=16'hc426;
26771: douta=16'hcc26;
26772: douta=16'hcc46;
26773: douta=16'hcc47;
26774: douta=16'hcc47;
26775: douta=16'hc426;
26776: douta=16'hcc47;
26777: douta=16'hcc46;
26778: douta=16'hcc46;
26779: douta=16'hcc46;
26780: douta=16'hcc46;
26781: douta=16'hcc46;
26782: douta=16'hcc46;
26783: douta=16'hcc46;
26784: douta=16'hcc47;
26785: douta=16'hcc46;
26786: douta=16'hcc47;
26787: douta=16'hcc46;
26788: douta=16'hd467;
26789: douta=16'hd467;
26790: douta=16'hd467;
26791: douta=16'hd467;
26792: douta=16'hd467;
26793: douta=16'hd467;
26794: douta=16'hd467;
26795: douta=16'hcc67;
26796: douta=16'hd467;
26797: douta=16'hd487;
26798: douta=16'hd487;
26799: douta=16'hd487;
26800: douta=16'hd467;
26801: douta=16'hd467;
26802: douta=16'hd467;
26803: douta=16'hd487;
26804: douta=16'hd467;
26805: douta=16'hd487;
26806: douta=16'hd468;
26807: douta=16'hd488;
26808: douta=16'hd488;
26809: douta=16'hd466;
26810: douta=16'hb4ce;
26811: douta=16'hce76;
26812: douta=16'hd468;
26813: douta=16'hcc87;
26814: douta=16'he486;
26815: douta=16'hacd1;
26816: douta=16'hacd1;
26817: douta=16'hb511;
26818: douta=16'hc573;
26819: douta=16'hde37;
26820: douta=16'hd616;
26821: douta=16'hde57;
26822: douta=16'hcdd5;
26823: douta=16'hc596;
26824: douta=16'hbd75;
26825: douta=16'hacf3;
26826: douta=16'h9c93;
26827: douta=16'h9452;
26828: douta=16'h9473;
26829: douta=16'h9473;
26830: douta=16'h8c12;
26831: douta=16'h83f1;
26832: douta=16'h7bb0;
26833: douta=16'h7390;
26834: douta=16'h7bd0;
26835: douta=16'h738e;
26836: douta=16'h41a6;
26837: douta=16'h49a5;
26838: douta=16'h3944;
26839: douta=16'h5227;
26840: douta=16'h5a88;
26841: douta=16'h6288;
26842: douta=16'h7b6b;
26843: douta=16'h6aea;
26844: douta=16'h732a;
26845: douta=16'h83cd;
26846: douta=16'h8c0d;
26847: douta=16'h9c4f;
26848: douta=16'hacf0;
26849: douta=16'hbd31;
26850: douta=16'hbd31;
26851: douta=16'hc551;
26852: douta=16'hc572;
26853: douta=16'hc572;
26854: douta=16'hbd52;
26855: douta=16'hb4d1;
26856: douta=16'ha4b1;
26857: douta=16'h83f0;
26858: douta=16'h6b6f;
26859: douta=16'h5b0e;
26860: douta=16'h39e9;
26861: douta=16'h31a8;
26862: douta=16'h2126;
26863: douta=16'h2106;
26864: douta=16'h2968;
26865: douta=16'h2988;
26866: douta=16'h832c;
26867: douta=16'h51a5;
26868: douta=16'h4a07;
26869: douta=16'h5aab;
26870: douta=16'h6b4e;
26871: douta=16'h6b6f;
26872: douta=16'h7432;
26873: douta=16'h7c73;
26874: douta=16'h7c73;
26875: douta=16'h7c73;
26876: douta=16'h7452;
26877: douta=16'h6bd0;
26878: douta=16'h5b2d;
26879: douta=16'h52cb;
26880: douta=16'hf6f9;
26881: douta=16'hde37;
26882: douta=16'hde37;
26883: douta=16'ha4b3;
26884: douta=16'hacf5;
26885: douta=16'hb514;
26886: douta=16'hcdb5;
26887: douta=16'hb555;
26888: douta=16'h9494;
26889: douta=16'h9cb4;
26890: douta=16'h8c94;
26891: douta=16'h94b5;
26892: douta=16'h8c95;
26893: douta=16'h8433;
26894: douta=16'h8c95;
26895: douta=16'h8475;
26896: douta=16'h3a4a;
26897: douta=16'h20c3;
26898: douta=16'h20c3;
26899: douta=16'h20c3;
26900: douta=16'h20c3;
26901: douta=16'h18a3;
26902: douta=16'h1882;
26903: douta=16'h1882;
26904: douta=16'h1882;
26905: douta=16'h2082;
26906: douta=16'h2082;
26907: douta=16'h20a2;
26908: douta=16'h20a2;
26909: douta=16'h2082;
26910: douta=16'h20a2;
26911: douta=16'h28c2;
26912: douta=16'h28e2;
26913: douta=16'h28c2;
26914: douta=16'h30e3;
26915: douta=16'h30e3;
26916: douta=16'h30e2;
26917: douta=16'h2967;
26918: douta=16'h28e4;
26919: douta=16'h4943;
26920: douta=16'h4963;
26921: douta=16'h4963;
26922: douta=16'h5184;
26923: douta=16'h51a3;
26924: douta=16'h59a4;
26925: douta=16'h61c4;
26926: douta=16'ha555;
26927: douta=16'h61a3;
26928: douta=16'h6a24;
26929: douta=16'h4164;
26930: douta=16'h51a4;
26931: douta=16'h7244;
26932: douta=16'h7a44;
26933: douta=16'h7a64;
26934: douta=16'h7a64;
26935: douta=16'h7a64;
26936: douta=16'h7a84;
26937: douta=16'h7a64;
26938: douta=16'h82a4;
26939: douta=16'h8ac5;
26940: douta=16'h8ac4;
26941: douta=16'h92e5;
26942: douta=16'h9305;
26943: douta=16'h9b25;
26944: douta=16'ha346;
26945: douta=16'ha345;
26946: douta=16'ha365;
26947: douta=16'hab65;
26948: douta=16'hb3a5;
26949: douta=16'hb3a5;
26950: douta=16'hb3a5;
26951: douta=16'hbbc5;
26952: douta=16'hbbc5;
26953: douta=16'hbbc6;
26954: douta=16'hbbe6;
26955: douta=16'hbc06;
26956: douta=16'hc406;
26957: douta=16'hc406;
26958: douta=16'hc406;
26959: douta=16'hc426;
26960: douta=16'hc426;
26961: douta=16'hc426;
26962: douta=16'hc426;
26963: douta=16'hcc26;
26964: douta=16'hcc46;
26965: douta=16'hcc26;
26966: douta=16'hcc46;
26967: douta=16'hcc46;
26968: douta=16'hcc26;
26969: douta=16'hcc46;
26970: douta=16'hcc46;
26971: douta=16'hcc46;
26972: douta=16'hcc46;
26973: douta=16'hcc46;
26974: douta=16'hcc46;
26975: douta=16'hcc47;
26976: douta=16'hcc46;
26977: douta=16'hcc47;
26978: douta=16'hcc46;
26979: douta=16'hcc47;
26980: douta=16'hd467;
26981: douta=16'hd467;
26982: douta=16'hd467;
26983: douta=16'hd467;
26984: douta=16'hcc67;
26985: douta=16'hd467;
26986: douta=16'hcc47;
26987: douta=16'hd468;
26988: douta=16'hd468;
26989: douta=16'hd487;
26990: douta=16'hd467;
26991: douta=16'hd487;
26992: douta=16'hd467;
26993: douta=16'hd467;
26994: douta=16'hd487;
26995: douta=16'hd487;
26996: douta=16'hd487;
26997: douta=16'hd467;
26998: douta=16'hd487;
26999: douta=16'hd488;
27000: douta=16'hd488;
27001: douta=16'hd467;
27002: douta=16'hb4ce;
27003: douta=16'hce76;
27004: douta=16'hd488;
27005: douta=16'hd487;
27006: douta=16'hd467;
27007: douta=16'h944f;
27008: douta=16'ha4b1;
27009: douta=16'hacd1;
27010: douta=16'hc594;
27011: douta=16'hcdf5;
27012: douta=16'hc5b5;
27013: douta=16'hc5b6;
27014: douta=16'hbd96;
27015: douta=16'hb556;
27016: douta=16'ha4f5;
27017: douta=16'h9493;
27018: douta=16'h9c94;
27019: douta=16'h7bf1;
27020: douta=16'h83f1;
27021: douta=16'h83f0;
27022: douta=16'h7bd0;
27023: douta=16'h83f0;
27024: douta=16'h734d;
27025: douta=16'h4a27;
27026: douta=16'h2903;
27027: douta=16'h3123;
27028: douta=16'h732b;
27029: douta=16'h62ca;
27030: douta=16'h6aea;
27031: douta=16'h730a;
27032: douta=16'h730a;
27033: douta=16'h732a;
27034: douta=16'h8bee;
27035: douta=16'h8c0e;
27036: douta=16'h942e;
27037: douta=16'h9c8f;
27038: douta=16'h9c6f;
27039: douta=16'ha4af;
27040: douta=16'hbd51;
27041: douta=16'hc572;
27042: douta=16'hc572;
27043: douta=16'hcdb3;
27044: douta=16'hd5d4;
27045: douta=16'hcdb3;
27046: douta=16'hc573;
27047: douta=16'hacd2;
27048: douta=16'ha4b1;
27049: douta=16'h8410;
27050: douta=16'h632e;
27051: douta=16'h5aec;
27052: douta=16'h4aad;
27053: douta=16'h426c;
27054: douta=16'h31c9;
27055: douta=16'h2126;
27056: douta=16'h1905;
27057: douta=16'h2126;
27058: douta=16'h0062;
27059: douta=16'h10e5;
27060: douta=16'h52ab;
27061: douta=16'h6b6e;
27062: douta=16'h632c;
27063: douta=16'h5acb;
27064: douta=16'h5289;
27065: douta=16'h5228;
27066: douta=16'h49e7;
27067: douta=16'h49a5;
27068: douta=16'h4985;
27069: douta=16'h4965;
27070: douta=16'h4985;
27071: douta=16'h5185;
27072: douta=16'he697;
27073: douta=16'hde77;
27074: douta=16'hcdd6;
27075: douta=16'ha4d4;
27076: douta=16'hacf5;
27077: douta=16'hc595;
27078: douta=16'hc595;
27079: douta=16'hb555;
27080: douta=16'h9453;
27081: douta=16'h9cd5;
27082: douta=16'h8c74;
27083: douta=16'h94b5;
27084: douta=16'h8c74;
27085: douta=16'h8433;
27086: douta=16'h8475;
27087: douta=16'h8c74;
27088: douta=16'h18a2;
27089: douta=16'h20c3;
27090: douta=16'h20c3;
27091: douta=16'h20c3;
27092: douta=16'h20c3;
27093: douta=16'h18a3;
27094: douta=16'h1882;
27095: douta=16'h1882;
27096: douta=16'h1882;
27097: douta=16'h2082;
27098: douta=16'h2082;
27099: douta=16'h20a2;
27100: douta=16'h20a2;
27101: douta=16'h20a2;
27102: douta=16'h20c2;
27103: douta=16'h20c2;
27104: douta=16'h20c2;
27105: douta=16'h28e2;
27106: douta=16'h30e3;
27107: douta=16'h3103;
27108: douta=16'h3103;
27109: douta=16'h2947;
27110: douta=16'h3103;
27111: douta=16'h4963;
27112: douta=16'h4963;
27113: douta=16'h4963;
27114: douta=16'h5184;
27115: douta=16'h51a4;
27116: douta=16'h59c4;
27117: douta=16'h61c4;
27118: douta=16'had74;
27119: douta=16'h61a3;
27120: douta=16'h6a04;
27121: douta=16'h4964;
27122: douta=16'h5184;
27123: douta=16'h7224;
27124: douta=16'h7a44;
27125: douta=16'h7a64;
27126: douta=16'h7a85;
27127: douta=16'h7a44;
27128: douta=16'h7a64;
27129: douta=16'h7a64;
27130: douta=16'h82a4;
27131: douta=16'h8ac4;
27132: douta=16'h8ac4;
27133: douta=16'h92e5;
27134: douta=16'h9305;
27135: douta=16'h9b26;
27136: douta=16'ha346;
27137: douta=16'ha345;
27138: douta=16'hab65;
27139: douta=16'hab85;
27140: douta=16'hb3a5;
27141: douta=16'hb3a5;
27142: douta=16'hb3a6;
27143: douta=16'hbbc5;
27144: douta=16'hbbc5;
27145: douta=16'hbbe6;
27146: douta=16'hbbe6;
27147: douta=16'hbbe5;
27148: douta=16'hc406;
27149: douta=16'hc406;
27150: douta=16'hc406;
27151: douta=16'hc426;
27152: douta=16'hc426;
27153: douta=16'hc426;
27154: douta=16'hcc26;
27155: douta=16'hcc26;
27156: douta=16'hcc46;
27157: douta=16'hcc26;
27158: douta=16'hcc47;
27159: douta=16'hcc26;
27160: douta=16'hcc46;
27161: douta=16'hcc46;
27162: douta=16'hcc46;
27163: douta=16'hcc46;
27164: douta=16'hcc46;
27165: douta=16'hcc46;
27166: douta=16'hcc46;
27167: douta=16'hcc46;
27168: douta=16'hcc67;
27169: douta=16'hcc47;
27170: douta=16'hcc47;
27171: douta=16'hcc67;
27172: douta=16'hd467;
27173: douta=16'hd467;
27174: douta=16'hd467;
27175: douta=16'hd467;
27176: douta=16'hd467;
27177: douta=16'hcc67;
27178: douta=16'hd467;
27179: douta=16'hd468;
27180: douta=16'hd488;
27181: douta=16'hd487;
27182: douta=16'hd467;
27183: douta=16'hd467;
27184: douta=16'hd467;
27185: douta=16'hd487;
27186: douta=16'hd487;
27187: douta=16'hd467;
27188: douta=16'hd487;
27189: douta=16'hd467;
27190: douta=16'hd468;
27191: douta=16'hd488;
27192: douta=16'hd488;
27193: douta=16'hd467;
27194: douta=16'hb4ce;
27195: douta=16'hce56;
27196: douta=16'hd488;
27197: douta=16'hd487;
27198: douta=16'hd487;
27199: douta=16'h9430;
27200: douta=16'ha491;
27201: douta=16'ha472;
27202: douta=16'hc553;
27203: douta=16'hc5b5;
27204: douta=16'hc595;
27205: douta=16'hb575;
27206: douta=16'had36;
27207: douta=16'had56;
27208: douta=16'h9cd4;
27209: douta=16'h8433;
27210: douta=16'h8433;
27211: douta=16'h7b90;
27212: douta=16'h83d0;
27213: douta=16'h7b8f;
27214: douta=16'h7b6e;
27215: douta=16'h6aeb;
27216: douta=16'h49e5;
27217: douta=16'h4185;
27218: douta=16'h5247;
27219: douta=16'h5a88;
27220: douta=16'h9c6f;
27221: douta=16'h838c;
27222: douta=16'h730b;
27223: douta=16'h7b4b;
27224: douta=16'h836b;
27225: douta=16'h834b;
27226: douta=16'h940e;
27227: douta=16'h9c6f;
27228: douta=16'hacd0;
27229: douta=16'hacd0;
27230: douta=16'hacaf;
27231: douta=16'hb510;
27232: douta=16'hcdb3;
27233: douta=16'hcdb3;
27234: douta=16'hcdb3;
27235: douta=16'hcdb4;
27236: douta=16'hcdd4;
27237: douta=16'hcdb3;
27238: douta=16'hcd93;
27239: douta=16'hb512;
27240: douta=16'hacd2;
27241: douta=16'h8c30;
27242: douta=16'h6b6f;
27243: douta=16'h5b0d;
27244: douta=16'h52cd;
27245: douta=16'h4a8d;
27246: douta=16'h3a4c;
27247: douta=16'h2967;
27248: douta=16'h10a4;
27249: douta=16'h1905;
27250: douta=16'h1083;
27251: douta=16'h18e5;
27252: douta=16'h2925;
27253: douta=16'h5226;
27254: douta=16'h49c6;
27255: douta=16'h49a5;
27256: douta=16'h4985;
27257: douta=16'h4985;
27258: douta=16'h4985;
27259: douta=16'h4985;
27260: douta=16'h49a5;
27261: douta=16'h51a5;
27262: douta=16'h51c5;
27263: douta=16'h49a5;
27264: douta=16'hcdb5;
27265: douta=16'he677;
27266: douta=16'hacd4;
27267: douta=16'ha4b3;
27268: douta=16'hcdd5;
27269: douta=16'hd5d6;
27270: douta=16'hb555;
27271: douta=16'ha4f5;
27272: douta=16'h9c94;
27273: douta=16'h9493;
27274: douta=16'h8c94;
27275: douta=16'h9495;
27276: douta=16'h8c94;
27277: douta=16'h8454;
27278: douta=16'h8c95;
27279: douta=16'ha558;
27280: douta=16'h20c3;
27281: douta=16'h20a3;
27282: douta=16'h20c3;
27283: douta=16'h20c3;
27284: douta=16'h18c3;
27285: douta=16'h20c3;
27286: douta=16'h1882;
27287: douta=16'h1881;
27288: douta=16'h1881;
27289: douta=16'h20a2;
27290: douta=16'h20a2;
27291: douta=16'h20a2;
27292: douta=16'h20a2;
27293: douta=16'h20c2;
27294: douta=16'h20a2;
27295: douta=16'h28c2;
27296: douta=16'h28e2;
27297: douta=16'h30e3;
27298: douta=16'h3103;
27299: douta=16'h3903;
27300: douta=16'h3144;
27301: douta=16'h1905;
27302: douta=16'h4143;
27303: douta=16'h4963;
27304: douta=16'h4983;
27305: douta=16'h51a4;
27306: douta=16'h5184;
27307: douta=16'h51a4;
27308: douta=16'h59c4;
27309: douta=16'h5983;
27310: douta=16'h9cb0;
27311: douta=16'h6a03;
27312: douta=16'h6a24;
27313: douta=16'h7264;
27314: douta=16'h49a4;
27315: douta=16'h7a83;
27316: douta=16'h7a64;
27317: douta=16'h7a64;
27318: douta=16'h7a84;
27319: douta=16'h7a84;
27320: douta=16'h7a64;
27321: douta=16'h8284;
27322: douta=16'h8284;
27323: douta=16'h8aa4;
27324: douta=16'h8ac5;
27325: douta=16'h92e4;
27326: douta=16'h9325;
27327: douta=16'h9b45;
27328: douta=16'ha366;
27329: douta=16'ha345;
27330: douta=16'hab65;
27331: douta=16'hb385;
27332: douta=16'hb3a6;
27333: douta=16'hb3a5;
27334: douta=16'hb3a6;
27335: douta=16'hbbc5;
27336: douta=16'hbbe6;
27337: douta=16'hbbe6;
27338: douta=16'hbbe6;
27339: douta=16'hbbe5;
27340: douta=16'hc406;
27341: douta=16'hc407;
27342: douta=16'hc407;
27343: douta=16'hc406;
27344: douta=16'hc426;
27345: douta=16'hc426;
27346: douta=16'hc426;
27347: douta=16'hc426;
27348: douta=16'hc426;
27349: douta=16'hcc46;
27350: douta=16'hcc26;
27351: douta=16'hcc26;
27352: douta=16'hcc46;
27353: douta=16'hcc46;
27354: douta=16'hcc46;
27355: douta=16'hcc46;
27356: douta=16'hcc47;
27357: douta=16'hcc47;
27358: douta=16'hcc47;
27359: douta=16'hcc67;
27360: douta=16'hcc46;
27361: douta=16'hcc47;
27362: douta=16'hd467;
27363: douta=16'hcc47;
27364: douta=16'hd467;
27365: douta=16'hcc67;
27366: douta=16'hd467;
27367: douta=16'hd468;
27368: douta=16'hd467;
27369: douta=16'hcc67;
27370: douta=16'hd468;
27371: douta=16'hd487;
27372: douta=16'hd487;
27373: douta=16'hd467;
27374: douta=16'hd487;
27375: douta=16'hd467;
27376: douta=16'hd487;
27377: douta=16'hd467;
27378: douta=16'hd468;
27379: douta=16'hd488;
27380: douta=16'hd488;
27381: douta=16'hd467;
27382: douta=16'hd488;
27383: douta=16'hcc68;
27384: douta=16'hd468;
27385: douta=16'hd487;
27386: douta=16'hb4ce;
27387: douta=16'hce76;
27388: douta=16'hd468;
27389: douta=16'hd488;
27390: douta=16'hcc87;
27391: douta=16'hcc69;
27392: douta=16'h942f;
27393: douta=16'h9c92;
27394: douta=16'h9c93;
27395: douta=16'h9473;
27396: douta=16'h9c93;
27397: douta=16'h8432;
27398: douta=16'h8c53;
27399: douta=16'h8c32;
27400: douta=16'h7bd2;
27401: douta=16'h736e;
27402: douta=16'h736f;
27403: douta=16'h6aeb;
27404: douta=16'h3984;
27405: douta=16'h3944;
27406: douta=16'h734c;
27407: douta=16'h734b;
27408: douta=16'h6b0a;
27409: douta=16'h732b;
27410: douta=16'h736b;
27411: douta=16'h7b8b;
27412: douta=16'h8bed;
27413: douta=16'hacb0;
27414: douta=16'ha490;
27415: douta=16'ha48f;
27416: douta=16'h9c4e;
27417: douta=16'ha46e;
27418: douta=16'haccf;
27419: douta=16'hbd31;
27420: douta=16'hc572;
27421: douta=16'hcdb4;
27422: douta=16'hd5d4;
27423: douta=16'hd5f4;
27424: douta=16'hde15;
27425: douta=16'hddf4;
27426: douta=16'hd5d4;
27427: douta=16'hc593;
27428: douta=16'hcd94;
27429: douta=16'hc573;
27430: douta=16'hbd33;
27431: douta=16'hbd53;
27432: douta=16'hb513;
27433: douta=16'h9472;
27434: douta=16'h8431;
27435: douta=16'h634e;
27436: douta=16'h4a6b;
27437: douta=16'h426b;
27438: douta=16'h3a4c;
27439: douta=16'h62ec;
27440: douta=16'h0883;
27441: douta=16'h18c5;
27442: douta=16'h2147;
27443: douta=16'h18e5;
27444: douta=16'h1946;
27445: douta=16'h59e6;
27446: douta=16'h51c6;
27447: douta=16'h51c5;
27448: douta=16'h51c6;
27449: douta=16'h51c6;
27450: douta=16'h51c6;
27451: douta=16'h51c5;
27452: douta=16'h51a6;
27453: douta=16'h51c6;
27454: douta=16'h51c6;
27455: douta=16'h59e6;
27456: douta=16'hbd12;
27457: douta=16'hcdd6;
27458: douta=16'hb535;
27459: douta=16'had14;
27460: douta=16'hd616;
27461: douta=16'hc595;
27462: douta=16'hb554;
27463: douta=16'h9494;
27464: douta=16'h9474;
27465: douta=16'h94b4;
27466: douta=16'h94b5;
27467: douta=16'h9495;
27468: douta=16'h8474;
27469: douta=16'h8c94;
27470: douta=16'h9d59;
27471: douta=16'h6b90;
27472: douta=16'h20c3;
27473: douta=16'h20a3;
27474: douta=16'h20c3;
27475: douta=16'h20c3;
27476: douta=16'h20c3;
27477: douta=16'h20e3;
27478: douta=16'h1881;
27479: douta=16'h20a2;
27480: douta=16'h18a2;
27481: douta=16'h20a2;
27482: douta=16'h20a2;
27483: douta=16'h20a2;
27484: douta=16'h2082;
27485: douta=16'h20c2;
27486: douta=16'h28e2;
27487: douta=16'h28c2;
27488: douta=16'h28e3;
27489: douta=16'h28e2;
27490: douta=16'h3103;
27491: douta=16'h3103;
27492: douta=16'h3986;
27493: douta=16'h10c5;
27494: douta=16'h4963;
27495: douta=16'h4963;
27496: douta=16'h5184;
27497: douta=16'h5184;
27498: douta=16'h59a4;
27499: douta=16'h59c4;
27500: douta=16'h61e4;
27501: douta=16'h59a3;
27502: douta=16'h940c;
27503: douta=16'h6a24;
27504: douta=16'h6a24;
27505: douta=16'h7a64;
27506: douta=16'h6204;
27507: douta=16'h7a64;
27508: douta=16'h7a84;
27509: douta=16'h7a84;
27510: douta=16'h7a84;
27511: douta=16'h7a64;
27512: douta=16'h8285;
27513: douta=16'h7a64;
27514: douta=16'h82a5;
27515: douta=16'h8ac4;
27516: douta=16'h8ac5;
27517: douta=16'h9305;
27518: douta=16'h9325;
27519: douta=16'h9b45;
27520: douta=16'ha345;
27521: douta=16'ha345;
27522: douta=16'hab65;
27523: douta=16'hb385;
27524: douta=16'hb3a6;
27525: douta=16'hb3a6;
27526: douta=16'hbbc6;
27527: douta=16'hbbc6;
27528: douta=16'hbbe6;
27529: douta=16'hbbe6;
27530: douta=16'hbbe5;
27531: douta=16'hbc06;
27532: douta=16'hc406;
27533: douta=16'hc405;
27534: douta=16'hc426;
27535: douta=16'hc426;
27536: douta=16'hc426;
27537: douta=16'hc426;
27538: douta=16'hc426;
27539: douta=16'hcc46;
27540: douta=16'hcc46;
27541: douta=16'hcc26;
27542: douta=16'hcc46;
27543: douta=16'hcc47;
27544: douta=16'hcc47;
27545: douta=16'hcc47;
27546: douta=16'hcc47;
27547: douta=16'hcc47;
27548: douta=16'hcc46;
27549: douta=16'hcc46;
27550: douta=16'hcc67;
27551: douta=16'hcc67;
27552: douta=16'hcc47;
27553: douta=16'hcc46;
27554: douta=16'hd467;
27555: douta=16'hd467;
27556: douta=16'hd468;
27557: douta=16'hd467;
27558: douta=16'hd467;
27559: douta=16'hcc67;
27560: douta=16'hd467;
27561: douta=16'hd467;
27562: douta=16'hcc67;
27563: douta=16'hd487;
27564: douta=16'hd467;
27565: douta=16'hd487;
27566: douta=16'hd467;
27567: douta=16'hd467;
27568: douta=16'hd467;
27569: douta=16'hd467;
27570: douta=16'hd487;
27571: douta=16'hd487;
27572: douta=16'hd487;
27573: douta=16'hd488;
27574: douta=16'hd488;
27575: douta=16'hd488;
27576: douta=16'hd487;
27577: douta=16'hd467;
27578: douta=16'haccd;
27579: douta=16'hd677;
27580: douta=16'hd467;
27581: douta=16'hcc68;
27582: douta=16'hd468;
27583: douta=16'hd485;
27584: douta=16'hc468;
27585: douta=16'h9430;
27586: douta=16'h8bf1;
27587: douta=16'h83f1;
27588: douta=16'h83d1;
27589: douta=16'h7bf1;
27590: douta=16'h738f;
27591: douta=16'h8c33;
27592: douta=16'h4a26;
27593: douta=16'h49e6;
27594: douta=16'h3964;
27595: douta=16'h4a06;
27596: douta=16'h5a68;
27597: douta=16'h62aa;
27598: douta=16'h8bcd;
27599: douta=16'h6b0a;
27600: douta=16'h838d;
27601: douta=16'h83ad;
27602: douta=16'h83cd;
27603: douta=16'h93ee;
27604: douta=16'h5268;
27605: douta=16'h942f;
27606: douta=16'hac8f;
27607: douta=16'hb4d0;
27608: douta=16'hb4f0;
27609: douta=16'hbd51;
27610: douta=16'hcd92;
27611: douta=16'hd5d3;
27612: douta=16'hcdb3;
27613: douta=16'hcdd3;
27614: douta=16'hd615;
27615: douta=16'hd614;
27616: douta=16'hd5f4;
27617: douta=16'hd5b3;
27618: douta=16'hcd73;
27619: douta=16'hb4f3;
27620: douta=16'hb4f3;
27621: douta=16'hacf3;
27622: douta=16'hacd3;
27623: douta=16'ha4b3;
27624: douta=16'ha4d3;
27625: douta=16'h9cd3;
27626: douta=16'h8c93;
27627: douta=16'h7c32;
27628: douta=16'h5b0e;
27629: douta=16'h422a;
27630: douta=16'h2987;
27631: douta=16'h52ac;
27632: douta=16'h1927;
27633: douta=16'h2127;
27634: douta=16'h2105;
27635: douta=16'h18c5;
27636: douta=16'h2168;
27637: douta=16'h51c5;
27638: douta=16'h59e6;
27639: douta=16'h51c6;
27640: douta=16'h51c5;
27641: douta=16'h59e6;
27642: douta=16'h51c6;
27643: douta=16'h59e6;
27644: douta=16'h59e6;
27645: douta=16'h59c6;
27646: douta=16'h59e6;
27647: douta=16'h59e6;
27648: douta=16'hcd54;
27649: douta=16'hc575;
27650: douta=16'hb534;
27651: douta=16'hacf4;
27652: douta=16'hcdb5;
27653: douta=16'hbd75;
27654: douta=16'hb555;
27655: douta=16'h8c73;
27656: douta=16'h9474;
27657: douta=16'h94b4;
27658: douta=16'h94d5;
27659: douta=16'h8c94;
27660: douta=16'h8454;
27661: douta=16'h8474;
27662: douta=16'h9517;
27663: douta=16'h31c6;
27664: douta=16'h20c2;
27665: douta=16'h20a3;
27666: douta=16'h20c3;
27667: douta=16'h20a3;
27668: douta=16'h20a3;
27669: douta=16'h20c3;
27670: douta=16'h20a2;
27671: douta=16'h20a2;
27672: douta=16'h20a2;
27673: douta=16'h20c2;
27674: douta=16'h20a2;
27675: douta=16'h20a2;
27676: douta=16'h20a2;
27677: douta=16'h20a2;
27678: douta=16'h28c2;
27679: douta=16'h28c2;
27680: douta=16'h28e2;
27681: douta=16'h30e3;
27682: douta=16'h3103;
27683: douta=16'h3903;
27684: douta=16'h41c8;
27685: douta=16'h10a4;
27686: douta=16'h4963;
27687: douta=16'h4964;
27688: douta=16'h5184;
27689: douta=16'h5184;
27690: douta=16'h59a4;
27691: douta=16'h59c4;
27692: douta=16'h61c3;
27693: douta=16'h61c4;
27694: douta=16'h8b8a;
27695: douta=16'h7244;
27696: douta=16'h6a04;
27697: douta=16'h7244;
27698: douta=16'h7224;
27699: douta=16'h6a04;
27700: douta=16'h7a64;
27701: douta=16'h7aa4;
27702: douta=16'h7a84;
27703: douta=16'h82a5;
27704: douta=16'h8285;
27705: douta=16'h82a4;
27706: douta=16'h82a4;
27707: douta=16'h8ac5;
27708: douta=16'h8ac4;
27709: douta=16'h9305;
27710: douta=16'h9325;
27711: douta=16'ha346;
27712: douta=16'ha345;
27713: douta=16'ha366;
27714: douta=16'hab85;
27715: douta=16'hb385;
27716: douta=16'hb3a6;
27717: douta=16'hb3a5;
27718: douta=16'hbbc6;
27719: douta=16'hbbc6;
27720: douta=16'hbbe6;
27721: douta=16'hbbe5;
27722: douta=16'hbbe5;
27723: douta=16'hbbe5;
27724: douta=16'hbc06;
27725: douta=16'hc426;
27726: douta=16'hc405;
27727: douta=16'hc426;
27728: douta=16'hc426;
27729: douta=16'hc426;
27730: douta=16'hc426;
27731: douta=16'hcc46;
27732: douta=16'hcc47;
27733: douta=16'hcc26;
27734: douta=16'hc446;
27735: douta=16'hcc47;
27736: douta=16'hcc46;
27737: douta=16'hcc46;
27738: douta=16'hcc47;
27739: douta=16'hcc67;
27740: douta=16'hcc47;
27741: douta=16'hcc67;
27742: douta=16'hcc67;
27743: douta=16'hcc67;
27744: douta=16'hd467;
27745: douta=16'hcc67;
27746: douta=16'hd467;
27747: douta=16'hd467;
27748: douta=16'hcc67;
27749: douta=16'hcc67;
27750: douta=16'hcc67;
27751: douta=16'hd467;
27752: douta=16'hd467;
27753: douta=16'hd467;
27754: douta=16'hd467;
27755: douta=16'hd467;
27756: douta=16'hd487;
27757: douta=16'hd487;
27758: douta=16'hd467;
27759: douta=16'hd467;
27760: douta=16'hd467;
27761: douta=16'hd467;
27762: douta=16'hd487;
27763: douta=16'hd488;
27764: douta=16'hd488;
27765: douta=16'hd488;
27766: douta=16'hd487;
27767: douta=16'hd487;
27768: douta=16'hd487;
27769: douta=16'hd468;
27770: douta=16'hb50e;
27771: douta=16'hceb7;
27772: douta=16'hcc68;
27773: douta=16'hcc88;
27774: douta=16'hd487;
27775: douta=16'hcc68;
27776: douta=16'hdca5;
27777: douta=16'h83d1;
27778: douta=16'h8bf1;
27779: douta=16'h736f;
27780: douta=16'h7b90;
27781: douta=16'h734e;
27782: douta=16'h734e;
27783: douta=16'h5a8a;
27784: douta=16'h3965;
27785: douta=16'h49c5;
27786: douta=16'h5206;
27787: douta=16'h6aea;
27788: douta=16'h62e9;
27789: douta=16'h7b6c;
27790: douta=16'h7b4c;
27791: douta=16'h732b;
27792: douta=16'h940e;
27793: douta=16'h940e;
27794: douta=16'h9c2e;
27795: douta=16'ha46f;
27796: douta=16'h5a69;
27797: douta=16'h838c;
27798: douta=16'ha490;
27799: douta=16'hbd11;
27800: douta=16'hc551;
27801: douta=16'hc572;
27802: douta=16'hd5d4;
27803: douta=16'hd5f4;
27804: douta=16'hde15;
27805: douta=16'hcd93;
27806: douta=16'hd5b3;
27807: douta=16'hd5b4;
27808: douta=16'hc553;
27809: douta=16'hb513;
27810: douta=16'hb4f3;
27811: douta=16'hacd3;
27812: douta=16'ha4d4;
27813: douta=16'ha4d4;
27814: douta=16'h94b5;
27815: douta=16'h9cb4;
27816: douta=16'h94b4;
27817: douta=16'h94d4;
27818: douta=16'h94b4;
27819: douta=16'h8453;
27820: douta=16'h7cb6;
27821: douta=16'h7434;
27822: douta=16'h4a8d;
27823: douta=16'h39e8;
27824: douta=16'h2988;
27825: douta=16'h2968;
27826: douta=16'h18c4;
27827: douta=16'h10a4;
27828: douta=16'h1946;
27829: douta=16'h59e6;
27830: douta=16'h51e6;
27831: douta=16'h59e6;
27832: douta=16'h59e6;
27833: douta=16'h59e6;
27834: douta=16'h51c6;
27835: douta=16'h59e6;
27836: douta=16'h59e6;
27837: douta=16'h6206;
27838: douta=16'h6206;
27839: douta=16'h6206;
27840: douta=16'hde16;
27841: douta=16'hb514;
27842: douta=16'hb555;
27843: douta=16'hb555;
27844: douta=16'hbd75;
27845: douta=16'hbd55;
27846: douta=16'had35;
27847: douta=16'h9473;
27848: douta=16'h9cb4;
27849: douta=16'h94b5;
27850: douta=16'h94b5;
27851: douta=16'h8c74;
27852: douta=16'h8433;
27853: douta=16'h9d58;
27854: douta=16'h0800;
27855: douta=16'h20c3;
27856: douta=16'h20c3;
27857: douta=16'h20a3;
27858: douta=16'h20c3;
27859: douta=16'h20c3;
27860: douta=16'h20c3;
27861: douta=16'h20a2;
27862: douta=16'h1881;
27863: douta=16'h1881;
27864: douta=16'h2082;
27865: douta=16'h20a2;
27866: douta=16'h20a2;
27867: douta=16'h20a2;
27868: douta=16'h20a2;
27869: douta=16'h20c2;
27870: douta=16'h20c2;
27871: douta=16'h28e2;
27872: douta=16'h30e3;
27873: douta=16'h3103;
27874: douta=16'h3923;
27875: douta=16'h3902;
27876: douta=16'h3a09;
27877: douta=16'h20a4;
27878: douta=16'h4984;
27879: douta=16'h4964;
27880: douta=16'h51a4;
27881: douta=16'h51a4;
27882: douta=16'h59a4;
27883: douta=16'h61c4;
27884: douta=16'h61c3;
27885: douta=16'h6267;
27886: douta=16'h6a04;
27887: douta=16'h7224;
27888: douta=16'h7224;
27889: douta=16'h7244;
27890: douta=16'h8285;
27891: douta=16'h4984;
27892: douta=16'h8284;
27893: douta=16'h7a64;
27894: douta=16'h8284;
27895: douta=16'h8285;
27896: douta=16'h8284;
27897: douta=16'h82a4;
27898: douta=16'h8ac5;
27899: douta=16'h8ac5;
27900: douta=16'h8ac4;
27901: douta=16'h9305;
27902: douta=16'h9b26;
27903: douta=16'ha346;
27904: douta=16'ha345;
27905: douta=16'hab85;
27906: douta=16'hab65;
27907: douta=16'hb3a5;
27908: douta=16'hb3a6;
27909: douta=16'hb3a5;
27910: douta=16'hbbc6;
27911: douta=16'hbbe6;
27912: douta=16'hbbe6;
27913: douta=16'hbc06;
27914: douta=16'hbc06;
27915: douta=16'hc406;
27916: douta=16'hc406;
27917: douta=16'hc406;
27918: douta=16'hc426;
27919: douta=16'hc426;
27920: douta=16'hc426;
27921: douta=16'hc426;
27922: douta=16'hc426;
27923: douta=16'hc426;
27924: douta=16'hc446;
27925: douta=16'hc446;
27926: douta=16'hcc47;
27927: douta=16'hcc47;
27928: douta=16'hcc67;
27929: douta=16'hcc47;
27930: douta=16'hcc47;
27931: douta=16'hcc47;
27932: douta=16'hcc47;
27933: douta=16'hcc67;
27934: douta=16'hcc67;
27935: douta=16'hcc67;
27936: douta=16'hcc47;
27937: douta=16'hcc67;
27938: douta=16'hcc67;
27939: douta=16'hcc67;
27940: douta=16'hcc67;
27941: douta=16'hd467;
27942: douta=16'hd467;
27943: douta=16'hd467;
27944: douta=16'hcc67;
27945: douta=16'hd488;
27946: douta=16'hd487;
27947: douta=16'hd487;
27948: douta=16'hd487;
27949: douta=16'hd487;
27950: douta=16'hd487;
27951: douta=16'hd487;
27952: douta=16'hcc67;
27953: douta=16'hd488;
27954: douta=16'hd488;
27955: douta=16'hd487;
27956: douta=16'hcc87;
27957: douta=16'hd488;
27958: douta=16'hd467;
27959: douta=16'hd466;
27960: douta=16'hcc66;
27961: douta=16'hd423;
27962: douta=16'ha48c;
27963: douta=16'hce76;
27964: douta=16'hcc69;
27965: douta=16'hccaa;
27966: douta=16'hd52d;
27967: douta=16'hd5f2;
27968: douta=16'he634;
27969: douta=16'hf6f8;
27970: douta=16'h83af;
27971: douta=16'h5a69;
27972: douta=16'h49e7;
27973: douta=16'h62ca;
27974: douta=16'h6b0b;
27975: douta=16'h6aea;
27976: douta=16'h6b0b;
27977: douta=16'h942f;
27978: douta=16'h9c4e;
27979: douta=16'h942f;
27980: douta=16'h942e;
27981: douta=16'hb510;
27982: douta=16'ha48f;
27983: douta=16'hcdd3;
27984: douta=16'hb511;
27985: douta=16'hbd31;
27986: douta=16'hc552;
27987: douta=16'hcdb3;
27988: douta=16'hbd52;
27989: douta=16'h62ca;
27990: douta=16'hacd1;
27991: douta=16'hcdb3;
27992: douta=16'hd5b3;
27993: douta=16'hcdb3;
27994: douta=16'hd5b3;
27995: douta=16'hcd53;
27996: douta=16'hb4f2;
27997: douta=16'h9cb3;
27998: douta=16'ha4d4;
27999: douta=16'h9cb4;
28000: douta=16'h94b4;
28001: douta=16'h8c93;
28002: douta=16'h8c73;
28003: douta=16'h8433;
28004: douta=16'h7bf1;
28005: douta=16'h7bf2;
28006: douta=16'h736e;
28007: douta=16'h5289;
28008: douta=16'h49e7;
28009: douta=16'h2081;
28010: douta=16'h20c2;
28011: douta=16'h4a06;
28012: douta=16'h5228;
28013: douta=16'h526a;
28014: douta=16'h5aee;
28015: douta=16'h29eb;
28016: douta=16'h62ee;
28017: douta=16'h0863;
28018: douta=16'h10a3;
28019: douta=16'h18e4;
28020: douta=16'h0001;
28021: douta=16'h59c5;
28022: douta=16'h59e6;
28023: douta=16'h59e7;
28024: douta=16'h59e6;
28025: douta=16'h6206;
28026: douta=16'h6206;
28027: douta=16'h6206;
28028: douta=16'h6226;
28029: douta=16'h6206;
28030: douta=16'h6206;
28031: douta=16'h6a26;
28032: douta=16'he678;
28033: douta=16'hbd34;
28034: douta=16'had15;
28035: douta=16'hcdb5;
28036: douta=16'hbd75;
28037: douta=16'hbd55;
28038: douta=16'ha4f5;
28039: douta=16'h9473;
28040: douta=16'ha4f5;
28041: douta=16'h94d5;
28042: douta=16'h8c75;
28043: douta=16'h8453;
28044: douta=16'h8454;
28045: douta=16'h52cc;
28046: douta=16'h20c3;
28047: douta=16'h20c3;
28048: douta=16'h20e3;
28049: douta=16'h20c3;
28050: douta=16'h20c3;
28051: douta=16'h20a3;
28052: douta=16'h20c3;
28053: douta=16'h1881;
28054: douta=16'h2082;
28055: douta=16'h20a2;
28056: douta=16'h1881;
28057: douta=16'h20a2;
28058: douta=16'h20a2;
28059: douta=16'h20a2;
28060: douta=16'h20c2;
28061: douta=16'h28c2;
28062: douta=16'h28e3;
28063: douta=16'h28e2;
28064: douta=16'h30e2;
28065: douta=16'h30e2;
28066: douta=16'h3123;
28067: douta=16'h3903;
28068: douta=16'h3209;
28069: douta=16'h3104;
28070: douta=16'h4964;
28071: douta=16'h4964;
28072: douta=16'h59a4;
28073: douta=16'h59a4;
28074: douta=16'h59c4;
28075: douta=16'h61e4;
28076: douta=16'h61c3;
28077: douta=16'h6b0a;
28078: douta=16'h69e3;
28079: douta=16'h7224;
28080: douta=16'h7244;
28081: douta=16'h7244;
28082: douta=16'h7a44;
28083: douta=16'h4164;
28084: douta=16'h7a85;
28085: douta=16'h7aa5;
28086: douta=16'h7a64;
28087: douta=16'h8285;
28088: douta=16'h8285;
28089: douta=16'h82a4;
28090: douta=16'h8ac5;
28091: douta=16'h8ac5;
28092: douta=16'h8ac5;
28093: douta=16'h9305;
28094: douta=16'h9b25;
28095: douta=16'ha346;
28096: douta=16'ha366;
28097: douta=16'hab66;
28098: douta=16'hab85;
28099: douta=16'hb3a5;
28100: douta=16'hb3c6;
28101: douta=16'hb3c6;
28102: douta=16'hbbc6;
28103: douta=16'hbbe6;
28104: douta=16'hbbe6;
28105: douta=16'hbbe5;
28106: douta=16'hc405;
28107: douta=16'hbbe5;
28108: douta=16'hc406;
28109: douta=16'hc406;
28110: douta=16'hc406;
28111: douta=16'hc426;
28112: douta=16'hc426;
28113: douta=16'hc426;
28114: douta=16'hc426;
28115: douta=16'hcc26;
28116: douta=16'hc426;
28117: douta=16'hcc27;
28118: douta=16'hcc47;
28119: douta=16'hcc67;
28120: douta=16'hcc67;
28121: douta=16'hcc47;
28122: douta=16'hcc67;
28123: douta=16'hcc48;
28124: douta=16'hcc68;
28125: douta=16'hcc67;
28126: douta=16'hcc67;
28127: douta=16'hcc67;
28128: douta=16'hd467;
28129: douta=16'hcc87;
28130: douta=16'hcc87;
28131: douta=16'hd488;
28132: douta=16'hd467;
28133: douta=16'hd468;
28134: douta=16'hd468;
28135: douta=16'hcc67;
28136: douta=16'hcc67;
28137: douta=16'hcc68;
28138: douta=16'hd468;
28139: douta=16'hd487;
28140: douta=16'hd467;
28141: douta=16'hd466;
28142: douta=16'hcc45;
28143: douta=16'hcc25;
28144: douta=16'hcc23;
28145: douta=16'hcc25;
28146: douta=16'hcc47;
28147: douta=16'hcccb;
28148: douta=16'hd52e;
28149: douta=16'hd5b1;
28150: douta=16'he675;
28151: douta=16'he6b6;
28152: douta=16'hef19;
28153: douta=16'hf7bc;
28154: douta=16'hf79b;
28155: douta=16'hf77a;
28156: douta=16'hff9b;
28157: douta=16'hf799;
28158: douta=16'hef17;
28159: douta=16'he652;
28160: douta=16'he612;
28161: douta=16'hd5ae;
28162: douta=16'h93ce;
28163: douta=16'h7b6c;
28164: douta=16'h83cd;
28165: douta=16'h734b;
28166: douta=16'h7b6c;
28167: douta=16'h734c;
28168: douta=16'h8bee;
28169: douta=16'h944f;
28170: douta=16'h940e;
28171: douta=16'hb4d0;
28172: douta=16'hacaf;
28173: douta=16'hb4f0;
28174: douta=16'hde55;
28175: douta=16'hde35;
28176: douta=16'hbd12;
28177: douta=16'hd614;
28178: douta=16'hd5f4;
28179: douta=16'hcdb4;
28180: douta=16'hd5f4;
28181: douta=16'hc5d4;
28182: douta=16'hacd1;
28183: douta=16'hd5d4;
28184: douta=16'hd5b4;
28185: douta=16'hc554;
28186: douta=16'h9c92;
28187: douta=16'h9453;
28188: douta=16'h8452;
28189: douta=16'h8452;
28190: douta=16'h7bf1;
28191: douta=16'h8c53;
28192: douta=16'h7bd2;
28193: douta=16'h7bd1;
28194: douta=16'h7390;
28195: douta=16'h4a07;
28196: douta=16'h49e7;
28197: douta=16'h2903;
28198: douta=16'h1881;
28199: douta=16'h3144;
28200: douta=16'h3965;
28201: douta=16'h62ca;
28202: douta=16'h6aea;
28203: douta=16'h7b8d;
28204: douta=16'h52cd;
28205: douta=16'h52cd;
28206: douta=16'h52cd;
28207: douta=16'h5310;
28208: douta=16'h6b4f;
28209: douta=16'h4aef;
28210: douta=16'h2968;
28211: douta=16'h2127;
28212: douta=16'h08a4;
28213: douta=16'h7267;
28214: douta=16'h6206;
28215: douta=16'h6206;
28216: douta=16'h6a26;
28217: douta=16'h61e6;
28218: douta=16'h61c5;
28219: douta=16'h59a5;
28220: douta=16'h59a5;
28221: douta=16'h61e5;
28222: douta=16'h6a89;
28223: douta=16'h7b4b;
28224: douta=16'he698;
28225: douta=16'hc575;
28226: douta=16'ha4b4;
28227: douta=16'hd5f6;
28228: douta=16'hbd54;
28229: douta=16'hb555;
28230: douta=16'h9cb4;
28231: douta=16'h9473;
28232: douta=16'h9cd5;
28233: douta=16'h94b5;
28234: douta=16'h8c74;
28235: douta=16'h8c54;
28236: douta=16'h8c54;
28237: douta=16'h18a3;
28238: douta=16'h20c3;
28239: douta=16'h20e3;
28240: douta=16'h20e3;
28241: douta=16'h20c3;
28242: douta=16'h20c3;
28243: douta=16'h20a3;
28244: douta=16'h20c3;
28245: douta=16'h1881;
28246: douta=16'h20a2;
28247: douta=16'h20a2;
28248: douta=16'h20a2;
28249: douta=16'h20a2;
28250: douta=16'h20a2;
28251: douta=16'h20a2;
28252: douta=16'h20a2;
28253: douta=16'h28e2;
28254: douta=16'h28e2;
28255: douta=16'h28e2;
28256: douta=16'h30e2;
28257: douta=16'h3103;
28258: douta=16'h3923;
28259: douta=16'h3923;
28260: douta=16'h3a09;
28261: douta=16'h3923;
28262: douta=16'h4984;
28263: douta=16'h4984;
28264: douta=16'h51a4;
28265: douta=16'h51a4;
28266: douta=16'h59c4;
28267: douta=16'h61e4;
28268: douta=16'h61e3;
28269: douta=16'h7b6c;
28270: douta=16'h69c3;
28271: douta=16'h7224;
28272: douta=16'h7244;
28273: douta=16'h7244;
28274: douta=16'h7a65;
28275: douta=16'h4984;
28276: douta=16'h7aa4;
28277: douta=16'h8284;
28278: douta=16'h7a64;
28279: douta=16'h8285;
28280: douta=16'h8285;
28281: douta=16'h82a4;
28282: douta=16'h8ac4;
28283: douta=16'h8ac5;
28284: douta=16'h8ac4;
28285: douta=16'h9305;
28286: douta=16'h9b26;
28287: douta=16'ha346;
28288: douta=16'ha366;
28289: douta=16'hab86;
28290: douta=16'hb385;
28291: douta=16'hb385;
28292: douta=16'hb3c6;
28293: douta=16'hb3c6;
28294: douta=16'hbbc6;
28295: douta=16'hbbe6;
28296: douta=16'hbbe6;
28297: douta=16'hc406;
28298: douta=16'hbc06;
28299: douta=16'hc406;
28300: douta=16'hc406;
28301: douta=16'hc406;
28302: douta=16'hc406;
28303: douta=16'hc426;
28304: douta=16'hc426;
28305: douta=16'hc446;
28306: douta=16'hc426;
28307: douta=16'hc426;
28308: douta=16'hc426;
28309: douta=16'hcc47;
28310: douta=16'hcc47;
28311: douta=16'hcc26;
28312: douta=16'hcc47;
28313: douta=16'hcc67;
28314: douta=16'hcc47;
28315: douta=16'hcc67;
28316: douta=16'hcc67;
28317: douta=16'hcc66;
28318: douta=16'hcc67;
28319: douta=16'hcc67;
28320: douta=16'hcc67;
28321: douta=16'hd467;
28322: douta=16'hcc68;
28323: douta=16'hd468;
28324: douta=16'hd467;
28325: douta=16'hcc87;
28326: douta=16'hcc87;
28327: douta=16'hd467;
28328: douta=16'hd466;
28329: douta=16'hd446;
28330: douta=16'hcc21;
28331: douta=16'hcc23;
28332: douta=16'hcc03;
28333: douta=16'hcc67;
28334: douta=16'hcc89;
28335: douta=16'hd52c;
28336: douta=16'hddd1;
28337: douta=16'he655;
28338: douta=16'he697;
28339: douta=16'hef59;
28340: douta=16'hf79c;
28341: douta=16'hffdd;
28342: douta=16'hfffd;
28343: douta=16'hffdc;
28344: douta=16'hff9b;
28345: douta=16'hf6f7;
28346: douta=16'he694;
28347: douta=16'he632;
28348: douta=16'hd56d;
28349: douta=16'hd52b;
28350: douta=16'hcc88;
28351: douta=16'hcc46;
28352: douta=16'hcc26;
28353: douta=16'hc404;
28354: douta=16'hc48c;
28355: douta=16'h83ad;
28356: douta=16'h8c0e;
28357: douta=16'h83cd;
28358: douta=16'h7b8c;
28359: douta=16'h83ce;
28360: douta=16'h944f;
28361: douta=16'h9c4e;
28362: douta=16'ha4af;
28363: douta=16'hb4f0;
28364: douta=16'hb510;
28365: douta=16'hb4f0;
28366: douta=16'hd616;
28367: douta=16'hcdb4;
28368: douta=16'hacd2;
28369: douta=16'hcdb4;
28370: douta=16'hde34;
28371: douta=16'hcdd4;
28372: douta=16'hacd2;
28373: douta=16'hd5f6;
28374: douta=16'hbd33;
28375: douta=16'hd5b3;
28376: douta=16'hb514;
28377: douta=16'ha4d4;
28378: douta=16'h8c53;
28379: douta=16'h8432;
28380: douta=16'h83f2;
28381: douta=16'h7bb1;
28382: douta=16'h73d1;
28383: douta=16'h7c12;
28384: douta=16'h738e;
28385: douta=16'h62cb;
28386: douta=16'h5248;
28387: douta=16'h1881;
28388: douta=16'h1081;
28389: douta=16'h2924;
28390: douta=16'h3985;
28391: douta=16'h5227;
28392: douta=16'h5248;
28393: douta=16'h734b;
28394: douta=16'h734b;
28395: douta=16'h4a07;
28396: douta=16'h2925;
28397: douta=16'h2104;
28398: douta=16'h2104;
28399: douta=16'h4ace;
28400: douta=16'h632f;
28401: douta=16'h4acf;
28402: douta=16'h2989;
28403: douta=16'h29aa;
28404: douta=16'h10a4;
28405: douta=16'h728a;
28406: douta=16'h7247;
28407: douta=16'h59a5;
28408: douta=16'h59e6;
28409: douta=16'h6a47;
28410: douta=16'h72ca;
28411: douta=16'h838d;
28412: douta=16'h8c0e;
28413: douta=16'h9cb0;
28414: douta=16'hb554;
28415: douta=16'hbdd5;
28416: douta=16'hc595;
28417: douta=16'hb535;
28418: douta=16'hbd75;
28419: douta=16'hcdb6;
28420: douta=16'hbd75;
28421: douta=16'ha4f5;
28422: douta=16'h8c52;
28423: douta=16'ha4d4;
28424: douta=16'h94b4;
28425: douta=16'h94d5;
28426: douta=16'h8474;
28427: douta=16'h8c95;
28428: douta=16'h94f7;
28429: douta=16'h20e3;
28430: douta=16'h20c3;
28431: douta=16'h20c3;
28432: douta=16'h20c3;
28433: douta=16'h20e3;
28434: douta=16'h20c3;
28435: douta=16'h20c3;
28436: douta=16'h20e3;
28437: douta=16'h1882;
28438: douta=16'h2082;
28439: douta=16'h1881;
28440: douta=16'h20a2;
28441: douta=16'h20a2;
28442: douta=16'h20a2;
28443: douta=16'h20c2;
28444: douta=16'h28e3;
28445: douta=16'h28c2;
28446: douta=16'h28e2;
28447: douta=16'h30e2;
28448: douta=16'h3103;
28449: douta=16'h3103;
28450: douta=16'h3903;
28451: douta=16'h41a6;
28452: douta=16'h31c9;
28453: douta=16'h4963;
28454: douta=16'h4984;
28455: douta=16'h5184;
28456: douta=16'h51a4;
28457: douta=16'h59a4;
28458: douta=16'h59c4;
28459: douta=16'h61e4;
28460: douta=16'h6a67;
28461: douta=16'h94b1;
28462: douta=16'h69e4;
28463: douta=16'h7a65;
28464: douta=16'h7244;
28465: douta=16'h7a64;
28466: douta=16'h7a64;
28467: douta=16'h8285;
28468: douta=16'h8ac5;
28469: douta=16'h8285;
28470: douta=16'h8284;
28471: douta=16'h82a4;
28472: douta=16'h8aa5;
28473: douta=16'h82a5;
28474: douta=16'h8aa4;
28475: douta=16'h8ac4;
28476: douta=16'h8ac5;
28477: douta=16'h9305;
28478: douta=16'h9b26;
28479: douta=16'ha346;
28480: douta=16'ha366;
28481: douta=16'hab66;
28482: douta=16'hb385;
28483: douta=16'hb3a6;
28484: douta=16'hb3c6;
28485: douta=16'hb3c6;
28486: douta=16'hbbc6;
28487: douta=16'hbbe6;
28488: douta=16'hbbe5;
28489: douta=16'hc406;
28490: douta=16'hc406;
28491: douta=16'hc406;
28492: douta=16'hc406;
28493: douta=16'hc406;
28494: douta=16'hc406;
28495: douta=16'hc426;
28496: douta=16'hc427;
28497: douta=16'hc427;
28498: douta=16'hc426;
28499: douta=16'hc446;
28500: douta=16'hc426;
28501: douta=16'hcc47;
28502: douta=16'hc447;
28503: douta=16'hcc47;
28504: douta=16'hcc47;
28505: douta=16'hcc47;
28506: douta=16'hcc47;
28507: douta=16'hcc25;
28508: douta=16'hcc25;
28509: douta=16'hcc04;
28510: douta=16'hcc24;
28511: douta=16'hcc25;
28512: douta=16'hcc69;
28513: douta=16'hd52d;
28514: douta=16'hd590;
28515: douta=16'hddd1;
28516: douta=16'he696;
28517: douta=16'hef39;
28518: douta=16'hf79c;
28519: douta=16'hfffd;
28520: douta=16'hfffd;
28521: douta=16'hffbc;
28522: douta=16'hf758;
28523: douta=16'hf6f7;
28524: douta=16'heed5;
28525: douta=16'he5d0;
28526: douta=16'hddae;
28527: douta=16'hdd4c;
28528: douta=16'hd4c9;
28529: douta=16'hd487;
28530: douta=16'hcc87;
28531: douta=16'hcc46;
28532: douta=16'hcc47;
28533: douta=16'hd488;
28534: douta=16'hd488;
28535: douta=16'hd488;
28536: douta=16'hd488;
28537: douta=16'hcc88;
28538: douta=16'hd488;
28539: douta=16'hd488;
28540: douta=16'hcc68;
28541: douta=16'hcc68;
28542: douta=16'hd467;
28543: douta=16'hd468;
28544: douta=16'hcc67;
28545: douta=16'hcc68;
28546: douta=16'hc46a;
28547: douta=16'h9c2f;
28548: douta=16'h8bed;
28549: douta=16'ha4d0;
28550: douta=16'ha490;
28551: douta=16'ha4b0;
28552: douta=16'hb511;
28553: douta=16'hbd32;
28554: douta=16'hc572;
28555: douta=16'hcdb4;
28556: douta=16'hcdd4;
28557: douta=16'hd5f4;
28558: douta=16'heed7;
28559: douta=16'hcd94;
28560: douta=16'hbd54;
28561: douta=16'hacf4;
28562: douta=16'h7bf2;
28563: douta=16'h6bb2;
28564: douta=16'hc574;
28565: douta=16'ha4b5;
28566: douta=16'ha4d3;
28567: douta=16'h8c74;
28568: douta=16'h8453;
28569: douta=16'h8433;
28570: douta=16'h6bd1;
28571: douta=16'h6b0d;
28572: douta=16'h4a08;
28573: douta=16'h2902;
28574: douta=16'h20e1;
28575: douta=16'h28e3;
28576: douta=16'h3985;
28577: douta=16'h3985;
28578: douta=16'h39a5;
28579: douta=16'h5247;
28580: douta=16'h6ac9;
28581: douta=16'h6aea;
28582: douta=16'h736c;
28583: douta=16'h7b8d;
28584: douta=16'h83cd;
28585: douta=16'h8bed;
28586: douta=16'h9c4e;
28587: douta=16'h9c2f;
28588: douta=16'h2967;
28589: douta=16'h2146;
28590: douta=16'h10c4;
28591: douta=16'h10e5;
28592: douta=16'h2967;
28593: douta=16'h1906;
28594: douta=16'h29a9;
28595: douta=16'h2147;
28596: douta=16'h2967;
28597: douta=16'h10e6;
28598: douta=16'h08a5;
28599: douta=16'h39a6;
28600: douta=16'h6266;
28601: douta=16'h6246;
28602: douta=16'h6226;
28603: douta=16'h6a26;
28604: douta=16'h6a46;
28605: douta=16'h7266;
28606: douta=16'h7267;
28607: douta=16'h7287;
28608: douta=16'hb514;
28609: douta=16'ha4f5;
28610: douta=16'hcdb6;
28611: douta=16'hc595;
28612: douta=16'had35;
28613: douta=16'h94b4;
28614: douta=16'h9c94;
28615: douta=16'ha4f5;
28616: douta=16'h94d5;
28617: douta=16'h9cd6;
28618: douta=16'h8c74;
28619: douta=16'h9d17;
28620: douta=16'h18a2;
28621: douta=16'h28e3;
28622: douta=16'h20e3;
28623: douta=16'h20e3;
28624: douta=16'h20c3;
28625: douta=16'h20e3;
28626: douta=16'h20c3;
28627: douta=16'h20e3;
28628: douta=16'h20c3;
28629: douta=16'h2082;
28630: douta=16'h2082;
28631: douta=16'h20a2;
28632: douta=16'h20a2;
28633: douta=16'h2082;
28634: douta=16'h20a2;
28635: douta=16'h20c2;
28636: douta=16'h20c2;
28637: douta=16'h28e2;
28638: douta=16'h28e2;
28639: douta=16'h3103;
28640: douta=16'h30e3;
28641: douta=16'h3103;
28642: douta=16'h3923;
28643: douta=16'h4209;
28644: douta=16'h2988;
28645: douta=16'h5164;
28646: douta=16'h51a4;
28647: douta=16'h51a4;
28648: douta=16'h59c4;
28649: douta=16'h59a4;
28650: douta=16'h61e4;
28651: douta=16'h61e4;
28652: douta=16'h6ac9;
28653: douta=16'had53;
28654: douta=16'h7245;
28655: douta=16'h7244;
28656: douta=16'h7244;
28657: douta=16'h7a44;
28658: douta=16'h7a64;
28659: douta=16'h8284;
28660: douta=16'h7244;
28661: douta=16'h8285;
28662: douta=16'h8285;
28663: douta=16'h82a4;
28664: douta=16'h8ac5;
28665: douta=16'h8ac5;
28666: douta=16'h8ac5;
28667: douta=16'h8ac5;
28668: douta=16'h8ac5;
28669: douta=16'h9b26;
28670: douta=16'ha326;
28671: douta=16'ha346;
28672: douta=16'hab86;
28673: douta=16'haba6;
28674: douta=16'hb385;
28675: douta=16'hb3a5;
28676: douta=16'hb3c6;
28677: douta=16'hbbc6;
28678: douta=16'hbbc6;
28679: douta=16'hbbe6;
28680: douta=16'hbbe6;
28681: douta=16'hc406;
28682: douta=16'hbc05;
28683: douta=16'hc406;
28684: douta=16'hc406;
28685: douta=16'hc426;
28686: douta=16'hc426;
28687: douta=16'hc426;
28688: douta=16'hc425;
28689: douta=16'hc405;
28690: douta=16'hc404;
28691: douta=16'hc3e3;
28692: douta=16'hc3e3;
28693: douta=16'hc405;
28694: douta=16'hc447;
28695: douta=16'hcc6a;
28696: douta=16'hd54e;
28697: douta=16'hddb0;
28698: douta=16'hde34;
28699: douta=16'heef8;
28700: douta=16'hf77b;
28701: douta=16'hf7bb;
28702: douta=16'hfffd;
28703: douta=16'hffdc;
28704: douta=16'hff9a;
28705: douta=16'hef16;
28706: douta=16'he694;
28707: douta=16'he653;
28708: douta=16'hddae;
28709: douta=16'hd52b;
28710: douta=16'hd4ca;
28711: douta=16'hcc87;
28712: douta=16'hcc45;
28713: douta=16'hcc46;
28714: douta=16'hcc46;
28715: douta=16'hcc47;
28716: douta=16'hcc67;
28717: douta=16'hd467;
28718: douta=16'hd467;
28719: douta=16'hd488;
28720: douta=16'hd487;
28721: douta=16'hd488;
28722: douta=16'hcc88;
28723: douta=16'hd488;
28724: douta=16'hd488;
28725: douta=16'hd488;
28726: douta=16'hcc88;
28727: douta=16'hcc88;
28728: douta=16'hd488;
28729: douta=16'hd488;
28730: douta=16'hcc88;
28731: douta=16'hd488;
28732: douta=16'hcc68;
28733: douta=16'hcc88;
28734: douta=16'hcc67;
28735: douta=16'hcc68;
28736: douta=16'hcc68;
28737: douta=16'hcc68;
28738: douta=16'hcc68;
28739: douta=16'h9c70;
28740: douta=16'h9c50;
28741: douta=16'h9c70;
28742: douta=16'ha4b0;
28743: douta=16'hb511;
28744: douta=16'hbd72;
28745: douta=16'hcd94;
28746: douta=16'hcdb4;
28747: douta=16'hd5f5;
28748: douta=16'hd5f5;
28749: douta=16'hcd93;
28750: douta=16'hb4f3;
28751: douta=16'hacf4;
28752: douta=16'hc555;
28753: douta=16'h94b4;
28754: douta=16'h8c74;
28755: douta=16'h73d1;
28756: douta=16'h6bb2;
28757: douta=16'h8433;
28758: douta=16'h73d2;
28759: douta=16'h6b91;
28760: douta=16'h4a6a;
28761: douta=16'h39c7;
28762: douta=16'h1881;
28763: douta=16'h2923;
28764: douta=16'h3965;
28765: douta=16'h41c5;
28766: douta=16'h5227;
28767: douta=16'h5207;
28768: douta=16'h6b0a;
28769: douta=16'h6ac9;
28770: douta=16'h6ae9;
28771: douta=16'h734b;
28772: douta=16'h7b4b;
28773: douta=16'h7b4b;
28774: douta=16'h9c4f;
28775: douta=16'ha46f;
28776: douta=16'hacaf;
28777: douta=16'hb4d0;
28778: douta=16'ha46f;
28779: douta=16'h9c6f;
28780: douta=16'h62ed;
28781: douta=16'h3a2b;
28782: douta=16'h2967;
28783: douta=16'h10c3;
28784: douta=16'h0882;
28785: douta=16'h08c3;
28786: douta=16'h10a4;
28787: douta=16'h10e5;
28788: douta=16'h2147;
28789: douta=16'h1906;
28790: douta=16'h1948;
28791: douta=16'h1905;
28792: douta=16'h7267;
28793: douta=16'h7286;
28794: douta=16'h7a67;
28795: douta=16'h7a87;
28796: douta=16'h7a87;
28797: douta=16'h7a87;
28798: douta=16'h7a86;
28799: douta=16'h7a87;
28800: douta=16'hb513;
28801: douta=16'ha4f5;
28802: douta=16'hcdf6;
28803: douta=16'hbd75;
28804: douta=16'ha4f4;
28805: douta=16'h8c73;
28806: douta=16'ha4d5;
28807: douta=16'ha4d5;
28808: douta=16'h94d5;
28809: douta=16'h9cd6;
28810: douta=16'h8474;
28811: douta=16'ha559;
28812: douta=16'h1040;
28813: douta=16'h20c3;
28814: douta=16'h20e3;
28815: douta=16'h20c3;
28816: douta=16'h20e3;
28817: douta=16'h20c3;
28818: douta=16'h20a3;
28819: douta=16'h20e3;
28820: douta=16'h20e3;
28821: douta=16'h2082;
28822: douta=16'h20a2;
28823: douta=16'h2082;
28824: douta=16'h20a2;
28825: douta=16'h20a2;
28826: douta=16'h20a2;
28827: douta=16'h20c2;
28828: douta=16'h28e2;
28829: douta=16'h28e2;
28830: douta=16'h28e2;
28831: douta=16'h30e3;
28832: douta=16'h30e3;
28833: douta=16'h3103;
28834: douta=16'h3924;
28835: douta=16'h422a;
28836: douta=16'h1926;
28837: douta=16'h5184;
28838: douta=16'h5184;
28839: douta=16'h5184;
28840: douta=16'h59c4;
28841: douta=16'h59c4;
28842: douta=16'h61c3;
28843: douta=16'h6a04;
28844: douta=16'h732b;
28845: douta=16'hb595;
28846: douta=16'h7224;
28847: douta=16'h7244;
28848: douta=16'h7a44;
28849: douta=16'h7a65;
28850: douta=16'h7a84;
28851: douta=16'h7a64;
28852: douta=16'h6a44;
28853: douta=16'h8284;
28854: douta=16'h8285;
28855: douta=16'h8aa4;
28856: douta=16'h8ac5;
28857: douta=16'h8aa4;
28858: douta=16'h92e5;
28859: douta=16'h8ac5;
28860: douta=16'h8ac5;
28861: douta=16'h9305;
28862: douta=16'h9b26;
28863: douta=16'ha346;
28864: douta=16'hab86;
28865: douta=16'hab66;
28866: douta=16'hb3a5;
28867: douta=16'hb3a6;
28868: douta=16'hb3c6;
28869: douta=16'hbbc6;
28870: douta=16'hbbe6;
28871: douta=16'hbbe6;
28872: douta=16'hbbe6;
28873: douta=16'hbc05;
28874: douta=16'hbbe5;
28875: douta=16'hc3e7;
28876: douta=16'hc3e5;
28877: douta=16'hc3c4;
28878: douta=16'hbbc3;
28879: douta=16'hc3c3;
28880: douta=16'hc3e4;
28881: douta=16'hc427;
28882: douta=16'hccaa;
28883: douta=16'hd52e;
28884: douta=16'hd56f;
28885: douta=16'hde13;
28886: douta=16'he696;
28887: douta=16'hef19;
28888: douta=16'hf7bc;
28889: douta=16'hf7bd;
28890: douta=16'hffdc;
28891: douta=16'hf77a;
28892: douta=16'hef17;
28893: douta=16'heef6;
28894: douta=16'hddf0;
28895: douta=16'hddcf;
28896: douta=16'hd54c;
28897: douta=16'hcca9;
28898: douta=16'hd487;
28899: douta=16'hcc67;
28900: douta=16'hcc25;
28901: douta=16'hcc46;
28902: douta=16'hcc46;
28903: douta=16'hd467;
28904: douta=16'hcc68;
28905: douta=16'hcc88;
28906: douta=16'hcc87;
28907: douta=16'hcc87;
28908: douta=16'hd487;
28909: douta=16'hd487;
28910: douta=16'hd487;
28911: douta=16'hd488;
28912: douta=16'hd488;
28913: douta=16'hcc88;
28914: douta=16'hcc88;
28915: douta=16'hcc88;
28916: douta=16'hd488;
28917: douta=16'hd488;
28918: douta=16'hcc88;
28919: douta=16'hd488;
28920: douta=16'hcc88;
28921: douta=16'hd488;
28922: douta=16'hcc88;
28923: douta=16'hcc68;
28924: douta=16'hcc68;
28925: douta=16'hd488;
28926: douta=16'hcc67;
28927: douta=16'hd468;
28928: douta=16'hcc69;
28929: douta=16'hcc67;
28930: douta=16'hd466;
28931: douta=16'h9c91;
28932: douta=16'h9c2f;
28933: douta=16'ha490;
28934: douta=16'ha4b0;
28935: douta=16'hbd32;
28936: douta=16'hc573;
28937: douta=16'hcdd4;
28938: douta=16'hcdb4;
28939: douta=16'hd5f4;
28940: douta=16'hcdb4;
28941: douta=16'hc553;
28942: douta=16'h9473;
28943: douta=16'h7c13;
28944: douta=16'ha4d4;
28945: douta=16'had16;
28946: douta=16'h7bf3;
28947: douta=16'h73d2;
28948: douta=16'h73d2;
28949: douta=16'h6b4f;
28950: douta=16'h6b4f;
28951: douta=16'h3186;
28952: douta=16'h2903;
28953: douta=16'h28e3;
28954: douta=16'h39a5;
28955: douta=16'h62a9;
28956: douta=16'h5a68;
28957: douta=16'h5227;
28958: douta=16'h5a47;
28959: douta=16'h4a06;
28960: douta=16'h83ac;
28961: douta=16'h836c;
28962: douta=16'h7b2b;
28963: douta=16'h8bcb;
28964: douta=16'h93ec;
28965: douta=16'ha44e;
28966: douta=16'ha46f;
28967: douta=16'haccf;
28968: douta=16'hb510;
28969: douta=16'hbd30;
28970: douta=16'hac8f;
28971: douta=16'h9c2f;
28972: douta=16'h6b4d;
28973: douta=16'h52ac;
28974: douta=16'h3209;
28975: douta=16'h2126;
28976: douta=16'h10a3;
28977: douta=16'h1083;
28978: douta=16'h10c3;
28979: douta=16'h10e4;
28980: douta=16'h1927;
28981: douta=16'h08a4;
28982: douta=16'h2188;
28983: douta=16'h08e6;
28984: douta=16'h7267;
28985: douta=16'h7a87;
28986: douta=16'h8287;
28987: douta=16'h7a87;
28988: douta=16'h7a87;
28989: douta=16'h82a7;
28990: douta=16'h7a87;
28991: douta=16'h7aa7;
28992: douta=16'hbd75;
28993: douta=16'hbd75;
28994: douta=16'hcdd6;
28995: douta=16'hc575;
28996: douta=16'h8c32;
28997: douta=16'h8c73;
28998: douta=16'h94b5;
28999: douta=16'h9cd5;
29000: douta=16'h9cf6;
29001: douta=16'h94d5;
29002: douta=16'ha579;
29003: douta=16'h5b0c;
29004: douta=16'h28e3;
29005: douta=16'h20c3;
29006: douta=16'h28e3;
29007: douta=16'h20a3;
29008: douta=16'h20c3;
29009: douta=16'h20e3;
29010: douta=16'h20c3;
29011: douta=16'h20e3;
29012: douta=16'h1882;
29013: douta=16'h20a2;
29014: douta=16'h1881;
29015: douta=16'h20a2;
29016: douta=16'h20a2;
29017: douta=16'h20a2;
29018: douta=16'h20c2;
29019: douta=16'h20c2;
29020: douta=16'h28c2;
29021: douta=16'h28c2;
29022: douta=16'h28e2;
29023: douta=16'h3103;
29024: douta=16'h3103;
29025: douta=16'h3103;
29026: douta=16'h41c7;
29027: douta=16'h424b;
29028: douta=16'h18e6;
29029: douta=16'h5184;
29030: douta=16'h5184;
29031: douta=16'h51a4;
29032: douta=16'h59c4;
29033: douta=16'h59c4;
29034: douta=16'h61e4;
29035: douta=16'h61c3;
29036: douta=16'h9491;
29037: douta=16'hb572;
29038: douta=16'h7245;
29039: douta=16'h7244;
29040: douta=16'h7a64;
29041: douta=16'h7a64;
29042: douta=16'h7a84;
29043: douta=16'h8285;
29044: douta=16'h51c4;
29045: douta=16'h82a4;
29046: douta=16'h7aa5;
29047: douta=16'h8aa5;
29048: douta=16'h8ac5;
29049: douta=16'h8ac5;
29050: douta=16'h8ae5;
29051: douta=16'h92e5;
29052: douta=16'h8ac5;
29053: douta=16'h92c4;
29054: douta=16'h9ae4;
29055: douta=16'h9ae4;
29056: douta=16'ha304;
29057: douta=16'ha344;
29058: douta=16'hab85;
29059: douta=16'hb408;
29060: douta=16'hc4ac;
29061: douta=16'hc4ee;
29062: douta=16'hd5b1;
29063: douta=16'hde54;
29064: douta=16'he6d7;
29065: douta=16'hf77a;
29066: douta=16'hf79a;
29067: douta=16'hf79a;
29068: douta=16'hef58;
29069: douta=16'heef6;
29070: douta=16'he6b5;
29071: douta=16'hddcf;
29072: douta=16'hd56e;
29073: douta=16'hd50b;
29074: douta=16'hc467;
29075: douta=16'hcc46;
29076: douta=16'hc425;
29077: douta=16'hc404;
29078: douta=16'hc405;
29079: douta=16'hcc25;
29080: douta=16'hcc47;
29081: douta=16'hcc47;
29082: douta=16'hcc68;
29083: douta=16'hcc68;
29084: douta=16'hcc68;
29085: douta=16'hcc67;
29086: douta=16'hcc68;
29087: douta=16'hcc68;
29088: douta=16'hcc68;
29089: douta=16'hcc68;
29090: douta=16'hd488;
29091: douta=16'hcc68;
29092: douta=16'hd468;
29093: douta=16'hcc68;
29094: douta=16'hd488;
29095: douta=16'hd488;
29096: douta=16'hd488;
29097: douta=16'hd488;
29098: douta=16'hd488;
29099: douta=16'hd488;
29100: douta=16'hd488;
29101: douta=16'hcc88;
29102: douta=16'hcc88;
29103: douta=16'hd488;
29104: douta=16'hd488;
29105: douta=16'hcc88;
29106: douta=16'hd488;
29107: douta=16'hd488;
29108: douta=16'hd489;
29109: douta=16'hd4a9;
29110: douta=16'hcc88;
29111: douta=16'hd488;
29112: douta=16'hd4a9;
29113: douta=16'hcc68;
29114: douta=16'hcc88;
29115: douta=16'hd488;
29116: douta=16'hd4a9;
29117: douta=16'hd488;
29118: douta=16'hcc67;
29119: douta=16'hd4c8;
29120: douta=16'hd4c9;
29121: douta=16'hd4c9;
29122: douta=16'hd468;
29123: douta=16'hac6f;
29124: douta=16'h9c91;
29125: douta=16'hacd2;
29126: douta=16'hb512;
29127: douta=16'hbd12;
29128: douta=16'hb513;
29129: douta=16'hb534;
29130: douta=16'hacf3;
29131: douta=16'h8c53;
29132: douta=16'h8433;
29133: douta=16'h7bf2;
29134: douta=16'h7bd1;
29135: douta=16'h6bb1;
29136: douta=16'h73b0;
29137: douta=16'h62cc;
29138: douta=16'h2903;
29139: douta=16'h3965;
29140: douta=16'h5226;
29141: douta=16'h41a5;
29142: douta=16'h5a68;
29143: douta=16'ha490;
29144: douta=16'h836c;
29145: douta=16'h836c;
29146: douta=16'h7b4b;
29147: douta=16'hacd1;
29148: douta=16'h9c4f;
29149: douta=16'ha46e;
29150: douta=16'ha46e;
29151: douta=16'ha46e;
29152: douta=16'h942d;
29153: douta=16'ha490;
29154: douta=16'hbd11;
29155: douta=16'hcdb3;
29156: douta=16'hcd93;
29157: douta=16'hcdb2;
29158: douta=16'hd5b3;
29159: douta=16'hd5d4;
29160: douta=16'hd5b3;
29161: douta=16'hc571;
29162: douta=16'hb4d0;
29163: douta=16'ha450;
29164: douta=16'h7bae;
29165: douta=16'h736e;
29166: douta=16'h4a6b;
29167: douta=16'h39e9;
29168: douta=16'h2146;
29169: douta=16'h2125;
29170: douta=16'h10c4;
29171: douta=16'h10a4;
29172: douta=16'h18e4;
29173: douta=16'h10a3;
29174: douta=16'h2168;
29175: douta=16'h1968;
29176: douta=16'h8ae7;
29177: douta=16'h82a7;
29178: douta=16'h82a7;
29179: douta=16'h82a7;
29180: douta=16'h82c7;
29181: douta=16'h82a7;
29182: douta=16'h8ac7;
29183: douta=16'h82a7;
29184: douta=16'had14;
29185: douta=16'hcdf6;
29186: douta=16'hc5b5;
29187: douta=16'hbd55;
29188: douta=16'h8c53;
29189: douta=16'ha557;
29190: douta=16'h94b4;
29191: douta=16'h9cd5;
29192: douta=16'h94d5;
29193: douta=16'h94b5;
29194: douta=16'h6b90;
29195: douta=16'h1060;
29196: douta=16'h20e3;
29197: douta=16'h28e3;
29198: douta=16'h20e3;
29199: douta=16'h20e3;
29200: douta=16'h20c3;
29201: douta=16'h20c3;
29202: douta=16'h20e3;
29203: douta=16'h20a2;
29204: douta=16'h1882;
29205: douta=16'h20a2;
29206: douta=16'h20a2;
29207: douta=16'h20a2;
29208: douta=16'h20a2;
29209: douta=16'h20a2;
29210: douta=16'h20c2;
29211: douta=16'h28e3;
29212: douta=16'h28e2;
29213: douta=16'h28e2;
29214: douta=16'h28e2;
29215: douta=16'h3123;
29216: douta=16'h3103;
29217: douta=16'h3923;
29218: douta=16'h422a;
29219: douta=16'h424a;
29220: douta=16'h18c5;
29221: douta=16'h5184;
29222: douta=16'h51a4;
29223: douta=16'h51a4;
29224: douta=16'h59c4;
29225: douta=16'h59c4;
29226: douta=16'h61e3;
29227: douta=16'h61a3;
29228: douta=16'hb594;
29229: douta=16'hacaf;
29230: douta=16'h7264;
29231: douta=16'h7244;
29232: douta=16'h7a85;
29233: douta=16'h7a85;
29234: douta=16'h7a85;
29235: douta=16'h7a64;
29236: douta=16'h6204;
29237: douta=16'h8244;
29238: douta=16'h7a24;
29239: douta=16'h82a5;
29240: douta=16'h82c6;
29241: douta=16'h9327;
29242: douta=16'ha40c;
29243: douta=16'hb4af;
29244: douta=16'hbd10;
29245: douta=16'hcdf3;
29246: douta=16'hde96;
29247: douta=16'he6f8;
29248: douta=16'hef59;
29249: douta=16'hf779;
29250: douta=16'hef37;
29251: douta=16'he6b5;
29252: douta=16'hde32;
29253: douta=16'hd5f0;
29254: douta=16'hcd2d;
29255: douta=16'hc4ca;
29256: douta=16'hc448;
29257: douta=16'hbc05;
29258: douta=16'hbbe5;
29259: douta=16'hbbc4;
29260: douta=16'hbbe5;
29261: douta=16'hc3e5;
29262: douta=16'hc405;
29263: douta=16'hc406;
29264: douta=16'hc427;
29265: douta=16'hcc47;
29266: douta=16'hcc48;
29267: douta=16'hcc47;
29268: douta=16'hcc47;
29269: douta=16'hcc46;
29270: douta=16'hcc47;
29271: douta=16'hcc48;
29272: douta=16'hcc67;
29273: douta=16'hcc47;
29274: douta=16'hcc67;
29275: douta=16'hcc68;
29276: douta=16'hcc48;
29277: douta=16'hcc68;
29278: douta=16'hcc68;
29279: douta=16'hcc68;
29280: douta=16'hcc68;
29281: douta=16'hcc67;
29282: douta=16'hcc68;
29283: douta=16'hcc68;
29284: douta=16'hcc88;
29285: douta=16'hcc68;
29286: douta=16'hcc68;
29287: douta=16'hd488;
29288: douta=16'hd488;
29289: douta=16'hd488;
29290: douta=16'hd488;
29291: douta=16'hd488;
29292: douta=16'hd488;
29293: douta=16'hd487;
29294: douta=16'hd488;
29295: douta=16'hd488;
29296: douta=16'hd488;
29297: douta=16'hcc88;
29298: douta=16'hd488;
29299: douta=16'hcc88;
29300: douta=16'hd488;
29301: douta=16'hd488;
29302: douta=16'hcc88;
29303: douta=16'hd488;
29304: douta=16'hd488;
29305: douta=16'hd4a9;
29306: douta=16'hcc68;
29307: douta=16'hd488;
29308: douta=16'hd488;
29309: douta=16'hd488;
29310: douta=16'hd487;
29311: douta=16'hcc25;
29312: douta=16'hcc25;
29313: douta=16'hcc45;
29314: douta=16'hcc87;
29315: douta=16'hccec;
29316: douta=16'ha490;
29317: douta=16'ha4b2;
29318: douta=16'hacd2;
29319: douta=16'hacd3;
29320: douta=16'ha4b3;
29321: douta=16'h9cb4;
29322: douta=16'h9494;
29323: douta=16'h8412;
29324: douta=16'h7bf2;
29325: douta=16'h8411;
29326: douta=16'h39a6;
29327: douta=16'h3944;
29328: douta=16'h28e3;
29329: douta=16'h4a05;
29330: douta=16'h72e9;
29331: douta=16'h6ae8;
29332: douta=16'h8bcc;
29333: douta=16'h8bcd;
29334: douta=16'h734a;
29335: douta=16'h41e6;
29336: douta=16'h9c6f;
29337: douta=16'h940d;
29338: douta=16'hb4f0;
29339: douta=16'h730b;
29340: douta=16'hc572;
29341: douta=16'hbd53;
29342: douta=16'hbd52;
29343: douta=16'hcd93;
29344: douta=16'hbd32;
29345: douta=16'hd5b3;
29346: douta=16'hd5b2;
29347: douta=16'hd5b3;
29348: douta=16'hd5b3;
29349: douta=16'hcd72;
29350: douta=16'hcd72;
29351: douta=16'hc532;
29352: douta=16'hc532;
29353: douta=16'hacb1;
29354: douta=16'hac91;
29355: douta=16'h8c10;
29356: douta=16'h9c71;
29357: douta=16'h8c10;
29358: douta=16'h6b4f;
29359: douta=16'h5b0d;
29360: douta=16'h3a2a;
29361: douta=16'h39e9;
29362: douta=16'h3a09;
29363: douta=16'h1906;
29364: douta=16'h10c4;
29365: douta=16'h1926;
29366: douta=16'h1128;
29367: douta=16'h3a6d;
29368: douta=16'h8aa6;
29369: douta=16'h8ac7;
29370: douta=16'h8ac7;
29371: douta=16'h8ac7;
29372: douta=16'h8ac7;
29373: douta=16'h8ac7;
29374: douta=16'h8ac7;
29375: douta=16'h8ae7;
29376: douta=16'had15;
29377: douta=16'hd616;
29378: douta=16'hc5b5;
29379: douta=16'hbd55;
29380: douta=16'h9494;
29381: douta=16'had57;
29382: douta=16'h9cd5;
29383: douta=16'h9cd5;
29384: douta=16'h94d5;
29385: douta=16'h8c74;
29386: douta=16'h4208;
29387: douta=16'h1040;
29388: douta=16'h28e3;
29389: douta=16'h20c3;
29390: douta=16'h20e3;
29391: douta=16'h20c3;
29392: douta=16'h20c3;
29393: douta=16'h20e3;
29394: douta=16'h20e3;
29395: douta=16'h20a3;
29396: douta=16'h1882;
29397: douta=16'h20a2;
29398: douta=16'h20a2;
29399: douta=16'h1881;
29400: douta=16'h20a2;
29401: douta=16'h20a2;
29402: douta=16'h28e2;
29403: douta=16'h28e3;
29404: douta=16'h28e2;
29405: douta=16'h28e2;
29406: douta=16'h30e2;
29407: douta=16'h3103;
29408: douta=16'h3903;
29409: douta=16'h3923;
29410: douta=16'h4a4b;
29411: douta=16'h3a09;
29412: douta=16'h18e5;
29413: douta=16'h5184;
29414: douta=16'h51a4;
29415: douta=16'h51a4;
29416: douta=16'h59c4;
29417: douta=16'h61e4;
29418: douta=16'h61e4;
29419: douta=16'h61c3;
29420: douta=16'hb594;
29421: douta=16'h9c2c;
29422: douta=16'h7a44;
29423: douta=16'h7224;
29424: douta=16'h7224;
29425: douta=16'h7203;
29426: douta=16'h7224;
29427: douta=16'h7224;
29428: douta=16'h7aa6;
29429: douta=16'h8b49;
29430: douta=16'h9beb;
29431: douta=16'hbd51;
29432: douta=16'hbd71;
29433: douta=16'hcdf3;
29434: douta=16'hdeb6;
29435: douta=16'hded6;
29436: douta=16'hded6;
29437: douta=16'hde95;
29438: douta=16'hde94;
29439: douta=16'hd631;
29440: douta=16'hc54d;
29441: douta=16'hc50c;
29442: douta=16'hc4aa;
29443: douta=16'hb3e7;
29444: douta=16'hb3c5;
29445: douta=16'hb3a4;
29446: douta=16'hb3a4;
29447: douta=16'hbba4;
29448: douta=16'hbbc4;
29449: douta=16'hc3e7;
29450: douta=16'hc3e7;
29451: douta=16'hc407;
29452: douta=16'hc406;
29453: douta=16'hc426;
29454: douta=16'hc426;
29455: douta=16'hc446;
29456: douta=16'hc446;
29457: douta=16'hc447;
29458: douta=16'hc446;
29459: douta=16'hcc48;
29460: douta=16'hcc47;
29461: douta=16'hcc47;
29462: douta=16'hcc67;
29463: douta=16'hcc47;
29464: douta=16'hcc67;
29465: douta=16'hcc68;
29466: douta=16'hcc67;
29467: douta=16'hcc48;
29468: douta=16'hcc68;
29469: douta=16'hcc68;
29470: douta=16'hcc88;
29471: douta=16'hcc68;
29472: douta=16'hcc88;
29473: douta=16'hcc67;
29474: douta=16'hd488;
29475: douta=16'hcc68;
29476: douta=16'hcc68;
29477: douta=16'hcc68;
29478: douta=16'hcc67;
29479: douta=16'hd488;
29480: douta=16'hd488;
29481: douta=16'hd488;
29482: douta=16'hcc67;
29483: douta=16'hd488;
29484: douta=16'hd488;
29485: douta=16'hd488;
29486: douta=16'hd488;
29487: douta=16'hd488;
29488: douta=16'hd488;
29489: douta=16'hd488;
29490: douta=16'hd488;
29491: douta=16'hd488;
29492: douta=16'hd488;
29493: douta=16'hd488;
29494: douta=16'hd488;
29495: douta=16'hcc88;
29496: douta=16'hd487;
29497: douta=16'hd467;
29498: douta=16'hcc25;
29499: douta=16'hcc46;
29500: douta=16'hcca9;
29501: douta=16'hccc9;
29502: douta=16'hcd0b;
29503: douta=16'hd58f;
29504: douta=16'hd5d0;
29505: douta=16'hde53;
29506: douta=16'heed7;
29507: douta=16'hffba;
29508: douta=16'he6d7;
29509: douta=16'ha492;
29510: douta=16'h9cb2;
29511: douta=16'ha4b3;
29512: douta=16'h9472;
29513: douta=16'h8c53;
29514: douta=16'h8c93;
29515: douta=16'h7bf2;
29516: douta=16'h738f;
29517: douta=16'h4a06;
29518: douta=16'h3124;
29519: douta=16'h41a5;
29520: douta=16'h5a68;
29521: douta=16'h7309;
29522: douta=16'h7b4a;
29523: douta=16'h7b2a;
29524: douta=16'h940d;
29525: douta=16'h940d;
29526: douta=16'ha46e;
29527: douta=16'h940e;
29528: douta=16'h6b0a;
29529: douta=16'h9c2e;
29530: douta=16'hde14;
29531: douta=16'h5a69;
29532: douta=16'hc573;
29533: douta=16'hc594;
29534: douta=16'hc573;
29535: douta=16'hbd12;
29536: douta=16'hbcf2;
29537: douta=16'ha471;
29538: douta=16'hb4f2;
29539: douta=16'hb4d2;
29540: douta=16'hb4d2;
29541: douta=16'hb4d2;
29542: douta=16'hacd2;
29543: douta=16'hacd2;
29544: douta=16'hacd3;
29545: douta=16'h9c71;
29546: douta=16'ha472;
29547: douta=16'h8c10;
29548: douta=16'h9451;
29549: douta=16'h8c11;
29550: douta=16'h73b0;
29551: douta=16'h6b6f;
29552: douta=16'h4a6c;
29553: douta=16'h3a4a;
29554: douta=16'h39e9;
29555: douta=16'h2188;
29556: douta=16'h2167;
29557: douta=16'h1905;
29558: douta=16'h1106;
29559: douta=16'h08e6;
29560: douta=16'h82a8;
29561: douta=16'h8ac7;
29562: douta=16'h8ae7;
29563: douta=16'h8b08;
29564: douta=16'h8ae7;
29565: douta=16'h8ac7;
29566: douta=16'h8ae7;
29567: douta=16'h8ae7;
29568: douta=16'had36;
29569: douta=16'hcdf6;
29570: douta=16'hc5b5;
29571: douta=16'had15;
29572: douta=16'had77;
29573: douta=16'ha516;
29574: douta=16'h9cf5;
29575: douta=16'h9cd5;
29576: douta=16'h8c74;
29577: douta=16'h8454;
29578: douta=16'h3a2a;
29579: douta=16'h4aac;
29580: douta=16'h39c8;
29581: douta=16'h20a2;
29582: douta=16'h20c2;
29583: douta=16'h20c3;
29584: douta=16'h20c3;
29585: douta=16'h28e3;
29586: douta=16'h20e3;
29587: douta=16'h1882;
29588: douta=16'h18a2;
29589: douta=16'h20a2;
29590: douta=16'h18a2;
29591: douta=16'h20c2;
29592: douta=16'h20a2;
29593: douta=16'h20c2;
29594: douta=16'h20c2;
29595: douta=16'h28e3;
29596: douta=16'h28e2;
29597: douta=16'h30e2;
29598: douta=16'h30e2;
29599: douta=16'h3103;
29600: douta=16'h3103;
29601: douta=16'h30e2;
29602: douta=16'h422a;
29603: douta=16'h2947;
29604: douta=16'h28e4;
29605: douta=16'h5184;
29606: douta=16'h51c4;
29607: douta=16'h5a05;
29608: douta=16'h7308;
29609: douta=16'h836a;
29610: douta=16'h93ec;
29611: douta=16'hb530;
29612: douta=16'hbd91;
29613: douta=16'hc5f3;
29614: douta=16'hce33;
29615: douta=16'hcdf2;
29616: douta=16'hc591;
29617: douta=16'hacee;
29618: douta=16'hac8d;
29619: douta=16'ha40b;
29620: douta=16'h9bea;
29621: douta=16'h49c4;
29622: douta=16'h9327;
29623: douta=16'h8284;
29624: douta=16'h8283;
29625: douta=16'h8284;
29626: douta=16'h8aa4;
29627: douta=16'h92c6;
29628: douta=16'h9306;
29629: douta=16'h9b26;
29630: douta=16'ha366;
29631: douta=16'ha386;
29632: douta=16'hab86;
29633: douta=16'hb3a6;
29634: douta=16'hb3a6;
29635: douta=16'hb3c6;
29636: douta=16'hbbc6;
29637: douta=16'hbbe6;
29638: douta=16'hbbe6;
29639: douta=16'hbbe6;
29640: douta=16'hbc06;
29641: douta=16'hc427;
29642: douta=16'hc427;
29643: douta=16'hc407;
29644: douta=16'hc427;
29645: douta=16'hcc47;
29646: douta=16'hc427;
29647: douta=16'hc426;
29648: douta=16'hc427;
29649: douta=16'hcc47;
29650: douta=16'hcc47;
29651: douta=16'hcc47;
29652: douta=16'hcc47;
29653: douta=16'hc447;
29654: douta=16'hcc47;
29655: douta=16'hcc48;
29656: douta=16'hcc67;
29657: douta=16'hcc68;
29658: douta=16'hcc47;
29659: douta=16'hcc68;
29660: douta=16'hcc68;
29661: douta=16'hcc69;
29662: douta=16'hcc88;
29663: douta=16'hcc88;
29664: douta=16'hcc67;
29665: douta=16'hcc68;
29666: douta=16'hd488;
29667: douta=16'hd488;
29668: douta=16'hcc67;
29669: douta=16'hcc68;
29670: douta=16'hcc87;
29671: douta=16'hd467;
29672: douta=16'hcc66;
29673: douta=16'hd446;
29674: douta=16'hcc45;
29675: douta=16'hcc25;
29676: douta=16'hcc45;
29677: douta=16'hcca9;
29678: douta=16'hcccb;
29679: douta=16'hd52d;
29680: douta=16'hddb1;
29681: douta=16'hde33;
29682: douta=16'he675;
29683: douta=16'hef18;
29684: douta=16'hf77b;
29685: douta=16'hf7bc;
29686: douta=16'hfffc;
29687: douta=16'hffdc;
29688: douta=16'hff9a;
29689: douta=16'hef17;
29690: douta=16'hf6d6;
29691: douta=16'hf75a;
29692: douta=16'hd50b;
29693: douta=16'hd50a;
29694: douta=16'hd4c9;
29695: douta=16'hcc67;
29696: douta=16'hcc46;
29697: douta=16'hcc47;
29698: douta=16'hd468;
29699: douta=16'hd447;
29700: douta=16'hcc68;
29701: douta=16'ha492;
29702: douta=16'h9472;
29703: douta=16'h8411;
29704: douta=16'h734e;
29705: douta=16'h5226;
29706: douta=16'h3163;
29707: douta=16'h5a68;
29708: douta=16'h732b;
29709: douta=16'h7b4b;
29710: douta=16'h7b4b;
29711: douta=16'h836b;
29712: douta=16'h9c4e;
29713: douta=16'ha44e;
29714: douta=16'ha46e;
29715: douta=16'hac8f;
29716: douta=16'hc531;
29717: douta=16'h940e;
29718: douta=16'hd5b3;
29719: douta=16'hc552;
29720: douta=16'hde16;
29721: douta=16'hd5b3;
29722: douta=16'h6b6f;
29723: douta=16'ha491;
29724: douta=16'h8390;
29725: douta=16'ha4b3;
29726: douta=16'ha473;
29727: douta=16'h9c72;
29728: douta=16'h8412;
29729: douta=16'h73b0;
29730: douta=16'h6b4f;
29731: douta=16'h7bd1;
29732: douta=16'h7bf1;
29733: douta=16'h8453;
29734: douta=16'h8453;
29735: douta=16'h8c94;
29736: douta=16'h8c75;
29737: douta=16'h9474;
29738: douta=16'h8c53;
29739: douta=16'h8c73;
29740: douta=16'h83f1;
29741: douta=16'h8c52;
29742: douta=16'h8c74;
29743: douta=16'h7c13;
29744: douta=16'h7c54;
29745: douta=16'h73f3;
29746: douta=16'h320a;
29747: douta=16'h3a2b;
29748: douta=16'h2947;
29749: douta=16'h2125;
29750: douta=16'h428b;
29751: douta=16'hb5b6;
29752: douta=16'h61c4;
29753: douta=16'h9309;
29754: douta=16'h92e8;
29755: douta=16'h9307;
29756: douta=16'h9307;
29757: douta=16'h9307;
29758: douta=16'h9308;
29759: douta=16'h9308;
29760: douta=16'had36;
29761: douta=16'hc5b5;
29762: douta=16'hbd95;
29763: douta=16'h9c94;
29764: douta=16'had57;
29765: douta=16'h9cf5;
29766: douta=16'h9cd5;
29767: douta=16'h9cd5;
29768: douta=16'h8433;
29769: douta=16'h94d7;
29770: douta=16'h20c3;
29771: douta=16'h20c3;
29772: douta=16'h2904;
29773: douta=16'h426b;
29774: douta=16'h426b;
29775: douta=16'h3a29;
29776: douta=16'h20c2;
29777: douta=16'h20a2;
29778: douta=16'h20e3;
29779: douta=16'h2082;
29780: douta=16'h20a2;
29781: douta=16'h1881;
29782: douta=16'h1881;
29783: douta=16'h1861;
29784: douta=16'h1881;
29785: douta=16'h2082;
29786: douta=16'h2082;
29787: douta=16'h28e3;
29788: douta=16'h3144;
29789: douta=16'h3965;
29790: douta=16'h41a5;
29791: douta=16'h5248;
29792: douta=16'h62c9;
29793: douta=16'h736c;
29794: douta=16'h39c8;
29795: douta=16'h1906;
29796: douta=16'h7b6c;
29797: douta=16'h948f;
29798: douta=16'h944e;
29799: douta=16'h942e;
29800: douta=16'h834a;
29801: douta=16'h7b29;
29802: douta=16'h72c7;
29803: douta=16'h6a45;
29804: douta=16'h7224;
29805: douta=16'h7224;
29806: douta=16'h7204;
29807: douta=16'h7203;
29808: douta=16'h7244;
29809: douta=16'h7a65;
29810: douta=16'h8285;
29811: douta=16'h82a5;
29812: douta=16'h82c5;
29813: douta=16'h51a4;
29814: douta=16'h7a65;
29815: douta=16'h8ae5;
29816: douta=16'h92e5;
29817: douta=16'h92c6;
29818: douta=16'h9306;
29819: douta=16'h9306;
29820: douta=16'h9306;
29821: douta=16'h9b46;
29822: douta=16'ha366;
29823: douta=16'hab87;
29824: douta=16'hab86;
29825: douta=16'hb3a6;
29826: douta=16'hb3a7;
29827: douta=16'hb3c7;
29828: douta=16'hbbe7;
29829: douta=16'hbbe7;
29830: douta=16'hbbe7;
29831: douta=16'hbbe6;
29832: douta=16'hc407;
29833: douta=16'hbc07;
29834: douta=16'hc407;
29835: douta=16'hc407;
29836: douta=16'hc426;
29837: douta=16'hc426;
29838: douta=16'hc427;
29839: douta=16'hc427;
29840: douta=16'hcc47;
29841: douta=16'hcc27;
29842: douta=16'hcc47;
29843: douta=16'hcc47;
29844: douta=16'hcc47;
29845: douta=16'hcc48;
29846: douta=16'hcc67;
29847: douta=16'hcc67;
29848: douta=16'hcc47;
29849: douta=16'hcc48;
29850: douta=16'hcc68;
29851: douta=16'hcc67;
29852: douta=16'hcc67;
29853: douta=16'hcc67;
29854: douta=16'hcc25;
29855: douta=16'hcc25;
29856: douta=16'hcc25;
29857: douta=16'hcc46;
29858: douta=16'hcc68;
29859: douta=16'hcca9;
29860: douta=16'hd52c;
29861: douta=16'hdd8f;
29862: douta=16'hde13;
29863: douta=16'he6b7;
29864: douta=16'heef8;
29865: douta=16'hf75a;
29866: douta=16'hf7bd;
29867: douta=16'hffdc;
29868: douta=16'hffdc;
29869: douta=16'hf77a;
29870: douta=16'hf738;
29871: douta=16'heed6;
29872: douta=16'he653;
29873: douta=16'hddcf;
29874: douta=16'hdd8f;
29875: douta=16'hd50b;
29876: douta=16'hcca9;
29877: douta=16'hcc67;
29878: douta=16'hcc46;
29879: douta=16'hcc26;
29880: douta=16'hcc66;
29881: douta=16'hd425;
29882: douta=16'had11;
29883: douta=16'hde97;
29884: douta=16'hd489;
29885: douta=16'hd4a9;
29886: douta=16'hd488;
29887: douta=16'hcc88;
29888: douta=16'hcc88;
29889: douta=16'hd489;
29890: douta=16'hcc69;
29891: douta=16'hcc68;
29892: douta=16'hdc87;
29893: douta=16'h83ae;
29894: douta=16'h62aa;
29895: douta=16'h4185;
29896: douta=16'h62a8;
29897: douta=16'h730a;
29898: douta=16'h7b4b;
29899: douta=16'h7b6b;
29900: douta=16'h8c0e;
29901: douta=16'h8c0d;
29902: douta=16'ha48f;
29903: douta=16'hacaf;
29904: douta=16'hb4f0;
29905: douta=16'hbd10;
29906: douta=16'hcd73;
29907: douta=16'hcdb4;
29908: douta=16'hacb0;
29909: douta=16'h8bad;
29910: douta=16'hddd4;
29911: douta=16'hcd93;
29912: douta=16'hacb3;
29913: douta=16'h9c52;
29914: douta=16'h8412;
29915: douta=16'h7390;
29916: douta=16'ha4b2;
29917: douta=16'h9452;
29918: douta=16'h8c32;
29919: douta=16'h83f1;
29920: douta=16'h7bb1;
29921: douta=16'h7390;
29922: douta=16'h6b4f;
29923: douta=16'h736f;
29924: douta=16'h738f;
29925: douta=16'h7390;
29926: douta=16'h7390;
29927: douta=16'h6b4f;
29928: douta=16'h736f;
29929: douta=16'h6b6f;
29930: douta=16'h73b1;
29931: douta=16'h73b0;
29932: douta=16'h73b1;
29933: douta=16'h6b70;
29934: douta=16'h7c12;
29935: douta=16'h7433;
29936: douta=16'h6370;
29937: douta=16'h6391;
29938: douta=16'h6350;
29939: douta=16'h3a2a;
29940: douta=16'h2147;
29941: douta=16'h2a4c;
29942: douta=16'hffff;
29943: douta=16'hffff;
29944: douta=16'h938e;
29945: douta=16'h9b49;
29946: douta=16'h9328;
29947: douta=16'h9307;
29948: douta=16'h9328;
29949: douta=16'h9307;
29950: douta=16'h9b28;
29951: douta=16'h9328;
29952: douta=16'hb556;
29953: douta=16'hcdb5;
29954: douta=16'hbd75;
29955: douta=16'h8c53;
29956: douta=16'ha516;
29957: douta=16'ha4f5;
29958: douta=16'h9cd5;
29959: douta=16'h9cb5;
29960: douta=16'h8c74;
29961: douta=16'h9d79;
29962: douta=16'h28e3;
29963: douta=16'h28e3;
29964: douta=16'h20a2;
29965: douta=16'h2924;
29966: douta=16'h320a;
29967: douta=16'h428c;
29968: douta=16'h3a4a;
29969: douta=16'h2925;
29970: douta=16'h2082;
29971: douta=16'h1881;
29972: douta=16'h1881;
29973: douta=16'h1881;
29974: douta=16'h20a3;
29975: douta=16'h2904;
29976: douta=16'h2924;
29977: douta=16'h39a6;
29978: douta=16'h39a7;
29979: douta=16'h4a29;
29980: douta=16'h52aa;
29981: douta=16'h630b;
29982: douta=16'h630b;
29983: douta=16'h734b;
29984: douta=16'h734b;
29985: douta=16'h734b;
29986: douta=16'h39c9;
29987: douta=16'h10e6;
29988: douta=16'h6247;
29989: douta=16'h5a25;
29990: douta=16'h5a05;
29991: douta=16'h59c4;
29992: douta=16'h59a3;
29993: douta=16'h59a3;
29994: douta=16'h61c4;
29995: douta=16'h69e3;
29996: douta=16'h7224;
29997: douta=16'h7244;
29998: douta=16'h7a64;
29999: douta=16'h7a64;
30000: douta=16'h8285;
30001: douta=16'h82a5;
30002: douta=16'h8285;
30003: douta=16'h82a5;
30004: douta=16'h8ac5;
30005: douta=16'h51c4;
30006: douta=16'h6a25;
30007: douta=16'h8ae5;
30008: douta=16'h9306;
30009: douta=16'h8ac5;
30010: douta=16'h92e6;
30011: douta=16'h9306;
30012: douta=16'h9326;
30013: douta=16'h9b46;
30014: douta=16'ha366;
30015: douta=16'hab87;
30016: douta=16'haba6;
30017: douta=16'haba6;
30018: douta=16'hb3c7;
30019: douta=16'hb3e6;
30020: douta=16'hbbe7;
30021: douta=16'hbbe6;
30022: douta=16'hbbe6;
30023: douta=16'hc3e7;
30024: douta=16'hc406;
30025: douta=16'hc427;
30026: douta=16'hc407;
30027: douta=16'hc427;
30028: douta=16'hcc27;
30029: douta=16'hc427;
30030: douta=16'hc427;
30031: douta=16'hcc47;
30032: douta=16'hcc47;
30033: douta=16'hcc47;
30034: douta=16'hcc47;
30035: douta=16'hcc48;
30036: douta=16'hcc47;
30037: douta=16'hcc47;
30038: douta=16'hcc47;
30039: douta=16'hcc47;
30040: douta=16'hc404;
30041: douta=16'hcc05;
30042: douta=16'hc403;
30043: douta=16'hcc25;
30044: douta=16'hc445;
30045: douta=16'hcc47;
30046: douta=16'hd52d;
30047: douta=16'hd56e;
30048: douta=16'hddd1;
30049: douta=16'hde74;
30050: douta=16'heed8;
30051: douta=16'hef19;
30052: douta=16'hf77c;
30053: douta=16'hffbc;
30054: douta=16'hffdc;
30055: douta=16'hf79a;
30056: douta=16'hf77a;
30057: douta=16'hef17;
30058: douta=16'he674;
30059: douta=16'he611;
30060: douta=16'hddef;
30061: douta=16'hd52c;
30062: douta=16'hd50b;
30063: douta=16'hcca9;
30064: douta=16'hcc67;
30065: douta=16'hcc46;
30066: douta=16'hcc47;
30067: douta=16'hcc47;
30068: douta=16'hd468;
30069: douta=16'hd468;
30070: douta=16'hd488;
30071: douta=16'hcc88;
30072: douta=16'hd488;
30073: douta=16'hd466;
30074: douta=16'had31;
30075: douta=16'hdeb8;
30076: douta=16'hcc68;
30077: douta=16'hd4a9;
30078: douta=16'hcc89;
30079: douta=16'hcc68;
30080: douta=16'hcc88;
30081: douta=16'hcc68;
30082: douta=16'hcc69;
30083: douta=16'hcc49;
30084: douta=16'hd468;
30085: douta=16'h49c5;
30086: douta=16'h4184;
30087: douta=16'h5227;
30088: douta=16'h838c;
30089: douta=16'h838c;
30090: douta=16'h8bcc;
30091: douta=16'h940d;
30092: douta=16'h9c8f;
30093: douta=16'h944e;
30094: douta=16'hbd30;
30095: douta=16'hbd10;
30096: douta=16'hbd11;
30097: douta=16'hc572;
30098: douta=16'hcd93;
30099: douta=16'hd5f4;
30100: douta=16'hcd93;
30101: douta=16'h940f;
30102: douta=16'hbd12;
30103: douta=16'hcd72;
30104: douta=16'ha492;
30105: douta=16'h9c92;
30106: douta=16'h8433;
30107: douta=16'h73b0;
30108: douta=16'h6b6f;
30109: douta=16'h83f1;
30110: douta=16'h8411;
30111: douta=16'h83d1;
30112: douta=16'h7bb1;
30113: douta=16'h6b4f;
30114: douta=16'h6b4f;
30115: douta=16'h6b4e;
30116: douta=16'h6b2e;
30117: douta=16'h6b4f;
30118: douta=16'h6b4e;
30119: douta=16'h6b0d;
30120: douta=16'h5a8b;
30121: douta=16'h6b2e;
30122: douta=16'h6b4f;
30123: douta=16'h6b4f;
30124: douta=16'h6b6f;
30125: douta=16'h6b4f;
30126: douta=16'h6370;
30127: douta=16'h7413;
30128: douta=16'h73f3;
30129: douta=16'h6391;
30130: douta=16'h7bf1;
30131: douta=16'h424c;
30132: douta=16'h2967;
30133: douta=16'h5b6e;
30134: douta=16'hffff;
30135: douta=16'hffff;
30136: douta=16'hd5b6;
30137: douta=16'h9309;
30138: douta=16'h9b28;
30139: douta=16'h9328;
30140: douta=16'h9b28;
30141: douta=16'h9b28;
30142: douta=16'h9b28;
30143: douta=16'h9b28;
30144: douta=16'hd5f6;
30145: douta=16'hc596;
30146: douta=16'had15;
30147: douta=16'h9cb4;
30148: douta=16'ha4f5;
30149: douta=16'ha4f5;
30150: douta=16'h9cd5;
30151: douta=16'h8434;
30152: douta=16'h94d6;
30153: douta=16'h3166;
30154: douta=16'h20e3;
30155: douta=16'h20e3;
30156: douta=16'h20c3;
30157: douta=16'h28e3;
30158: douta=16'h20e3;
30159: douta=16'h20c3;
30160: douta=16'h20a3;
30161: douta=16'h20c3;
30162: douta=16'h20e3;
30163: douta=16'h2103;
30164: douta=16'h2103;
30165: douta=16'h20a3;
30166: douta=16'h20c3;
30167: douta=16'h20a2;
30168: douta=16'h20a2;
30169: douta=16'h20a2;
30170: douta=16'h28a2;
30171: douta=16'h28c2;
30172: douta=16'h28c2;
30173: douta=16'h30e2;
30174: douta=16'h3102;
30175: douta=16'h3903;
30176: douta=16'h4123;
30177: douta=16'h4123;
30178: douta=16'h2947;
30179: douta=16'h0884;
30180: douta=16'h5184;
30181: douta=16'h59c4;
30182: douta=16'h59c4;
30183: douta=16'h59c4;
30184: douta=16'h61e4;
30185: douta=16'h6204;
30186: douta=16'h6a24;
30187: douta=16'h7224;
30188: douta=16'h7244;
30189: douta=16'h7a65;
30190: douta=16'h7a64;
30191: douta=16'h7a85;
30192: douta=16'h7a85;
30193: douta=16'h8285;
30194: douta=16'h82a6;
30195: douta=16'h8aa6;
30196: douta=16'h82c6;
30197: douta=16'h7a85;
30198: douta=16'h5184;
30199: douta=16'h8ac5;
30200: douta=16'h9306;
30201: douta=16'h9306;
30202: douta=16'h9306;
30203: douta=16'h9306;
30204: douta=16'h9326;
30205: douta=16'h9b26;
30206: douta=16'ha366;
30207: douta=16'hab87;
30208: douta=16'hb3c6;
30209: douta=16'hb3a6;
30210: douta=16'hb3c6;
30211: douta=16'hb3c7;
30212: douta=16'hbbe6;
30213: douta=16'hb3c6;
30214: douta=16'hbbe6;
30215: douta=16'hbbe6;
30216: douta=16'hbbc5;
30217: douta=16'hbba4;
30218: douta=16'hc3c4;
30219: douta=16'hbbc4;
30220: douta=16'hc426;
30221: douta=16'hc468;
30222: douta=16'hc4a9;
30223: douta=16'hd58f;
30224: douta=16'hd5d1;
30225: douta=16'hde54;
30226: douta=16'heef8;
30227: douta=16'hef59;
30228: douta=16'hf77a;
30229: douta=16'hf7bc;
30230: douta=16'hf7bb;
30231: douta=16'hf77a;
30232: douta=16'heef6;
30233: douta=16'he6b6;
30234: douta=16'he673;
30235: douta=16'hddaf;
30236: douta=16'hd54d;
30237: douta=16'hd52b;
30238: douta=16'hcca8;
30239: douta=16'hcc88;
30240: douta=16'hcc46;
30241: douta=16'hcc25;
30242: douta=16'hcc46;
30243: douta=16'hcc46;
30244: douta=16'hcc47;
30245: douta=16'hcc68;
30246: douta=16'hd488;
30247: douta=16'hcc88;
30248: douta=16'hcc88;
30249: douta=16'hcc88;
30250: douta=16'hd488;
30251: douta=16'hcc88;
30252: douta=16'hcc88;
30253: douta=16'hcc88;
30254: douta=16'hd488;
30255: douta=16'hcc88;
30256: douta=16'hd4a9;
30257: douta=16'hcc68;
30258: douta=16'hd469;
30259: douta=16'hd488;
30260: douta=16'hcc69;
30261: douta=16'hd488;
30262: douta=16'hd488;
30263: douta=16'hd488;
30264: douta=16'hd4a9;
30265: douta=16'hd487;
30266: douta=16'had11;
30267: douta=16'hdeb8;
30268: douta=16'hcc88;
30269: douta=16'hcc88;
30270: douta=16'hcc88;
30271: douta=16'hcc68;
30272: douta=16'hcc68;
30273: douta=16'hcc68;
30274: douta=16'hcc68;
30275: douta=16'hcc69;
30276: douta=16'hcc68;
30277: douta=16'h730a;
30278: douta=16'h8bac;
30279: douta=16'h8bee;
30280: douta=16'hacb0;
30281: douta=16'hac90;
30282: douta=16'ha490;
30283: douta=16'hc552;
30284: douta=16'hbd11;
30285: douta=16'hc553;
30286: douta=16'hcdb4;
30287: douta=16'hd5d4;
30288: douta=16'hd5b4;
30289: douta=16'hc573;
30290: douta=16'hbd12;
30291: douta=16'hacd3;
30292: douta=16'h8c12;
30293: douta=16'h8bf1;
30294: douta=16'h9452;
30295: douta=16'h83b0;
30296: douta=16'h8c53;
30297: douta=16'h9474;
30298: douta=16'h7bf2;
30299: douta=16'h7390;
30300: douta=16'h632f;
30301: douta=16'h6b2e;
30302: douta=16'h734f;
30303: douta=16'h630d;
30304: douta=16'h630e;
30305: douta=16'h6b2e;
30306: douta=16'h630e;
30307: douta=16'h5acd;
30308: douta=16'h528c;
30309: douta=16'h734f;
30310: douta=16'h62cd;
30311: douta=16'h62ed;
30312: douta=16'h5a6b;
30313: douta=16'h528a;
30314: douta=16'h49e9;
30315: douta=16'h7b6f;
30316: douta=16'h62ac;
30317: douta=16'h62ed;
30318: douta=16'h5b0e;
30319: douta=16'h320b;
30320: douta=16'h8433;
30321: douta=16'h7390;
30322: douta=16'h6bb3;
30323: douta=16'h5b72;
30324: douta=16'h53d3;
30325: douta=16'hffff;
30326: douta=16'hfeba;
30327: douta=16'hee58;
30328: douta=16'hab49;
30329: douta=16'ha349;
30330: douta=16'h9b29;
30331: douta=16'h9b48;
30332: douta=16'h9b48;
30333: douta=16'h9b48;
30334: douta=16'h9b48;
30335: douta=16'h9b48;
30336: douta=16'hde16;
30337: douta=16'hbd55;
30338: douta=16'h9494;
30339: douta=16'had36;
30340: douta=16'ha515;
30341: douta=16'ha4f5;
30342: douta=16'h9cd5;
30343: douta=16'h8cb6;
30344: douta=16'h31c7;
30345: douta=16'h1040;
30346: douta=16'h28e3;
30347: douta=16'h28e3;
30348: douta=16'h28e3;
30349: douta=16'h28e3;
30350: douta=16'h20e3;
30351: douta=16'h20e3;
30352: douta=16'h20e3;
30353: douta=16'h20e3;
30354: douta=16'h20e3;
30355: douta=16'h20a2;
30356: douta=16'h20a2;
30357: douta=16'h20a2;
30358: douta=16'h20a2;
30359: douta=16'h20a2;
30360: douta=16'h20a2;
30361: douta=16'h28e2;
30362: douta=16'h28e3;
30363: douta=16'h30e3;
30364: douta=16'h3103;
30365: douta=16'h3123;
30366: douta=16'h3903;
30367: douta=16'h4123;
30368: douta=16'h4144;
30369: douta=16'h4165;
30370: douta=16'h2126;
30371: douta=16'h18a5;
30372: douta=16'h59a4;
30373: douta=16'h51a4;
30374: douta=16'h61e4;
30375: douta=16'h61c4;
30376: douta=16'h6204;
30377: douta=16'h6a04;
30378: douta=16'h6a04;
30379: douta=16'h7244;
30380: douta=16'h7a64;
30381: douta=16'h7a64;
30382: douta=16'h7a85;
30383: douta=16'h8286;
30384: douta=16'h82a5;
30385: douta=16'h82a6;
30386: douta=16'h82a5;
30387: douta=16'h82c6;
30388: douta=16'h8ac6;
30389: douta=16'h9326;
30390: douta=16'h61e5;
30391: douta=16'h9306;
30392: douta=16'h9306;
30393: douta=16'h9305;
30394: douta=16'h92e6;
30395: douta=16'h9326;
30396: douta=16'h9306;
30397: douta=16'h9b05;
30398: douta=16'ha326;
30399: douta=16'ha325;
30400: douta=16'hab45;
30401: douta=16'hab64;
30402: douta=16'hab85;
30403: douta=16'hbc08;
30404: douta=16'hc4ac;
30405: douta=16'hc50d;
30406: douta=16'hd5b1;
30407: douta=16'hde53;
30408: douta=16'he6d6;
30409: douta=16'hef7a;
30410: douta=16'hf77a;
30411: douta=16'hf7bb;
30412: douta=16'hf77a;
30413: douta=16'hef38;
30414: douta=16'heef6;
30415: douta=16'hde32;
30416: douta=16'hddf1;
30417: douta=16'hd58e;
30418: douta=16'hccea;
30419: douta=16'hcca8;
30420: douta=16'hc468;
30421: douta=16'hc425;
30422: douta=16'hcc25;
30423: douta=16'hcc25;
30424: douta=16'hcc46;
30425: douta=16'hcc46;
30426: douta=16'hcc67;
30427: douta=16'hcc68;
30428: douta=16'hcc67;
30429: douta=16'hcc68;
30430: douta=16'hd488;
30431: douta=16'hcc67;
30432: douta=16'hcc68;
30433: douta=16'hcc68;
30434: douta=16'hd488;
30435: douta=16'hcc68;
30436: douta=16'hcc68;
30437: douta=16'hcc88;
30438: douta=16'hcc88;
30439: douta=16'hcc88;
30440: douta=16'hcc88;
30441: douta=16'hd488;
30442: douta=16'hcc88;
30443: douta=16'hcc88;
30444: douta=16'hcc88;
30445: douta=16'hd4a9;
30446: douta=16'hcc88;
30447: douta=16'hd4a9;
30448: douta=16'hcc88;
30449: douta=16'hd4a9;
30450: douta=16'hd489;
30451: douta=16'hd489;
30452: douta=16'hd4a9;
30453: douta=16'hd4a9;
30454: douta=16'hd4a9;
30455: douta=16'hd488;
30456: douta=16'hd488;
30457: douta=16'hd487;
30458: douta=16'had31;
30459: douta=16'hded7;
30460: douta=16'hcc68;
30461: douta=16'hcc68;
30462: douta=16'hcc88;
30463: douta=16'hcc88;
30464: douta=16'hcc88;
30465: douta=16'hcc88;
30466: douta=16'hd488;
30467: douta=16'hcc68;
30468: douta=16'hcc88;
30469: douta=16'h8bad;
30470: douta=16'h8bcd;
30471: douta=16'h93ee;
30472: douta=16'hbd32;
30473: douta=16'hbd12;
30474: douta=16'hbd33;
30475: douta=16'hc573;
30476: douta=16'hbd73;
30477: douta=16'hcdb5;
30478: douta=16'hd5d4;
30479: douta=16'hcd92;
30480: douta=16'hcd73;
30481: douta=16'hb4d3;
30482: douta=16'h8c32;
30483: douta=16'h9453;
30484: douta=16'h9473;
30485: douta=16'h8c32;
30486: douta=16'h7bb0;
30487: douta=16'h6b4f;
30488: douta=16'h7bb0;
30489: douta=16'h732f;
30490: douta=16'h6b2e;
30491: douta=16'h630e;
30492: douta=16'h632e;
30493: douta=16'h8432;
30494: douta=16'h736f;
30495: douta=16'h62ed;
30496: douta=16'h4a2a;
30497: douta=16'h5acc;
30498: douta=16'h62cc;
30499: douta=16'h5a8b;
30500: douta=16'h526a;
30501: douta=16'h41e8;
30502: douta=16'h736f;
30503: douta=16'h8c32;
30504: douta=16'h9453;
30505: douta=16'h8c74;
30506: douta=16'h8432;
30507: douta=16'h6b4f;
30508: douta=16'h6b2e;
30509: douta=16'h634e;
30510: douta=16'h9c92;
30511: douta=16'ha575;
30512: douta=16'h6c94;
30513: douta=16'h8557;
30514: douta=16'hcdb3;
30515: douta=16'hddb2;
30516: douta=16'hc388;
30517: douta=16'h9ac4;
30518: douta=16'ha368;
30519: douta=16'ha368;
30520: douta=16'h9b47;
30521: douta=16'ha369;
30522: douta=16'ha369;
30523: douta=16'h9b48;
30524: douta=16'h9b48;
30525: douta=16'h9b48;
30526: douta=16'h9b48;
30527: douta=16'h9b48;
30528: douta=16'hd616;
30529: douta=16'hbd96;
30530: douta=16'h8433;
30531: douta=16'hb577;
30532: douta=16'ha4f5;
30533: douta=16'h9cf5;
30534: douta=16'ha4d5;
30535: douta=16'ha539;
30536: douta=16'h1881;
30537: douta=16'h28e3;
30538: douta=16'h28e3;
30539: douta=16'h28e3;
30540: douta=16'h20e3;
30541: douta=16'h20c3;
30542: douta=16'h20c3;
30543: douta=16'h28e3;
30544: douta=16'h20e3;
30545: douta=16'h20c3;
30546: douta=16'h20e3;
30547: douta=16'h20c2;
30548: douta=16'h2082;
30549: douta=16'h20a2;
30550: douta=16'h20a2;
30551: douta=16'h20a2;
30552: douta=16'h20a2;
30553: douta=16'h28e3;
30554: douta=16'h28e3;
30555: douta=16'h30e3;
30556: douta=16'h3123;
30557: douta=16'h3103;
30558: douta=16'h3923;
30559: douta=16'h4143;
30560: douta=16'h4143;
30561: douta=16'h4185;
30562: douta=16'h1905;
30563: douta=16'h20c5;
30564: douta=16'h51a4;
30565: douta=16'h59e4;
30566: douta=16'h59c4;
30567: douta=16'h61c4;
30568: douta=16'h61e4;
30569: douta=16'h69e4;
30570: douta=16'h6a04;
30571: douta=16'h7244;
30572: douta=16'h7a65;
30573: douta=16'h7a65;
30574: douta=16'h7a85;
30575: douta=16'h82a5;
30576: douta=16'h8285;
30577: douta=16'h8aa6;
30578: douta=16'h8aa6;
30579: douta=16'h82c6;
30580: douta=16'h8ac6;
30581: douta=16'h9306;
30582: douta=16'h6a25;
30583: douta=16'h8ac4;
30584: douta=16'h8ac4;
30585: douta=16'h8aa4;
30586: douta=16'h8a84;
30587: douta=16'h8aa5;
30588: douta=16'h8ac6;
30589: douta=16'h9b67;
30590: douta=16'ha3e8;
30591: douta=16'hb46b;
30592: douta=16'hcd4f;
30593: douta=16'hcd90;
30594: douta=16'hde13;
30595: douta=16'he6b6;
30596: douta=16'hef38;
30597: douta=16'hef59;
30598: douta=16'hf77a;
30599: douta=16'hef59;
30600: douta=16'heef7;
30601: douta=16'he653;
30602: douta=16'hde32;
30603: douta=16'hd5d0;
30604: douta=16'hcd2d;
30605: douta=16'hccca;
30606: douta=16'hcca9;
30607: douta=16'hc425;
30608: douta=16'hc425;
30609: douta=16'hc404;
30610: douta=16'hcc07;
30611: douta=16'hcc27;
30612: douta=16'hcc26;
30613: douta=16'hcc67;
30614: douta=16'hcc67;
30615: douta=16'hcc67;
30616: douta=16'hcc67;
30617: douta=16'hcc67;
30618: douta=16'hcc67;
30619: douta=16'hcc67;
30620: douta=16'hcc67;
30621: douta=16'hcc68;
30622: douta=16'hcc68;
30623: douta=16'hcc68;
30624: douta=16'hd488;
30625: douta=16'hcc68;
30626: douta=16'hcc68;
30627: douta=16'hcc68;
30628: douta=16'hcc68;
30629: douta=16'hcc88;
30630: douta=16'hcc88;
30631: douta=16'hd488;
30632: douta=16'hcc88;
30633: douta=16'hcc88;
30634: douta=16'hd488;
30635: douta=16'hcc88;
30636: douta=16'hcc88;
30637: douta=16'hd488;
30638: douta=16'hcc88;
30639: douta=16'hcc88;
30640: douta=16'hcc88;
30641: douta=16'hd488;
30642: douta=16'hd4a9;
30643: douta=16'hd488;
30644: douta=16'hcc88;
30645: douta=16'hd488;
30646: douta=16'hcc88;
30647: douta=16'hd488;
30648: douta=16'hd488;
30649: douta=16'hd487;
30650: douta=16'had31;
30651: douta=16'he6d8;
30652: douta=16'hcc88;
30653: douta=16'hcc88;
30654: douta=16'hcc68;
30655: douta=16'hcc88;
30656: douta=16'hcc88;
30657: douta=16'hcc88;
30658: douta=16'hcc88;
30659: douta=16'hcc88;
30660: douta=16'hcc68;
30661: douta=16'h93ee;
30662: douta=16'h940e;
30663: douta=16'h940e;
30664: douta=16'hbd32;
30665: douta=16'hbd32;
30666: douta=16'hc573;
30667: douta=16'hbd33;
30668: douta=16'hc594;
30669: douta=16'hcdd5;
30670: douta=16'hc553;
30671: douta=16'hbd13;
30672: douta=16'hb4d3;
30673: douta=16'ha492;
30674: douta=16'h8412;
30675: douta=16'h8432;
30676: douta=16'h83f1;
30677: douta=16'h8412;
30678: douta=16'h7390;
30679: douta=16'h632e;
30680: douta=16'h7bb0;
30681: douta=16'h736f;
30682: douta=16'h6b2e;
30683: douta=16'h62ed;
30684: douta=16'h6b4e;
30685: douta=16'h7c12;
30686: douta=16'h6b6f;
30687: douta=16'h6b0d;
30688: douta=16'h526c;
30689: douta=16'h526b;
30690: douta=16'h52ab;
30691: douta=16'h6b2e;
30692: douta=16'h736f;
30693: douta=16'h8bf0;
30694: douta=16'h8c73;
30695: douta=16'h632f;
30696: douta=16'h528d;
30697: douta=16'h7bb1;
30698: douta=16'h630e;
30699: douta=16'h52ce;
30700: douta=16'h9d55;
30701: douta=16'hc67a;
30702: douta=16'hf7ff;
30703: douta=16'hffff;
30704: douta=16'hfefa;
30705: douta=16'hf636;
30706: douta=16'hbb47;
30707: douta=16'h9aa3;
30708: douta=16'h9b47;
30709: douta=16'ha388;
30710: douta=16'ha368;
30711: douta=16'ha368;
30712: douta=16'ha368;
30713: douta=16'ha368;
30714: douta=16'ha349;
30715: douta=16'ha348;
30716: douta=16'ha348;
30717: douta=16'h9b48;
30718: douta=16'ha348;
30719: douta=16'h9b48;
30720: douta=16'hcdb5;
30721: douta=16'had15;
30722: douta=16'h9473;
30723: douta=16'ha515;
30724: douta=16'ha4d5;
30725: douta=16'ha4f5;
30726: douta=16'h94d5;
30727: douta=16'h6370;
30728: douta=16'h39e8;
30729: douta=16'h3166;
30730: douta=16'h20a2;
30731: douta=16'h28e3;
30732: douta=16'h28e3;
30733: douta=16'h20e3;
30734: douta=16'h20e3;
30735: douta=16'h20e3;
30736: douta=16'h20e3;
30737: douta=16'h20c3;
30738: douta=16'h20a2;
30739: douta=16'h20a2;
30740: douta=16'h20a2;
30741: douta=16'h20c2;
30742: douta=16'h20a2;
30743: douta=16'h20a2;
30744: douta=16'h20a2;
30745: douta=16'h28e3;
30746: douta=16'h28e3;
30747: douta=16'h28e2;
30748: douta=16'h3103;
30749: douta=16'h3123;
30750: douta=16'h3923;
30751: douta=16'h3923;
30752: douta=16'h4143;
30753: douta=16'h49e8;
30754: douta=16'h10a5;
30755: douta=16'h3924;
30756: douta=16'h59a4;
30757: douta=16'h59c4;
30758: douta=16'h59c4;
30759: douta=16'h61c4;
30760: douta=16'h61c4;
30761: douta=16'h61c3;
30762: douta=16'h69c3;
30763: douta=16'h6a03;
30764: douta=16'h7223;
30765: douta=16'h7244;
30766: douta=16'h82e7;
30767: douta=16'h8b49;
30768: douta=16'h9beb;
30769: douta=16'hb4ce;
30770: douta=16'hb50f;
30771: douta=16'hc5b1;
30772: douta=16'hd633;
30773: douta=16'hd653;
30774: douta=16'he6f5;
30775: douta=16'hcdf2;
30776: douta=16'hc5b1;
30777: douta=16'hbd4f;
30778: douta=16'hb4ad;
30779: douta=16'ha40a;
30780: douta=16'ha3ca;
30781: douta=16'ha387;
30782: douta=16'ha386;
30783: douta=16'ha345;
30784: douta=16'hab65;
30785: douta=16'hab65;
30786: douta=16'hb385;
30787: douta=16'hb3a6;
30788: douta=16'hbbe6;
30789: douta=16'hbbe6;
30790: douta=16'hbbe7;
30791: douta=16'hbc07;
30792: douta=16'hc407;
30793: douta=16'hc426;
30794: douta=16'hc426;
30795: douta=16'hc428;
30796: douta=16'hc447;
30797: douta=16'hc447;
30798: douta=16'hc447;
30799: douta=16'hc447;
30800: douta=16'hc447;
30801: douta=16'hcc67;
30802: douta=16'hcc47;
30803: douta=16'hcc47;
30804: douta=16'hcc47;
30805: douta=16'hcc48;
30806: douta=16'hcc67;
30807: douta=16'hcc67;
30808: douta=16'hcc67;
30809: douta=16'hcc67;
30810: douta=16'hcc68;
30811: douta=16'hcc68;
30812: douta=16'hcc68;
30813: douta=16'hcc68;
30814: douta=16'hcc68;
30815: douta=16'hcc67;
30816: douta=16'hcc68;
30817: douta=16'hcc68;
30818: douta=16'hcc68;
30819: douta=16'hcc68;
30820: douta=16'hd488;
30821: douta=16'hcc68;
30822: douta=16'hcc88;
30823: douta=16'hcc88;
30824: douta=16'hcc88;
30825: douta=16'hcc68;
30826: douta=16'hcc88;
30827: douta=16'hd488;
30828: douta=16'hd489;
30829: douta=16'hcc88;
30830: douta=16'hd488;
30831: douta=16'hcc88;
30832: douta=16'hd489;
30833: douta=16'hd489;
30834: douta=16'hd488;
30835: douta=16'hd4a9;
30836: douta=16'hd4a9;
30837: douta=16'hd488;
30838: douta=16'hcc88;
30839: douta=16'hcc88;
30840: douta=16'hcc88;
30841: douta=16'hd487;
30842: douta=16'had32;
30843: douta=16'hdeb7;
30844: douta=16'hcc88;
30845: douta=16'hcc88;
30846: douta=16'hcc88;
30847: douta=16'hd489;
30848: douta=16'hcc89;
30849: douta=16'hcc88;
30850: douta=16'hcc88;
30851: douta=16'hcc88;
30852: douta=16'hcc69;
30853: douta=16'h9430;
30854: douta=16'h940f;
30855: douta=16'h9c50;
30856: douta=16'hb513;
30857: douta=16'hb533;
30858: douta=16'hacf3;
30859: douta=16'hb513;
30860: douta=16'hacd4;
30861: douta=16'h9c93;
30862: douta=16'h8c53;
30863: douta=16'h8412;
30864: douta=16'h8432;
30865: douta=16'h7bf2;
30866: douta=16'h8412;
30867: douta=16'h8433;
30868: douta=16'h630e;
30869: douta=16'h6b2e;
30870: douta=16'h62ed;
30871: douta=16'h630d;
30872: douta=16'h62cd;
30873: douta=16'h62ed;
30874: douta=16'h630e;
30875: douta=16'h62ed;
30876: douta=16'h62ed;
30877: douta=16'h7b8f;
30878: douta=16'h83d0;
30879: douta=16'h9c92;
30880: douta=16'ha493;
30881: douta=16'h838f;
30882: douta=16'h734e;
30883: douta=16'h83f0;
30884: douta=16'h6b4f;
30885: douta=16'h4a2a;
30886: douta=16'h8473;
30887: douta=16'hae18;
30888: douta=16'hc73d;
30889: douta=16'hffff;
30890: douta=16'hf636;
30891: douta=16'hd44d;
30892: douta=16'haac4;
30893: douta=16'h9ac4;
30894: douta=16'ha388;
30895: douta=16'ha388;
30896: douta=16'hab88;
30897: douta=16'ha388;
30898: douta=16'ha368;
30899: douta=16'hab88;
30900: douta=16'ha368;
30901: douta=16'ha368;
30902: douta=16'hab88;
30903: douta=16'hab68;
30904: douta=16'ha368;
30905: douta=16'ha368;
30906: douta=16'ha368;
30907: douta=16'ha368;
30908: douta=16'ha368;
30909: douta=16'ha368;
30910: douta=16'ha368;
30911: douta=16'ha369;
30912: douta=16'hc5b6;
30913: douta=16'h9494;
30914: douta=16'ha515;
30915: douta=16'ha4f5;
30916: douta=16'ha4f5;
30917: douta=16'ha4f5;
30918: douta=16'h8475;
30919: douta=16'h1020;
30920: douta=16'h3125;
30921: douta=16'h31a6;
30922: douta=16'h4aac;
30923: douta=16'h424b;
30924: douta=16'h3165;
30925: douta=16'h2082;
30926: douta=16'h28c3;
30927: douta=16'h20c3;
30928: douta=16'h20c3;
30929: douta=16'h20e3;
30930: douta=16'h1882;
30931: douta=16'h20a2;
30932: douta=16'h20a2;
30933: douta=16'h20c2;
30934: douta=16'h20a2;
30935: douta=16'h20a2;
30936: douta=16'h20c2;
30937: douta=16'h28e3;
30938: douta=16'h28e2;
30939: douta=16'h28e2;
30940: douta=16'h30e2;
30941: douta=16'h3103;
30942: douta=16'h30e2;
30943: douta=16'h3902;
30944: douta=16'h3902;
30945: douta=16'h4a4a;
30946: douta=16'h18c4;
30947: douta=16'h51c5;
30948: douta=16'h6246;
30949: douta=16'h7329;
30950: douta=16'h838b;
30951: douta=16'h8bcc;
30952: douta=16'hacef;
30953: douta=16'had30;
30954: douta=16'hbdb2;
30955: douta=16'hd675;
30956: douta=16'hbd71;
30957: douta=16'hbd51;
30958: douta=16'haccd;
30959: douta=16'ha44c;
30960: douta=16'h9bca;
30961: douta=16'h8b27;
30962: douta=16'h8b07;
30963: douta=16'h8ae6;
30964: douta=16'h8285;
30965: douta=16'h8285;
30966: douta=16'h8aa5;
30967: douta=16'h92e5;
30968: douta=16'h92c5;
30969: douta=16'h9306;
30970: douta=16'h9305;
30971: douta=16'h9306;
30972: douta=16'h9b27;
30973: douta=16'ha366;
30974: douta=16'hab86;
30975: douta=16'haba7;
30976: douta=16'hb3c7;
30977: douta=16'hb3c7;
30978: douta=16'hbbc7;
30979: douta=16'hbbe6;
30980: douta=16'hbbe7;
30981: douta=16'hc3e7;
30982: douta=16'hbc07;
30983: douta=16'hbc06;
30984: douta=16'hc427;
30985: douta=16'hc426;
30986: douta=16'hc447;
30987: douta=16'hc426;
30988: douta=16'hc447;
30989: douta=16'hc448;
30990: douta=16'hc448;
30991: douta=16'hcc47;
30992: douta=16'hcc47;
30993: douta=16'hcc47;
30994: douta=16'hcc67;
30995: douta=16'hcc67;
30996: douta=16'hcc47;
30997: douta=16'hcc68;
30998: douta=16'hcc48;
30999: douta=16'hcc68;
31000: douta=16'hcc48;
31001: douta=16'hcc48;
31002: douta=16'hcc68;
31003: douta=16'hcc68;
31004: douta=16'hcc68;
31005: douta=16'hcc68;
31006: douta=16'hcc68;
31007: douta=16'hcc68;
31008: douta=16'hcc68;
31009: douta=16'hcc68;
31010: douta=16'hcc68;
31011: douta=16'hcc68;
31012: douta=16'hcc68;
31013: douta=16'hcc68;
31014: douta=16'hd488;
31015: douta=16'hd488;
31016: douta=16'hd488;
31017: douta=16'hcc88;
31018: douta=16'hcc69;
31019: douta=16'hcc88;
31020: douta=16'hcc88;
31021: douta=16'hd4a9;
31022: douta=16'hd4a9;
31023: douta=16'hd488;
31024: douta=16'hd489;
31025: douta=16'hd489;
31026: douta=16'hd4a9;
31027: douta=16'hd4a9;
31028: douta=16'hd488;
31029: douta=16'hd488;
31030: douta=16'hd4a9;
31031: douta=16'hd4a9;
31032: douta=16'hd488;
31033: douta=16'hd488;
31034: douta=16'had32;
31035: douta=16'hdeb7;
31036: douta=16'hcc88;
31037: douta=16'hd488;
31038: douta=16'hcc88;
31039: douta=16'hcc89;
31040: douta=16'hcc89;
31041: douta=16'hcc88;
31042: douta=16'hcc89;
31043: douta=16'hcc69;
31044: douta=16'hcc89;
31045: douta=16'h9c0f;
31046: douta=16'h8bef;
31047: douta=16'h9c51;
31048: douta=16'h9452;
31049: douta=16'ha4d4;
31050: douta=16'ha4d4;
31051: douta=16'h9cb3;
31052: douta=16'h9452;
31053: douta=16'h8432;
31054: douta=16'h73b0;
31055: douta=16'h6b90;
31056: douta=16'h6b6f;
31057: douta=16'h6b70;
31058: douta=16'h630e;
31059: douta=16'h630e;
31060: douta=16'h630e;
31061: douta=16'h630e;
31062: douta=16'h62cd;
31063: douta=16'h62cd;
31064: douta=16'h62ed;
31065: douta=16'h6b0d;
31066: douta=16'h8c11;
31067: douta=16'h8bf1;
31068: douta=16'h9452;
31069: douta=16'h6b4e;
31070: douta=16'h7bb0;
31071: douta=16'h7bb0;
31072: douta=16'h6acd;
31073: douta=16'h6b0d;
31074: douta=16'h6b8f;
31075: douta=16'hefff;
31076: douta=16'hffff;
31077: douta=16'hffff;
31078: douta=16'hed71;
31079: douta=16'hbb87;
31080: douta=16'hb305;
31081: douta=16'ha367;
31082: douta=16'haba8;
31083: douta=16'haba8;
31084: douta=16'ha388;
31085: douta=16'haba8;
31086: douta=16'hab88;
31087: douta=16'hab88;
31088: douta=16'ha388;
31089: douta=16'ha388;
31090: douta=16'hab88;
31091: douta=16'hab88;
31092: douta=16'hab89;
31093: douta=16'hab89;
31094: douta=16'ha388;
31095: douta=16'haba8;
31096: douta=16'hab88;
31097: douta=16'ha368;
31098: douta=16'ha368;
31099: douta=16'ha368;
31100: douta=16'ha368;
31101: douta=16'ha368;
31102: douta=16'hab68;
31103: douta=16'ha368;
31104: douta=16'hc596;
31105: douta=16'h8c53;
31106: douta=16'had36;
31107: douta=16'ha4f5;
31108: douta=16'ha515;
31109: douta=16'ha4f5;
31110: douta=16'h8cd6;
31111: douta=16'h1861;
31112: douta=16'h20c2;
31113: douta=16'h28c3;
31114: douta=16'h39c8;
31115: douta=16'h426b;
31116: douta=16'h42cd;
31117: douta=16'h3187;
31118: douta=16'h2082;
31119: douta=16'h2082;
31120: douta=16'h20c3;
31121: douta=16'h20e3;
31122: douta=16'h2082;
31123: douta=16'h20a2;
31124: douta=16'h20a2;
31125: douta=16'h20a2;
31126: douta=16'h20a2;
31127: douta=16'h2082;
31128: douta=16'h20a2;
31129: douta=16'h20a1;
31130: douta=16'h20a1;
31131: douta=16'h28c2;
31132: douta=16'h3123;
31133: douta=16'h4165;
31134: douta=16'h41a5;
31135: douta=16'h5227;
31136: douta=16'h62a9;
31137: douta=16'h4a29;
31138: douta=16'h3146;
31139: douta=16'h942f;
31140: douta=16'h9c8f;
31141: douta=16'ha4f1;
31142: douta=16'ha4f0;
31143: douta=16'hacf0;
31144: douta=16'h9c8e;
31145: douta=16'h9c6d;
31146: douta=16'h940c;
31147: douta=16'hb510;
31148: douta=16'h7aa6;
31149: douta=16'h7aa6;
31150: douta=16'h7a64;
31151: douta=16'h7a44;
31152: douta=16'h7a44;
31153: douta=16'h7a64;
31154: douta=16'h8284;
31155: douta=16'h8aa5;
31156: douta=16'h8ac5;
31157: douta=16'h8ae6;
31158: douta=16'h92e6;
31159: douta=16'h9b27;
31160: douta=16'h9306;
31161: douta=16'h9326;
31162: douta=16'h9307;
31163: douta=16'h9306;
31164: douta=16'h9b26;
31165: douta=16'ha367;
31166: douta=16'hab86;
31167: douta=16'hab87;
31168: douta=16'hb3c7;
31169: douta=16'hb3c7;
31170: douta=16'hb3c6;
31171: douta=16'hbbe6;
31172: douta=16'hbbe7;
31173: douta=16'hbc07;
31174: douta=16'hc406;
31175: douta=16'hbc06;
31176: douta=16'hbc07;
31177: douta=16'hc407;
31178: douta=16'hc427;
31179: douta=16'hc427;
31180: douta=16'hc447;
31181: douta=16'hc427;
31182: douta=16'hc448;
31183: douta=16'hcc47;
31184: douta=16'hc447;
31185: douta=16'hc447;
31186: douta=16'hcc47;
31187: douta=16'hcc47;
31188: douta=16'hcc47;
31189: douta=16'hcc47;
31190: douta=16'hcc68;
31191: douta=16'hcc67;
31192: douta=16'hcc68;
31193: douta=16'hcc68;
31194: douta=16'hcc48;
31195: douta=16'hcc47;
31196: douta=16'hcc88;
31197: douta=16'hcc68;
31198: douta=16'hcc68;
31199: douta=16'hcc68;
31200: douta=16'hcc68;
31201: douta=16'hcc68;
31202: douta=16'hcc68;
31203: douta=16'hcc68;
31204: douta=16'hd488;
31205: douta=16'hcc68;
31206: douta=16'hcc88;
31207: douta=16'hcc68;
31208: douta=16'hcc68;
31209: douta=16'hcc88;
31210: douta=16'hd489;
31211: douta=16'hcc88;
31212: douta=16'hcc88;
31213: douta=16'hcc88;
31214: douta=16'hd488;
31215: douta=16'hcc88;
31216: douta=16'hd489;
31217: douta=16'hd489;
31218: douta=16'hd4a9;
31219: douta=16'hcc88;
31220: douta=16'hcc88;
31221: douta=16'hd4a9;
31222: douta=16'hd488;
31223: douta=16'hd488;
31224: douta=16'hcc88;
31225: douta=16'hd488;
31226: douta=16'had32;
31227: douta=16'hdeb8;
31228: douta=16'hcc88;
31229: douta=16'hcc89;
31230: douta=16'hcc88;
31231: douta=16'hcc89;
31232: douta=16'hcc89;
31233: douta=16'hcc88;
31234: douta=16'hcc89;
31235: douta=16'hcc69;
31236: douta=16'hcc69;
31237: douta=16'ha42d;
31238: douta=16'h83f0;
31239: douta=16'h9431;
31240: douta=16'h9c73;
31241: douta=16'h9452;
31242: douta=16'h8c73;
31243: douta=16'h8c53;
31244: douta=16'h7bf2;
31245: douta=16'h7bd1;
31246: douta=16'h6b6f;
31247: douta=16'h6b2e;
31248: douta=16'h6b4f;
31249: douta=16'h6b4f;
31250: douta=16'h6b4f;
31251: douta=16'h5acd;
31252: douta=16'h5aee;
31253: douta=16'h62ad;
31254: douta=16'h62cd;
31255: douta=16'h8c32;
31256: douta=16'h7bd0;
31257: douta=16'h8c11;
31258: douta=16'h9c72;
31259: douta=16'h422a;
31260: douta=16'h9432;
31261: douta=16'h62ad;
31262: douta=16'h5aad;
31263: douta=16'h73b0;
31264: douta=16'h8c93;
31265: douta=16'hc71c;
31266: douta=16'hefff;
31267: douta=16'hff1a;
31268: douta=16'hf5d4;
31269: douta=16'hcbca;
31270: douta=16'ha2e3;
31271: douta=16'ha3a7;
31272: douta=16'habc8;
31273: douta=16'haba8;
31274: douta=16'hb3a8;
31275: douta=16'hb3c8;
31276: douta=16'haba8;
31277: douta=16'hab88;
31278: douta=16'hab88;
31279: douta=16'hab89;
31280: douta=16'hab88;
31281: douta=16'hb3a8;
31282: douta=16'haba9;
31283: douta=16'hab89;
31284: douta=16'haba8;
31285: douta=16'hab88;
31286: douta=16'hab88;
31287: douta=16'hab88;
31288: douta=16'hab88;
31289: douta=16'hab88;
31290: douta=16'hab89;
31291: douta=16'ha368;
31292: douta=16'ha368;
31293: douta=16'ha368;
31294: douta=16'hab68;
31295: douta=16'ha368;
31296: douta=16'hb536;
31297: douta=16'h8c53;
31298: douta=16'ha4f5;
31299: douta=16'had36;
31300: douta=16'h9cf5;
31301: douta=16'h8c95;
31302: douta=16'h8cf7;
31303: douta=16'h28e3;
31304: douta=16'h2903;
31305: douta=16'h28e3;
31306: douta=16'h28e3;
31307: douta=16'h2903;
31308: douta=16'h20c3;
31309: douta=16'h20a2;
31310: douta=16'h2924;
31311: douta=16'h2966;
31312: douta=16'h4aac;
31313: douta=16'h31a8;
31314: douta=16'h39c8;
31315: douta=16'h39e8;
31316: douta=16'h3a08;
31317: douta=16'h39c7;
31318: douta=16'h39c7;
31319: douta=16'h39c7;
31320: douta=16'h39a6;
31321: douta=16'h41a6;
31322: douta=16'h39a5;
31323: douta=16'h3985;
31324: douta=16'h3944;
31325: douta=16'h3944;
31326: douta=16'h3943;
31327: douta=16'h3922;
31328: douta=16'h3923;
31329: douta=16'h4a4a;
31330: douta=16'h3944;
31331: douta=16'h59a3;
31332: douta=16'h59a4;
31333: douta=16'h61e4;
31334: douta=16'h59c4;
31335: douta=16'h61e4;
31336: douta=16'h6204;
31337: douta=16'h6a04;
31338: douta=16'h7265;
31339: douta=16'h82e7;
31340: douta=16'h7a84;
31341: douta=16'h7a85;
31342: douta=16'h7a85;
31343: douta=16'h82a5;
31344: douta=16'h82a5;
31345: douta=16'h8aa5;
31346: douta=16'h8aa5;
31347: douta=16'h8ac6;
31348: douta=16'h8ac6;
31349: douta=16'h8ae7;
31350: douta=16'h9307;
31351: douta=16'h9b47;
31352: douta=16'h9306;
31353: douta=16'h9306;
31354: douta=16'h9326;
31355: douta=16'h9326;
31356: douta=16'h9327;
31357: douta=16'ha367;
31358: douta=16'hab86;
31359: douta=16'haba7;
31360: douta=16'hb3c6;
31361: douta=16'hb3c7;
31362: douta=16'hbbe7;
31363: douta=16'hbbe7;
31364: douta=16'hbbe7;
31365: douta=16'hbc07;
31366: douta=16'hbc07;
31367: douta=16'hc407;
31368: douta=16'hc407;
31369: douta=16'hc447;
31370: douta=16'hc427;
31371: douta=16'hc427;
31372: douta=16'hc428;
31373: douta=16'hc448;
31374: douta=16'hc428;
31375: douta=16'hcc47;
31376: douta=16'hc447;
31377: douta=16'hcc47;
31378: douta=16'hcc67;
31379: douta=16'hcc68;
31380: douta=16'hcc67;
31381: douta=16'hcc47;
31382: douta=16'hcc68;
31383: douta=16'hcc48;
31384: douta=16'hcc68;
31385: douta=16'hcc68;
31386: douta=16'hcc68;
31387: douta=16'hcc68;
31388: douta=16'hcc68;
31389: douta=16'hcc68;
31390: douta=16'hcc68;
31391: douta=16'hcc68;
31392: douta=16'hcc68;
31393: douta=16'hcc68;
31394: douta=16'hcc68;
31395: douta=16'hcc68;
31396: douta=16'hcc88;
31397: douta=16'hcc88;
31398: douta=16'hcc88;
31399: douta=16'hcc88;
31400: douta=16'hcc88;
31401: douta=16'hcc89;
31402: douta=16'hd4aa;
31403: douta=16'hd489;
31404: douta=16'hd489;
31405: douta=16'hd488;
31406: douta=16'hcc88;
31407: douta=16'hcc89;
31408: douta=16'hd489;
31409: douta=16'hcc89;
31410: douta=16'hcc88;
31411: douta=16'hcc88;
31412: douta=16'hd488;
31413: douta=16'hcc89;
31414: douta=16'hd4a9;
31415: douta=16'hcc88;
31416: douta=16'hd489;
31417: douta=16'hd488;
31418: douta=16'had53;
31419: douta=16'hdeb7;
31420: douta=16'hcc89;
31421: douta=16'hcc89;
31422: douta=16'hcc89;
31423: douta=16'hcc89;
31424: douta=16'hcc69;
31425: douta=16'hd489;
31426: douta=16'hcc69;
31427: douta=16'hcc69;
31428: douta=16'hcc69;
31429: douta=16'hd486;
31430: douta=16'hb44d;
31431: douta=16'h9430;
31432: douta=16'h83d0;
31433: douta=16'h7bd1;
31434: douta=16'h83f1;
31435: douta=16'h73b0;
31436: douta=16'h7bb1;
31437: douta=16'h6b4f;
31438: douta=16'h630e;
31439: douta=16'h62cd;
31440: douta=16'h62ed;
31441: douta=16'h734e;
31442: douta=16'h8411;
31443: douta=16'h9472;
31444: douta=16'h83d0;
31445: douta=16'h7baf;
31446: douta=16'h5a8c;
31447: douta=16'h628c;
31448: douta=16'h630d;
31449: douta=16'h8431;
31450: douta=16'hdf5d;
31451: douta=16'hffff;
31452: douta=16'hffff;
31453: douta=16'hfeb9;
31454: douta=16'hedf4;
31455: douta=16'hcba8;
31456: douta=16'hb344;
31457: douta=16'hb3e8;
31458: douta=16'hb3e8;
31459: douta=16'hb3c8;
31460: douta=16'hb3c8;
31461: douta=16'hb3a8;
31462: douta=16'hb3a8;
31463: douta=16'hb3c8;
31464: douta=16'hb3c8;
31465: douta=16'hb3c8;
31466: douta=16'hb3c8;
31467: douta=16'hb3c8;
31468: douta=16'haba8;
31469: douta=16'haba8;
31470: douta=16'hb3c9;
31471: douta=16'hb3c8;
31472: douta=16'hb3a8;
31473: douta=16'hb3c8;
31474: douta=16'haba8;
31475: douta=16'hab88;
31476: douta=16'hab89;
31477: douta=16'hab88;
31478: douta=16'hab88;
31479: douta=16'hab89;
31480: douta=16'hab88;
31481: douta=16'hab89;
31482: douta=16'hab89;
31483: douta=16'ha368;
31484: douta=16'ha368;
31485: douta=16'ha368;
31486: douta=16'hab88;
31487: douta=16'hab68;
31488: douta=16'ha4f6;
31489: douta=16'ha4f5;
31490: douta=16'h9cb4;
31491: douta=16'had36;
31492: douta=16'h8cb6;
31493: douta=16'h8c96;
31494: douta=16'h634f;
31495: douta=16'h2903;
31496: douta=16'h28e3;
31497: douta=16'h28e3;
31498: douta=16'h28e3;
31499: douta=16'h28e3;
31500: douta=16'h28e3;
31501: douta=16'h28e3;
31502: douta=16'h20a3;
31503: douta=16'h20c3;
31504: douta=16'h20a3;
31505: douta=16'h20c3;
31506: douta=16'h20a2;
31507: douta=16'h20a2;
31508: douta=16'h2082;
31509: douta=16'h20a2;
31510: douta=16'h20a2;
31511: douta=16'h20c2;
31512: douta=16'h20a2;
31513: douta=16'h30e2;
31514: douta=16'h30e2;
31515: douta=16'h3103;
31516: douta=16'h3103;
31517: douta=16'h4143;
31518: douta=16'h3923;
31519: douta=16'h4143;
31520: douta=16'h49a6;
31521: douta=16'h39e8;
31522: douta=16'h4985;
31523: douta=16'h59c4;
31524: douta=16'h59c4;
31525: douta=16'h59e4;
31526: douta=16'h61e4;
31527: douta=16'h6204;
31528: douta=16'h6a24;
31529: douta=16'h6a04;
31530: douta=16'h6a87;
31531: douta=16'h7244;
31532: douta=16'h7a84;
31533: douta=16'h7a64;
31534: douta=16'h7a85;
31535: douta=16'h82a5;
31536: douta=16'h82a5;
31537: douta=16'h8aa5;
31538: douta=16'h8ac6;
31539: douta=16'h8ac6;
31540: douta=16'h8ae6;
31541: douta=16'h8ac6;
31542: douta=16'h8ac6;
31543: douta=16'h9b26;
31544: douta=16'h9306;
31545: douta=16'h9b47;
31546: douta=16'h9326;
31547: douta=16'h9326;
31548: douta=16'h9b27;
31549: douta=16'ha367;
31550: douta=16'ha386;
31551: douta=16'haba7;
31552: douta=16'hb3c6;
31553: douta=16'hb3c7;
31554: douta=16'hbbc7;
31555: douta=16'hbbe7;
31556: douta=16'hbbe7;
31557: douta=16'hbbe7;
31558: douta=16'hbc07;
31559: douta=16'hc407;
31560: douta=16'hc407;
31561: douta=16'hc427;
31562: douta=16'hc427;
31563: douta=16'hc427;
31564: douta=16'hc427;
31565: douta=16'hc428;
31566: douta=16'hc428;
31567: douta=16'hcc47;
31568: douta=16'hcc47;
31569: douta=16'hcc47;
31570: douta=16'hcc47;
31571: douta=16'hcc47;
31572: douta=16'hcc68;
31573: douta=16'hcc67;
31574: douta=16'hcc68;
31575: douta=16'hcc68;
31576: douta=16'hcc48;
31577: douta=16'hcc48;
31578: douta=16'hcc68;
31579: douta=16'hcc68;
31580: douta=16'hcc68;
31581: douta=16'hcc68;
31582: douta=16'hcc68;
31583: douta=16'hcc68;
31584: douta=16'hcc68;
31585: douta=16'hcc69;
31586: douta=16'hcc69;
31587: douta=16'hcc88;
31588: douta=16'hcc88;
31589: douta=16'hcc88;
31590: douta=16'hcc88;
31591: douta=16'hcc89;
31592: douta=16'hcc89;
31593: douta=16'hcc88;
31594: douta=16'hcc68;
31595: douta=16'hcc88;
31596: douta=16'hcc88;
31597: douta=16'hd488;
31598: douta=16'hd488;
31599: douta=16'hcc89;
31600: douta=16'hcc89;
31601: douta=16'hcc89;
31602: douta=16'hd488;
31603: douta=16'hd488;
31604: douta=16'hcc88;
31605: douta=16'hd489;
31606: douta=16'hcc89;
31607: douta=16'hcc89;
31608: douta=16'hcc89;
31609: douta=16'hd488;
31610: douta=16'had33;
31611: douta=16'hdeb7;
31612: douta=16'hcc89;
31613: douta=16'hcc89;
31614: douta=16'hcc69;
31615: douta=16'hcc89;
31616: douta=16'hcc89;
31617: douta=16'hcc69;
31618: douta=16'hcc69;
31619: douta=16'hcc68;
31620: douta=16'hcc49;
31621: douta=16'hcc69;
31622: douta=16'hdc86;
31623: douta=16'h7bf1;
31624: douta=16'h8411;
31625: douta=16'h7390;
31626: douta=16'h738f;
31627: douta=16'h6b4f;
31628: douta=16'h6b4f;
31629: douta=16'h5aed;
31630: douta=16'h422b;
31631: douta=16'h62ee;
31632: douta=16'h528d;
31633: douta=16'h7bb0;
31634: douta=16'h7b90;
31635: douta=16'h7b90;
31636: douta=16'h6b4f;
31637: douta=16'h8431;
31638: douta=16'hadd7;
31639: douta=16'hffff;
31640: douta=16'hffff;
31641: douta=16'hff9c;
31642: douta=16'hdd0e;
31643: douta=16'hcbc7;
31644: douta=16'hbb64;
31645: douta=16'hbc08;
31646: douta=16'hbc08;
31647: douta=16'hbc09;
31648: douta=16'hbbe9;
31649: douta=16'hb3c9;
31650: douta=16'hbbe9;
31651: douta=16'hb3c8;
31652: douta=16'hbbc9;
31653: douta=16'hb3e9;
31654: douta=16'hb3e9;
31655: douta=16'hb3c8;
31656: douta=16'hb3c8;
31657: douta=16'hb3c8;
31658: douta=16'hb3a8;
31659: douta=16'hb3c8;
31660: douta=16'hb3c8;
31661: douta=16'hb3a8;
31662: douta=16'hb3a8;
31663: douta=16'hb3c8;
31664: douta=16'hb3c8;
31665: douta=16'hb3a8;
31666: douta=16'hb3c8;
31667: douta=16'haba8;
31668: douta=16'hb3a8;
31669: douta=16'hab88;
31670: douta=16'hab88;
31671: douta=16'hab89;
31672: douta=16'hab88;
31673: douta=16'hab88;
31674: douta=16'hab89;
31675: douta=16'ha368;
31676: douta=16'hab88;
31677: douta=16'ha368;
31678: douta=16'hab68;
31679: douta=16'ha368;
31680: douta=16'h9cb5;
31681: douta=16'ha516;
31682: douta=16'ha4f4;
31683: douta=16'had16;
31684: douta=16'h8cb6;
31685: douta=16'h94d6;
31686: douta=16'h422a;
31687: douta=16'h2903;
31688: douta=16'h28e3;
31689: douta=16'h28e3;
31690: douta=16'h28e3;
31691: douta=16'h28e3;
31692: douta=16'h20e3;
31693: douta=16'h28e3;
31694: douta=16'h20c3;
31695: douta=16'h20c3;
31696: douta=16'h20c3;
31697: douta=16'h2082;
31698: douta=16'h20a2;
31699: douta=16'h20a3;
31700: douta=16'h20a3;
31701: douta=16'h20c2;
31702: douta=16'h20c2;
31703: douta=16'h20c2;
31704: douta=16'h20c2;
31705: douta=16'h30e3;
31706: douta=16'h3103;
31707: douta=16'h3103;
31708: douta=16'h3923;
31709: douta=16'h4124;
31710: douta=16'h4123;
31711: douta=16'h4163;
31712: douta=16'h49c7;
31713: douta=16'h31a8;
31714: douta=16'h51a5;
31715: douta=16'h59c4;
31716: douta=16'h59c4;
31717: douta=16'h61e4;
31718: douta=16'h61e4;
31719: douta=16'h6204;
31720: douta=16'h6a04;
31721: douta=16'h7224;
31722: douta=16'h72c9;
31723: douta=16'h7203;
31724: douta=16'h7a64;
31725: douta=16'h7a84;
31726: douta=16'h7a85;
31727: douta=16'h82c6;
31728: douta=16'h82a5;
31729: douta=16'h8aa5;
31730: douta=16'h8aa5;
31731: douta=16'h8aa5;
31732: douta=16'h8ae6;
31733: douta=16'h8ac6;
31734: douta=16'h8ae6;
31735: douta=16'h9b26;
31736: douta=16'h9326;
31737: douta=16'h9b47;
31738: douta=16'h9306;
31739: douta=16'h9326;
31740: douta=16'h9327;
31741: douta=16'ha367;
31742: douta=16'hab87;
31743: douta=16'hab87;
31744: douta=16'hb3c6;
31745: douta=16'hb3c7;
31746: douta=16'hbbe8;
31747: douta=16'hbbe7;
31748: douta=16'hbbe7;
31749: douta=16'hbbe7;
31750: douta=16'hbbe7;
31751: douta=16'hc407;
31752: douta=16'hc427;
31753: douta=16'hc427;
31754: douta=16'hc428;
31755: douta=16'hc427;
31756: douta=16'hc427;
31757: douta=16'hc428;
31758: douta=16'hc428;
31759: douta=16'hcc47;
31760: douta=16'hcc47;
31761: douta=16'hcc47;
31762: douta=16'hcc47;
31763: douta=16'hcc67;
31764: douta=16'hcc67;
31765: douta=16'hcc68;
31766: douta=16'hcc67;
31767: douta=16'hcc67;
31768: douta=16'hcc68;
31769: douta=16'hcc48;
31770: douta=16'hcc68;
31771: douta=16'hcc68;
31772: douta=16'hcc68;
31773: douta=16'hcc68;
31774: douta=16'hcc48;
31775: douta=16'hcc68;
31776: douta=16'hcc68;
31777: douta=16'hcc69;
31778: douta=16'hcc69;
31779: douta=16'hcc89;
31780: douta=16'hcc88;
31781: douta=16'hcc88;
31782: douta=16'hcc88;
31783: douta=16'hcc89;
31784: douta=16'hcc89;
31785: douta=16'hcc89;
31786: douta=16'hcc89;
31787: douta=16'hd489;
31788: douta=16'hcc89;
31789: douta=16'hd489;
31790: douta=16'hd489;
31791: douta=16'hcc89;
31792: douta=16'hcc89;
31793: douta=16'hd489;
31794: douta=16'hd488;
31795: douta=16'hcc89;
31796: douta=16'hd489;
31797: douta=16'hd489;
31798: douta=16'hcc89;
31799: douta=16'hcc69;
31800: douta=16'hcc89;
31801: douta=16'hd488;
31802: douta=16'had53;
31803: douta=16'he6b7;
31804: douta=16'hcc89;
31805: douta=16'hcc89;
31806: douta=16'hcc69;
31807: douta=16'hcc89;
31808: douta=16'hcc89;
31809: douta=16'hcc89;
31810: douta=16'hcc89;
31811: douta=16'hcc89;
31812: douta=16'hcc69;
31813: douta=16'hcc69;
31814: douta=16'hd487;
31815: douta=16'h7bd0;
31816: douta=16'h83f0;
31817: douta=16'h7390;
31818: douta=16'h6b6e;
31819: douta=16'h6b2e;
31820: douta=16'h528c;
31821: douta=16'h528c;
31822: douta=16'h83f1;
31823: douta=16'h9473;
31824: douta=16'h31cb;
31825: douta=16'h62ed;
31826: douta=16'h62cd;
31827: douta=16'h630e;
31828: douta=16'hc69b;
31829: douta=16'hef9f;
31830: douta=16'hffff;
31831: douta=16'he615;
31832: douta=16'hd48c;
31833: douta=16'hcc09;
31834: douta=16'hbb85;
31835: douta=16'hbc28;
31836: douta=16'hc429;
31837: douta=16'hbc09;
31838: douta=16'hbc08;
31839: douta=16'hbbe8;
31840: douta=16'hbc09;
31841: douta=16'hbbe9;
31842: douta=16'hbbe9;
31843: douta=16'hbbe9;
31844: douta=16'hb3e9;
31845: douta=16'hb3e8;
31846: douta=16'hbbe9;
31847: douta=16'hb3e9;
31848: douta=16'hb3c9;
31849: douta=16'hb3c8;
31850: douta=16'hb3e9;
31851: douta=16'hb3a8;
31852: douta=16'hb3c8;
31853: douta=16'hb3a8;
31854: douta=16'hb3a8;
31855: douta=16'hb3a9;
31856: douta=16'hb3c9;
31857: douta=16'hb3c8;
31858: douta=16'hb3c8;
31859: douta=16'haba8;
31860: douta=16'hab88;
31861: douta=16'hab88;
31862: douta=16'haba9;
31863: douta=16'hab89;
31864: douta=16'hab88;
31865: douta=16'hab88;
31866: douta=16'hab88;
31867: douta=16'hab88;
31868: douta=16'ha368;
31869: douta=16'hab68;
31870: douta=16'ha368;
31871: douta=16'ha368;
31872: douta=16'h9c94;
31873: douta=16'ha516;
31874: douta=16'hb555;
31875: douta=16'ha516;
31876: douta=16'h94f6;
31877: douta=16'h9518;
31878: douta=16'h1861;
31879: douta=16'h28e3;
31880: douta=16'h28e3;
31881: douta=16'h28e3;
31882: douta=16'h20c2;
31883: douta=16'h28e3;
31884: douta=16'h28e3;
31885: douta=16'h28e3;
31886: douta=16'h20c3;
31887: douta=16'h20c3;
31888: douta=16'h20e3;
31889: douta=16'h20a2;
31890: douta=16'h20c2;
31891: douta=16'h20a2;
31892: douta=16'h20c2;
31893: douta=16'h20c2;
31894: douta=16'h28c3;
31895: douta=16'h28e2;
31896: douta=16'h28c2;
31897: douta=16'h3103;
31898: douta=16'h3103;
31899: douta=16'h3103;
31900: douta=16'h3923;
31901: douta=16'h4143;
31902: douta=16'h4144;
31903: douta=16'h4964;
31904: douta=16'h4a49;
31905: douta=16'h1906;
31906: douta=16'h61c4;
31907: douta=16'h59c4;
31908: douta=16'h59c4;
31909: douta=16'h61e4;
31910: douta=16'h6204;
31911: douta=16'h6a04;
31912: douta=16'h7224;
31913: douta=16'h69e4;
31914: douta=16'h7bad;
31915: douta=16'h7a04;
31916: douta=16'h7a84;
31917: douta=16'h7a64;
31918: douta=16'h7a85;
31919: douta=16'h82a5;
31920: douta=16'h8aa5;
31921: douta=16'h8ac6;
31922: douta=16'h8aa5;
31923: douta=16'h8aa5;
31924: douta=16'h8ac6;
31925: douta=16'h8ae6;
31926: douta=16'h9307;
31927: douta=16'h9b47;
31928: douta=16'h9327;
31929: douta=16'h9b26;
31930: douta=16'h92e6;
31931: douta=16'h9327;
31932: douta=16'h9326;
31933: douta=16'hab87;
31934: douta=16'hab86;
31935: douta=16'haba7;
31936: douta=16'hb3e7;
31937: douta=16'hb3e6;
31938: douta=16'hb3e6;
31939: douta=16'hbbe7;
31940: douta=16'hbc07;
31941: douta=16'hbbe7;
31942: douta=16'hbc07;
31943: douta=16'hbc07;
31944: douta=16'hc407;
31945: douta=16'hc428;
31946: douta=16'hc427;
31947: douta=16'hc428;
31948: douta=16'hc448;
31949: douta=16'hc448;
31950: douta=16'hc448;
31951: douta=16'hcc47;
31952: douta=16'hcc47;
31953: douta=16'hc448;
31954: douta=16'hcc48;
31955: douta=16'hcc67;
31956: douta=16'hcc68;
31957: douta=16'hcc68;
31958: douta=16'hcc47;
31959: douta=16'hcc68;
31960: douta=16'hcc68;
31961: douta=16'hcc68;
31962: douta=16'hcc88;
31963: douta=16'hcc68;
31964: douta=16'hcc68;
31965: douta=16'hcc48;
31966: douta=16'hcc68;
31967: douta=16'hcc69;
31968: douta=16'hcc69;
31969: douta=16'hcc68;
31970: douta=16'hcc68;
31971: douta=16'hcc68;
31972: douta=16'hcc68;
31973: douta=16'hcc88;
31974: douta=16'hcc89;
31975: douta=16'hcc89;
31976: douta=16'hcc89;
31977: douta=16'hcc89;
31978: douta=16'hcc69;
31979: douta=16'hd489;
31980: douta=16'hcc89;
31981: douta=16'hd489;
31982: douta=16'hcc89;
31983: douta=16'hd489;
31984: douta=16'hd489;
31985: douta=16'hd489;
31986: douta=16'hd489;
31987: douta=16'hcc89;
31988: douta=16'hd489;
31989: douta=16'hd489;
31990: douta=16'hd4a9;
31991: douta=16'hcc89;
31992: douta=16'hcc88;
31993: douta=16'hd468;
31994: douta=16'had53;
31995: douta=16'he6b7;
31996: douta=16'hcc69;
31997: douta=16'hcc89;
31998: douta=16'hcc69;
31999: douta=16'hcc89;
32000: douta=16'hcc89;
32001: douta=16'hcc69;
32002: douta=16'hcc89;
32003: douta=16'hcc69;
32004: douta=16'hcc69;
32005: douta=16'hcc68;
32006: douta=16'hcc69;
32007: douta=16'hd487;
32008: douta=16'h7bf1;
32009: douta=16'h630e;
32010: douta=16'h8c74;
32011: douta=16'h94f6;
32012: douta=16'h7bd3;
32013: douta=16'h7bf1;
32014: douta=16'hdf7f;
32015: douta=16'he7ff;
32016: douta=16'hdfff;
32017: douta=16'hce18;
32018: douta=16'hc48e;
32019: douta=16'hc40a;
32020: douta=16'hc407;
32021: douta=16'hcc28;
32022: douta=16'hc449;
32023: douta=16'hc428;
32024: douta=16'hc429;
32025: douta=16'hc429;
32026: douta=16'hc429;
32027: douta=16'hc429;
32028: douta=16'hbc08;
32029: douta=16'hc429;
32030: douta=16'hbc09;
32031: douta=16'hbc09;
32032: douta=16'hbc09;
32033: douta=16'hbc09;
32034: douta=16'hbc09;
32035: douta=16'hbbe9;
32036: douta=16'hbc09;
32037: douta=16'hbbe9;
32038: douta=16'hbbe9;
32039: douta=16'hb3e8;
32040: douta=16'hb3e8;
32041: douta=16'hb3e8;
32042: douta=16'hb3e8;
32043: douta=16'hb3c8;
32044: douta=16'hb3a8;
32045: douta=16'hb3a8;
32046: douta=16'hb3c8;
32047: douta=16'hb3a9;
32048: douta=16'hb3a9;
32049: douta=16'hb3a8;
32050: douta=16'hb3c8;
32051: douta=16'haba8;
32052: douta=16'hb3a8;
32053: douta=16'haba9;
32054: douta=16'hab88;
32055: douta=16'hab89;
32056: douta=16'hab89;
32057: douta=16'hab88;
32058: douta=16'hab89;
32059: douta=16'hab89;
32060: douta=16'hab88;
32061: douta=16'ha389;
32062: douta=16'ha388;
32063: douta=16'ha388;
32064: douta=16'ha4f5;
32065: douta=16'h9cb4;
32066: douta=16'hbd75;
32067: douta=16'h94b5;
32068: douta=16'h8cb7;
32069: douta=16'h7c53;
32070: douta=16'h28e2;
32071: douta=16'h28e3;
32072: douta=16'h28e3;
32073: douta=16'h28e3;
32074: douta=16'h28e3;
32075: douta=16'h28e3;
32076: douta=16'h28e3;
32077: douta=16'h20c3;
32078: douta=16'h20c3;
32079: douta=16'h20a3;
32080: douta=16'h20c3;
32081: douta=16'h20a2;
32082: douta=16'h20a2;
32083: douta=16'h20c2;
32084: douta=16'h20c2;
32085: douta=16'h20c2;
32086: douta=16'h28e3;
32087: douta=16'h28e3;
32088: douta=16'h30e3;
32089: douta=16'h30e2;
32090: douta=16'h3103;
32091: douta=16'h3103;
32092: douta=16'h3923;
32093: douta=16'h4144;
32094: douta=16'h4143;
32095: douta=16'h4143;
32096: douta=16'h528b;
32097: douta=16'h10c5;
32098: douta=16'h59c4;
32099: douta=16'h59c4;
32100: douta=16'h59c4;
32101: douta=16'h61e4;
32102: douta=16'h6204;
32103: douta=16'h6a04;
32104: douta=16'h6a24;
32105: douta=16'h7203;
32106: douta=16'h9cb0;
32107: douta=16'h7a44;
32108: douta=16'h7a84;
32109: douta=16'h7a85;
32110: douta=16'h7a85;
32111: douta=16'h8aa6;
32112: douta=16'h8aa5;
32113: douta=16'h8ac6;
32114: douta=16'h8ac6;
32115: douta=16'h8ac6;
32116: douta=16'h8ac6;
32117: douta=16'h9307;
32118: douta=16'h9306;
32119: douta=16'h9b26;
32120: douta=16'h9b47;
32121: douta=16'h9b27;
32122: douta=16'h92e5;
32123: douta=16'h9326;
32124: douta=16'h9327;
32125: douta=16'hab87;
32126: douta=16'hab86;
32127: douta=16'hb3a7;
32128: douta=16'hb3c6;
32129: douta=16'hb3c7;
32130: douta=16'hb3c7;
32131: douta=16'hbbe7;
32132: douta=16'hbbe7;
32133: douta=16'hbc07;
32134: douta=16'hc407;
32135: douta=16'hbc07;
32136: douta=16'hc407;
32137: douta=16'hc428;
32138: douta=16'hc427;
32139: douta=16'hc428;
32140: douta=16'hc428;
32141: douta=16'hc448;
32142: douta=16'hc448;
32143: douta=16'hcc47;
32144: douta=16'hc447;
32145: douta=16'hcc67;
32146: douta=16'hcc48;
32147: douta=16'hcc67;
32148: douta=16'hcc47;
32149: douta=16'hcc67;
32150: douta=16'hcc68;
32151: douta=16'hcc47;
32152: douta=16'hcc67;
32153: douta=16'hcc68;
32154: douta=16'hcc68;
32155: douta=16'hcc68;
32156: douta=16'hcc68;
32157: douta=16'hcc68;
32158: douta=16'hcc68;
32159: douta=16'hcc68;
32160: douta=16'hcc68;
32161: douta=16'hcc88;
32162: douta=16'hcc68;
32163: douta=16'hcc68;
32164: douta=16'hcc69;
32165: douta=16'hd489;
32166: douta=16'hcc89;
32167: douta=16'hcc89;
32168: douta=16'hd489;
32169: douta=16'hd489;
32170: douta=16'hcc89;
32171: douta=16'hd48a;
32172: douta=16'hd489;
32173: douta=16'hcc89;
32174: douta=16'hd489;
32175: douta=16'hd489;
32176: douta=16'hcc89;
32177: douta=16'hcc69;
32178: douta=16'hcc89;
32179: douta=16'hcc8a;
32180: douta=16'hcc89;
32181: douta=16'hd489;
32182: douta=16'hcc89;
32183: douta=16'hcc89;
32184: douta=16'hd489;
32185: douta=16'hd468;
32186: douta=16'had33;
32187: douta=16'he6b7;
32188: douta=16'hcc69;
32189: douta=16'hcc89;
32190: douta=16'hcc69;
32191: douta=16'hcc69;
32192: douta=16'hcc69;
32193: douta=16'hcc89;
32194: douta=16'hcc69;
32195: douta=16'hcc69;
32196: douta=16'hcc69;
32197: douta=16'hcc69;
32198: douta=16'hcc69;
32199: douta=16'hc468;
32200: douta=16'hd447;
32201: douta=16'hc449;
32202: douta=16'hcc48;
32203: douta=16'hd468;
32204: douta=16'hd485;
32205: douta=16'hcc6b;
32206: douta=16'hbc4b;
32207: douta=16'hc428;
32208: douta=16'hc3a3;
32209: douta=16'hcc49;
32210: douta=16'hcc4a;
32211: douta=16'hc449;
32212: douta=16'hc449;
32213: douta=16'hc448;
32214: douta=16'hc428;
32215: douta=16'hc428;
32216: douta=16'hc449;
32217: douta=16'hc449;
32218: douta=16'hc429;
32219: douta=16'hbc08;
32220: douta=16'hc429;
32221: douta=16'hc429;
32222: douta=16'hbc09;
32223: douta=16'hbc09;
32224: douta=16'hbc09;
32225: douta=16'hbc09;
32226: douta=16'hbc09;
32227: douta=16'hbc09;
32228: douta=16'hbbe9;
32229: douta=16'hbbe9;
32230: douta=16'hbbe9;
32231: douta=16'hb3e9;
32232: douta=16'hb3e9;
32233: douta=16'hb3c9;
32234: douta=16'hb3c8;
32235: douta=16'hb3c9;
32236: douta=16'hb3c9;
32237: douta=16'hb3c8;
32238: douta=16'hb3a8;
32239: douta=16'hb3a8;
32240: douta=16'hb3c8;
32241: douta=16'hb3c9;
32242: douta=16'hb3c8;
32243: douta=16'hb3a8;
32244: douta=16'hb3a8;
32245: douta=16'hab89;
32246: douta=16'haba9;
32247: douta=16'hab89;
32248: douta=16'haba9;
32249: douta=16'haba8;
32250: douta=16'haba8;
32251: douta=16'haba8;
32252: douta=16'ha388;
32253: douta=16'ha388;
32254: douta=16'ha388;
32255: douta=16'ha389;
32256: douta=16'ha4d5;
32257: douta=16'h9cd4;
32258: douta=16'hb555;
32259: douta=16'h8c95;
32260: douta=16'h94f7;
32261: douta=16'h636f;
32262: douta=16'h28e3;
32263: douta=16'h28e3;
32264: douta=16'h28e3;
32265: douta=16'h28e3;
32266: douta=16'h28e3;
32267: douta=16'h28e3;
32268: douta=16'h28e3;
32269: douta=16'h20c3;
32270: douta=16'h20c3;
32271: douta=16'h20a3;
32272: douta=16'h20c3;
32273: douta=16'h20a2;
32274: douta=16'h20c2;
32275: douta=16'h20c2;
32276: douta=16'h20c2;
32277: douta=16'h28c3;
32278: douta=16'h28e2;
32279: douta=16'h28e3;
32280: douta=16'h30e3;
32281: douta=16'h3103;
32282: douta=16'h3103;
32283: douta=16'h3123;
32284: douta=16'h3944;
32285: douta=16'h4124;
32286: douta=16'h4164;
32287: douta=16'h4964;
32288: douta=16'h528b;
32289: douta=16'h10c5;
32290: douta=16'h59c4;
32291: douta=16'h59c4;
32292: douta=16'h61c4;
32293: douta=16'h61e4;
32294: douta=16'h6204;
32295: douta=16'h6a24;
32296: douta=16'h7224;
32297: douta=16'h6a03;
32298: douta=16'ha511;
32299: douta=16'h7a64;
32300: douta=16'h7a84;
32301: douta=16'h7a85;
32302: douta=16'h82a5;
32303: douta=16'h8aa6;
32304: douta=16'h8aa5;
32305: douta=16'h8ac6;
32306: douta=16'h8ac5;
32307: douta=16'h8ac6;
32308: douta=16'h8ac6;
32309: douta=16'h9306;
32310: douta=16'h9306;
32311: douta=16'h9306;
32312: douta=16'h9b46;
32313: douta=16'h9326;
32314: douta=16'h9306;
32315: douta=16'h9307;
32316: douta=16'h9326;
32317: douta=16'hab87;
32318: douta=16'haba7;
32319: douta=16'haba7;
32320: douta=16'hb3c6;
32321: douta=16'hb3c7;
32322: douta=16'hb3e6;
32323: douta=16'hbbe7;
32324: douta=16'hbc07;
32325: douta=16'hbbe7;
32326: douta=16'hbc07;
32327: douta=16'hbc07;
32328: douta=16'hbc07;
32329: douta=16'hc448;
32330: douta=16'hc427;
32331: douta=16'hc428;
32332: douta=16'hc448;
32333: douta=16'hc448;
32334: douta=16'hc428;
32335: douta=16'hc447;
32336: douta=16'hcc47;
32337: douta=16'hcc48;
32338: douta=16'hcc48;
32339: douta=16'hcc68;
32340: douta=16'hcc67;
32341: douta=16'hcc47;
32342: douta=16'hcc67;
32343: douta=16'hcc68;
32344: douta=16'hcc68;
32345: douta=16'hcc68;
32346: douta=16'hcc68;
32347: douta=16'hcc68;
32348: douta=16'hcc68;
32349: douta=16'hcc68;
32350: douta=16'hcc88;
32351: douta=16'hcc88;
32352: douta=16'hcc68;
32353: douta=16'hcc68;
32354: douta=16'hcc88;
32355: douta=16'hcc88;
32356: douta=16'hcc68;
32357: douta=16'hcc89;
32358: douta=16'hcc89;
32359: douta=16'hcc89;
32360: douta=16'hd489;
32361: douta=16'hcc89;
32362: douta=16'hcc89;
32363: douta=16'hd489;
32364: douta=16'hcc69;
32365: douta=16'hcc89;
32366: douta=16'hcc69;
32367: douta=16'hcc89;
32368: douta=16'hcc89;
32369: douta=16'hcc89;
32370: douta=16'hcc89;
32371: douta=16'hcc8a;
32372: douta=16'hcc69;
32373: douta=16'hd489;
32374: douta=16'hcc89;
32375: douta=16'hcc89;
32376: douta=16'hcc88;
32377: douta=16'hd468;
32378: douta=16'had53;
32379: douta=16'hde96;
32380: douta=16'hcc68;
32381: douta=16'hcc69;
32382: douta=16'hcc69;
32383: douta=16'hcc69;
32384: douta=16'hcc69;
32385: douta=16'hcc69;
32386: douta=16'hcc69;
32387: douta=16'hcc89;
32388: douta=16'hcc69;
32389: douta=16'hcc69;
32390: douta=16'hcc69;
32391: douta=16'hcc69;
32392: douta=16'hcc69;
32393: douta=16'hcc48;
32394: douta=16'hcc69;
32395: douta=16'hcc69;
32396: douta=16'hcc49;
32397: douta=16'hcc68;
32398: douta=16'hd447;
32399: douta=16'hcc68;
32400: douta=16'hcc49;
32401: douta=16'hc449;
32402: douta=16'hc448;
32403: douta=16'hc448;
32404: douta=16'hcc29;
32405: douta=16'hc448;
32406: douta=16'hc428;
32407: douta=16'hc428;
32408: douta=16'hc429;
32409: douta=16'hc429;
32410: douta=16'hc429;
32411: douta=16'hbc08;
32412: douta=16'hc429;
32413: douta=16'hc429;
32414: douta=16'hbc09;
32415: douta=16'hbc08;
32416: douta=16'hbc09;
32417: douta=16'hbc09;
32418: douta=16'hbc09;
32419: douta=16'hbbe9;
32420: douta=16'hbbe9;
32421: douta=16'hb3c9;
32422: douta=16'hb3e8;
32423: douta=16'hb3e9;
32424: douta=16'hb3e9;
32425: douta=16'hb3e9;
32426: douta=16'hb3c9;
32427: douta=16'hb3c8;
32428: douta=16'hb3c8;
32429: douta=16'hb3c8;
32430: douta=16'hb3a8;
32431: douta=16'hb3a8;
32432: douta=16'hb3a8;
32433: douta=16'hb3c8;
32434: douta=16'haba9;
32435: douta=16'hb3a8;
32436: douta=16'hb3c8;
32437: douta=16'haba9;
32438: douta=16'haba9;
32439: douta=16'haba9;
32440: douta=16'haba9;
32441: douta=16'haba8;
32442: douta=16'haba8;
32443: douta=16'ha388;
32444: douta=16'ha388;
32445: douta=16'ha388;
32446: douta=16'ha368;
32447: douta=16'ha368;
32448: douta=16'ha4f5;
32449: douta=16'ha4d4;
32450: douta=16'h9cf5;
32451: douta=16'h94d6;
32452: douta=16'h73b1;
32453: douta=16'h1881;
32454: douta=16'h2903;
32455: douta=16'h28e3;
32456: douta=16'h28e3;
32457: douta=16'h28e3;
32458: douta=16'h28e3;
32459: douta=16'h20c3;
32460: douta=16'h20c3;
32461: douta=16'h20c3;
32462: douta=16'h20c3;
32463: douta=16'h20c3;
32464: douta=16'h20a2;
32465: douta=16'h20a2;
32466: douta=16'h20c2;
32467: douta=16'h20a2;
32468: douta=16'h20a2;
32469: douta=16'h28c3;
32470: douta=16'h28e3;
32471: douta=16'h3103;
32472: douta=16'h3103;
32473: douta=16'h3103;
32474: douta=16'h3103;
32475: douta=16'h3923;
32476: douta=16'h4144;
32477: douta=16'h4163;
32478: douta=16'h4964;
32479: douta=16'h4985;
32480: douta=16'h4209;
32481: douta=16'h10c5;
32482: douta=16'h59a4;
32483: douta=16'h59c4;
32484: douta=16'h61e4;
32485: douta=16'h6204;
32486: douta=16'h6a04;
32487: douta=16'h6a04;
32488: douta=16'h6a24;
32489: douta=16'h7246;
32490: douta=16'hb572;
32491: douta=16'h7a64;
32492: douta=16'h7a85;
32493: douta=16'h7a85;
32494: douta=16'h82a5;
32495: douta=16'h82a6;
32496: douta=16'h8ac6;
32497: douta=16'h8ac6;
32498: douta=16'h8ac6;
32499: douta=16'h8ac6;
32500: douta=16'h8ac6;
32501: douta=16'h9306;
32502: douta=16'h9306;
32503: douta=16'h7266;
32504: douta=16'ha367;
32505: douta=16'h9326;
32506: douta=16'h9305;
32507: douta=16'h9305;
32508: douta=16'h9305;
32509: douta=16'ha366;
32510: douta=16'haba7;
32511: douta=16'hab87;
32512: douta=16'hb3c7;
32513: douta=16'hb3c7;
32514: douta=16'hbbe7;
32515: douta=16'hbbe7;
32516: douta=16'hbc07;
32517: douta=16'hbbe7;
32518: douta=16'hbc07;
32519: douta=16'hbc07;
32520: douta=16'hc428;
32521: douta=16'hc427;
32522: douta=16'hc427;
32523: douta=16'hc427;
32524: douta=16'hc427;
32525: douta=16'hc448;
32526: douta=16'hc448;
32527: douta=16'hcc47;
32528: douta=16'hc447;
32529: douta=16'hcc48;
32530: douta=16'hcc67;
32531: douta=16'hcc68;
32532: douta=16'hcc48;
32533: douta=16'hcc67;
32534: douta=16'hcc47;
32535: douta=16'hcc67;
32536: douta=16'hcc68;
32537: douta=16'hcc68;
32538: douta=16'hcc68;
32539: douta=16'hcc68;
32540: douta=16'hcc68;
32541: douta=16'hcc68;
32542: douta=16'hcc88;
32543: douta=16'hcc88;
32544: douta=16'hcc68;
32545: douta=16'hcc88;
32546: douta=16'hcc69;
32547: douta=16'hcc68;
32548: douta=16'hcc89;
32549: douta=16'hcc69;
32550: douta=16'hcc69;
32551: douta=16'hcc89;
32552: douta=16'hcc69;
32553: douta=16'hd489;
32554: douta=16'hcc69;
32555: douta=16'hd489;
32556: douta=16'hcc69;
32557: douta=16'hd48a;
32558: douta=16'hcc89;
32559: douta=16'hcc89;
32560: douta=16'hcc89;
32561: douta=16'hcc69;
32562: douta=16'hcc69;
32563: douta=16'hcc8a;
32564: douta=16'hcc89;
32565: douta=16'hcc8a;
32566: douta=16'hcc89;
32567: douta=16'hcc69;
32568: douta=16'hcc69;
32569: douta=16'hd468;
32570: douta=16'had73;
32571: douta=16'he696;
32572: douta=16'hcc69;
32573: douta=16'hcc69;
32574: douta=16'hcc69;
32575: douta=16'hcc89;
32576: douta=16'hcc69;
32577: douta=16'hcc69;
32578: douta=16'hcc69;
32579: douta=16'hcc69;
32580: douta=16'hcc69;
32581: douta=16'hcc69;
32582: douta=16'hcc69;
32583: douta=16'hcc69;
32584: douta=16'hcc68;
32585: douta=16'hcc6a;
32586: douta=16'hcc69;
32587: douta=16'hcc49;
32588: douta=16'hcc69;
32589: douta=16'hc468;
32590: douta=16'hc449;
32591: douta=16'hcc69;
32592: douta=16'hcc49;
32593: douta=16'hcc49;
32594: douta=16'hc449;
32595: douta=16'hc449;
32596: douta=16'hc449;
32597: douta=16'hc428;
32598: douta=16'hc428;
32599: douta=16'hc429;
32600: douta=16'hc429;
32601: douta=16'hc429;
32602: douta=16'hc429;
32603: douta=16'hc429;
32604: douta=16'hbc09;
32605: douta=16'hc429;
32606: douta=16'hc429;
32607: douta=16'hbc08;
32608: douta=16'hbc09;
32609: douta=16'hbc29;
32610: douta=16'hbc09;
32611: douta=16'hbbe9;
32612: douta=16'hbc09;
32613: douta=16'hbbe9;
32614: douta=16'hb3e8;
32615: douta=16'hbc09;
32616: douta=16'hb3e9;
32617: douta=16'hb3e9;
32618: douta=16'hb3e9;
32619: douta=16'hb3c8;
32620: douta=16'hb3c8;
32621: douta=16'hb3c9;
32622: douta=16'hb3c8;
32623: douta=16'hb3c8;
32624: douta=16'hb3c9;
32625: douta=16'hb3c8;
32626: douta=16'hb3c9;
32627: douta=16'haba9;
32628: douta=16'haba9;
32629: douta=16'haba9;
32630: douta=16'haba9;
32631: douta=16'haba9;
32632: douta=16'haba9;
32633: douta=16'haba9;
32634: douta=16'hab89;
32635: douta=16'ha388;
32636: douta=16'hab89;
32637: douta=16'ha388;
32638: douta=16'ha389;
32639: douta=16'ha368;
32640: douta=16'ha4d5;
32641: douta=16'hacf4;
32642: douta=16'h8c95;
32643: douta=16'h94d6;
32644: douta=16'h39a7;
32645: douta=16'h2082;
32646: douta=16'h2904;
32647: douta=16'h28e3;
32648: douta=16'h28e3;
32649: douta=16'h28e3;
32650: douta=16'h28e3;
32651: douta=16'h28e3;
32652: douta=16'h28e3;
32653: douta=16'h28e3;
32654: douta=16'h20c3;
32655: douta=16'h20a2;
32656: douta=16'h2082;
32657: douta=16'h20c2;
32658: douta=16'h20a2;
32659: douta=16'h20c2;
32660: douta=16'h28c3;
32661: douta=16'h28c3;
32662: douta=16'h28e3;
32663: douta=16'h28e2;
32664: douta=16'h28e2;
32665: douta=16'h3103;
32666: douta=16'h3103;
32667: douta=16'h3923;
32668: douta=16'h4123;
32669: douta=16'h4143;
32670: douta=16'h4143;
32671: douta=16'h41c7;
32672: douta=16'h31a7;
32673: douta=16'h20c4;
32674: douta=16'h59c4;
32675: douta=16'h59c4;
32676: douta=16'h61c4;
32677: douta=16'h6a24;
32678: douta=16'h6204;
32679: douta=16'h6a04;
32680: douta=16'h7223;
32681: douta=16'h6a46;
32682: douta=16'hb550;
32683: douta=16'h7a85;
32684: douta=16'h7a85;
32685: douta=16'h7a85;
32686: douta=16'h82a6;
32687: douta=16'h8aa6;
32688: douta=16'h8aa6;
32689: douta=16'h8ac6;
32690: douta=16'h8ac6;
32691: douta=16'h8ac6;
32692: douta=16'h9307;
32693: douta=16'h9306;
32694: douta=16'h9327;
32695: douta=16'h51e5;
32696: douta=16'h7265;
32697: douta=16'h92e4;
32698: douta=16'h8243;
32699: douta=16'h7a23;
32700: douta=16'h7202;
32701: douta=16'h92c4;
32702: douta=16'haba6;
32703: douta=16'hb3a7;
32704: douta=16'hb3c7;
32705: douta=16'hb3e7;
32706: douta=16'hbbe7;
32707: douta=16'hbc07;
32708: douta=16'hbc07;
32709: douta=16'hbc07;
32710: douta=16'hbc08;
32711: douta=16'hc428;
32712: douta=16'hbc07;
32713: douta=16'hc428;
32714: douta=16'hc427;
32715: douta=16'hc448;
32716: douta=16'hc448;
32717: douta=16'hc448;
32718: douta=16'hcc48;
32719: douta=16'hc448;
32720: douta=16'hc448;
32721: douta=16'hcc48;
32722: douta=16'hc448;
32723: douta=16'hcc68;
32724: douta=16'hcc68;
32725: douta=16'hcc67;
32726: douta=16'hcc68;
32727: douta=16'hcc67;
32728: douta=16'hcc67;
32729: douta=16'hcc68;
32730: douta=16'hcc68;
32731: douta=16'hcc67;
32732: douta=16'hcc68;
32733: douta=16'hcc68;
32734: douta=16'hcc68;
32735: douta=16'hcc68;
32736: douta=16'hcc88;
32737: douta=16'hcc68;
32738: douta=16'hcc89;
32739: douta=16'hcc68;
32740: douta=16'hcc69;
32741: douta=16'hcc89;
32742: douta=16'hcc69;
32743: douta=16'hcc69;
32744: douta=16'hcc89;
32745: douta=16'hcc89;
32746: douta=16'hcc69;
32747: douta=16'hcc89;
32748: douta=16'hcc89;
32749: douta=16'hcc89;
32750: douta=16'hcc69;
32751: douta=16'hcc89;
32752: douta=16'hcc89;
32753: douta=16'hcc89;
32754: douta=16'hcc89;
32755: douta=16'hd489;
32756: douta=16'hcc69;
32757: douta=16'hcc89;
32758: douta=16'hcc89;
32759: douta=16'hcc89;
32760: douta=16'hcc69;
32761: douta=16'hd468;
32762: douta=16'had73;
32763: douta=16'he6b7;
32764: douta=16'hcc69;
32765: douta=16'hcc69;
32766: douta=16'hcc69;
32767: douta=16'hcc69;
32768: douta=16'hcc69;
32769: douta=16'hcc69;
32770: douta=16'hcc69;
32771: douta=16'hcc69;
32772: douta=16'hcc69;
32773: douta=16'hcc69;
32774: douta=16'hcc69;
32775: douta=16'hcc69;
32776: douta=16'hcc69;
32777: douta=16'hcc69;
32778: douta=16'hcc49;
32779: douta=16'hcc69;
32780: douta=16'hcc69;
32781: douta=16'hcc49;
32782: douta=16'hcc69;
32783: douta=16'hcc69;
32784: douta=16'hc449;
32785: douta=16'hcc69;
32786: douta=16'hcc49;
32787: douta=16'hcc49;
32788: douta=16'hc449;
32789: douta=16'hc449;
32790: douta=16'hc428;
32791: douta=16'hc429;
32792: douta=16'hc429;
32793: douta=16'hc429;
32794: douta=16'hc429;
32795: douta=16'hc429;
32796: douta=16'hc429;
32797: douta=16'hc429;
32798: douta=16'hbc09;
32799: douta=16'hbc29;
32800: douta=16'hbc09;
32801: douta=16'hbc09;
32802: douta=16'hbc09;
32803: douta=16'hbbe9;
32804: douta=16'hbbe9;
32805: douta=16'hbbe9;
32806: douta=16'hb3e8;
32807: douta=16'hbbe9;
32808: douta=16'hb3e8;
32809: douta=16'hb3c8;
32810: douta=16'hb3e9;
32811: douta=16'hb3c8;
32812: douta=16'hb3c9;
32813: douta=16'hb3c8;
32814: douta=16'hb3c9;
32815: douta=16'hb3c9;
32816: douta=16'hb3c8;
32817: douta=16'hb3c8;
32818: douta=16'haba9;
32819: douta=16'haba9;
32820: douta=16'haba9;
32821: douta=16'haba9;
32822: douta=16'haba9;
32823: douta=16'haba9;
32824: douta=16'haba9;
32825: douta=16'hab88;
32826: douta=16'hab88;
32827: douta=16'hab89;
32828: douta=16'ha389;
32829: douta=16'ha389;
32830: douta=16'ha389;
32831: douta=16'ha368;
32832: douta=16'ha4f5;
32833: douta=16'ha4f5;
32834: douta=16'h8cb6;
32835: douta=16'h8c95;
32836: douta=16'h20c3;
32837: douta=16'h28c3;
32838: douta=16'h28e3;
32839: douta=16'h28e3;
32840: douta=16'h28e3;
32841: douta=16'h28e3;
32842: douta=16'h28e3;
32843: douta=16'h28e3;
32844: douta=16'h20c3;
32845: douta=16'h20a3;
32846: douta=16'h20e3;
32847: douta=16'h20c2;
32848: douta=16'h20a2;
32849: douta=16'h20a2;
32850: douta=16'h20a2;
32851: douta=16'h28e3;
32852: douta=16'h28c3;
32853: douta=16'h28c2;
32854: douta=16'h28e3;
32855: douta=16'h28e3;
32856: douta=16'h3103;
32857: douta=16'h3103;
32858: douta=16'h3103;
32859: douta=16'h3923;
32860: douta=16'h4124;
32861: douta=16'h4163;
32862: douta=16'h4964;
32863: douta=16'h4a08;
32864: douta=16'h2967;
32865: douta=16'h28e4;
32866: douta=16'h59c4;
32867: douta=16'h61c4;
32868: douta=16'h61c4;
32869: douta=16'h6204;
32870: douta=16'h6a24;
32871: douta=16'h6a24;
32872: douta=16'h7224;
32873: douta=16'h6aa8;
32874: douta=16'haccf;
32875: douta=16'h7a85;
32876: douta=16'h7a85;
32877: douta=16'h7a85;
32878: douta=16'h82a6;
32879: douta=16'h82c6;
32880: douta=16'h8ac6;
32881: douta=16'h82c6;
32882: douta=16'h8ac6;
32883: douta=16'h8ae6;
32884: douta=16'h8ae6;
32885: douta=16'h9306;
32886: douta=16'h9b27;
32887: douta=16'h7285;
32888: douta=16'h51c5;
32889: douta=16'ha3c9;
32890: douta=16'h93aa;
32891: douta=16'h940c;
32892: douta=16'ha46d;
32893: douta=16'h7329;
32894: douta=16'hbbe7;
32895: douta=16'hb3a7;
32896: douta=16'hb3c6;
32897: douta=16'hb3e7;
32898: douta=16'hbbe7;
32899: douta=16'hbbe7;
32900: douta=16'hbc07;
32901: douta=16'hbc08;
32902: douta=16'hc428;
32903: douta=16'hc428;
32904: douta=16'hc428;
32905: douta=16'hc428;
32906: douta=16'hc428;
32907: douta=16'hc428;
32908: douta=16'hc448;
32909: douta=16'hc448;
32910: douta=16'hcc48;
32911: douta=16'hc448;
32912: douta=16'hcc48;
32913: douta=16'hcc48;
32914: douta=16'hcc68;
32915: douta=16'hcc69;
32916: douta=16'hcc69;
32917: douta=16'hcc68;
32918: douta=16'hcc68;
32919: douta=16'hcc68;
32920: douta=16'hcc68;
32921: douta=16'hcc68;
32922: douta=16'hcc69;
32923: douta=16'hcc68;
32924: douta=16'hcc68;
32925: douta=16'hcc68;
32926: douta=16'hcc88;
32927: douta=16'hcc68;
32928: douta=16'hcc88;
32929: douta=16'hcc89;
32930: douta=16'hcc89;
32931: douta=16'hcc89;
32932: douta=16'hcc89;
32933: douta=16'hcc69;
32934: douta=16'hcc8a;
32935: douta=16'hcc89;
32936: douta=16'hcc69;
32937: douta=16'hcc69;
32938: douta=16'hcc69;
32939: douta=16'hcc69;
32940: douta=16'hcc89;
32941: douta=16'hcc69;
32942: douta=16'hcc89;
32943: douta=16'hcc89;
32944: douta=16'hcc8a;
32945: douta=16'hcc89;
32946: douta=16'hcc89;
32947: douta=16'hd489;
32948: douta=16'hd489;
32949: douta=16'hcc69;
32950: douta=16'hcc89;
32951: douta=16'hcc89;
32952: douta=16'hcc89;
32953: douta=16'hd468;
32954: douta=16'had73;
32955: douta=16'he696;
32956: douta=16'hcc69;
32957: douta=16'hcc68;
32958: douta=16'hcc69;
32959: douta=16'hcc69;
32960: douta=16'hcc69;
32961: douta=16'hcc69;
32962: douta=16'hcc69;
32963: douta=16'hcc69;
32964: douta=16'hcc69;
32965: douta=16'hcc69;
32966: douta=16'hcc69;
32967: douta=16'hcc69;
32968: douta=16'hcc69;
32969: douta=16'hcc69;
32970: douta=16'hcc69;
32971: douta=16'hcc69;
32972: douta=16'hcc69;
32973: douta=16'hcc69;
32974: douta=16'hc449;
32975: douta=16'hcc69;
32976: douta=16'hc449;
32977: douta=16'hcc49;
32978: douta=16'hcc49;
32979: douta=16'hcc49;
32980: douta=16'hc449;
32981: douta=16'hc449;
32982: douta=16'hc449;
32983: douta=16'hc429;
32984: douta=16'hc429;
32985: douta=16'hc429;
32986: douta=16'hc429;
32987: douta=16'hc429;
32988: douta=16'hc429;
32989: douta=16'hbc29;
32990: douta=16'hbc09;
32991: douta=16'hbc29;
32992: douta=16'hbc09;
32993: douta=16'hbc09;
32994: douta=16'hbbe9;
32995: douta=16'hbbe9;
32996: douta=16'hbbe9;
32997: douta=16'hbc09;
32998: douta=16'hbc09;
32999: douta=16'hb3e8;
33000: douta=16'hbbe9;
33001: douta=16'hb3e9;
33002: douta=16'hb3e9;
33003: douta=16'hb3c8;
33004: douta=16'hb3c9;
33005: douta=16'hb3c9;
33006: douta=16'hb3c9;
33007: douta=16'hb3c9;
33008: douta=16'hb3c9;
33009: douta=16'hb3c8;
33010: douta=16'habc9;
33011: douta=16'haba9;
33012: douta=16'hb3c8;
33013: douta=16'haba9;
33014: douta=16'haba9;
33015: douta=16'hab89;
33016: douta=16'haba9;
33017: douta=16'hab89;
33018: douta=16'haba9;
33019: douta=16'ha389;
33020: douta=16'hab89;
33021: douta=16'ha389;
33022: douta=16'hab89;
33023: douta=16'ha368;
33024: douta=16'hb556;
33025: douta=16'h94b5;
33026: douta=16'h94f6;
33027: douta=16'h94f7;
33028: douta=16'h2904;
33029: douta=16'h2904;
33030: douta=16'h20e3;
33031: douta=16'h2904;
33032: douta=16'h28e3;
33033: douta=16'h2903;
33034: douta=16'h28e3;
33035: douta=16'h28e3;
33036: douta=16'h20e3;
33037: douta=16'h20e3;
33038: douta=16'h20c3;
33039: douta=16'h20e3;
33040: douta=16'h20a2;
33041: douta=16'h20a2;
33042: douta=16'h20a2;
33043: douta=16'h20a2;
33044: douta=16'h20a2;
33045: douta=16'h28e3;
33046: douta=16'h28e3;
33047: douta=16'h28e3;
33048: douta=16'h3103;
33049: douta=16'h3123;
33050: douta=16'h3923;
33051: douta=16'h3943;
33052: douta=16'h4143;
33053: douta=16'h4964;
33054: douta=16'h4964;
33055: douta=16'h528b;
33056: douta=16'h10e5;
33057: douta=16'h4985;
33058: douta=16'h59c4;
33059: douta=16'h59c4;
33060: douta=16'h61e4;
33061: douta=16'h6a24;
33062: douta=16'h6a04;
33063: douta=16'h6a24;
33064: douta=16'h7265;
33065: douta=16'h83ee;
33066: douta=16'h8327;
33067: douta=16'h8286;
33068: douta=16'h8285;
33069: douta=16'h8285;
33070: douta=16'h82c6;
33071: douta=16'h82c6;
33072: douta=16'h82c6;
33073: douta=16'h8ac6;
33074: douta=16'h8b07;
33075: douta=16'h8ac6;
33076: douta=16'h9307;
33077: douta=16'h9306;
33078: douta=16'h9326;
33079: douta=16'h9b27;
33080: douta=16'ha347;
33081: douta=16'h93ee;
33082: douta=16'hde76;
33083: douta=16'hc551;
33084: douta=16'he696;
33085: douta=16'h6267;
33086: douta=16'hb3e7;
33087: douta=16'haba7;
33088: douta=16'hb3e7;
33089: douta=16'hb3e7;
33090: douta=16'hb3e7;
33091: douta=16'hbbe7;
33092: douta=16'hbc07;
33093: douta=16'hbc07;
33094: douta=16'hbc07;
33095: douta=16'hc407;
33096: douta=16'hc407;
33097: douta=16'hc428;
33098: douta=16'hc428;
33099: douta=16'hc428;
33100: douta=16'hc448;
33101: douta=16'hc448;
33102: douta=16'hc448;
33103: douta=16'hcc48;
33104: douta=16'hcc48;
33105: douta=16'hcc48;
33106: douta=16'hcc68;
33107: douta=16'hcc68;
33108: douta=16'hcc68;
33109: douta=16'hcc67;
33110: douta=16'hcc68;
33111: douta=16'hcc68;
33112: douta=16'hcc68;
33113: douta=16'hcc68;
33114: douta=16'hcc68;
33115: douta=16'hcc68;
33116: douta=16'hcc88;
33117: douta=16'hcc68;
33118: douta=16'hcc68;
33119: douta=16'hcc69;
33120: douta=16'hcc69;
33121: douta=16'hcc68;
33122: douta=16'hcc69;
33123: douta=16'hcc89;
33124: douta=16'hd489;
33125: douta=16'hcc69;
33126: douta=16'hcc89;
33127: douta=16'hcc89;
33128: douta=16'hcc69;
33129: douta=16'hcc89;
33130: douta=16'hcc89;
33131: douta=16'hcc8a;
33132: douta=16'hcc69;
33133: douta=16'hcc89;
33134: douta=16'hcc8a;
33135: douta=16'hcc89;
33136: douta=16'hcc89;
33137: douta=16'hcc8a;
33138: douta=16'hcc89;
33139: douta=16'hcc89;
33140: douta=16'hcc89;
33141: douta=16'hcc89;
33142: douta=16'hcc89;
33143: douta=16'hcc89;
33144: douta=16'hcc89;
33145: douta=16'hd488;
33146: douta=16'had74;
33147: douta=16'he696;
33148: douta=16'hcc89;
33149: douta=16'hcc89;
33150: douta=16'hcc69;
33151: douta=16'hcc69;
33152: douta=16'hcc69;
33153: douta=16'hcc69;
33154: douta=16'hcc69;
33155: douta=16'hcc69;
33156: douta=16'hcc69;
33157: douta=16'hcc69;
33158: douta=16'hcc69;
33159: douta=16'hcc69;
33160: douta=16'hcc69;
33161: douta=16'hcc69;
33162: douta=16'hcc69;
33163: douta=16'hcc69;
33164: douta=16'hcc49;
33165: douta=16'hcc69;
33166: douta=16'hc468;
33167: douta=16'hcc69;
33168: douta=16'hcc49;
33169: douta=16'hc449;
33170: douta=16'hc449;
33171: douta=16'hc449;
33172: douta=16'hc449;
33173: douta=16'hc449;
33174: douta=16'hc429;
33175: douta=16'hc429;
33176: douta=16'hc429;
33177: douta=16'hc429;
33178: douta=16'hc429;
33179: douta=16'hbc29;
33180: douta=16'hc429;
33181: douta=16'hc429;
33182: douta=16'hc429;
33183: douta=16'hbc09;
33184: douta=16'hc429;
33185: douta=16'hbc09;
33186: douta=16'hbc29;
33187: douta=16'hbc09;
33188: douta=16'hbbe9;
33189: douta=16'hbc09;
33190: douta=16'hbbe9;
33191: douta=16'hbc09;
33192: douta=16'hbbe9;
33193: douta=16'hb3e9;
33194: douta=16'hb3e9;
33195: douta=16'hb3c8;
33196: douta=16'hb3c9;
33197: douta=16'hb3c9;
33198: douta=16'hb3c9;
33199: douta=16'hb3c9;
33200: douta=16'hb3c9;
33201: douta=16'hb3c9;
33202: douta=16'haba9;
33203: douta=16'hb3c9;
33204: douta=16'haba9;
33205: douta=16'haba9;
33206: douta=16'haba9;
33207: douta=16'haba9;
33208: douta=16'haba9;
33209: douta=16'haba9;
33210: douta=16'haba8;
33211: douta=16'hab89;
33212: douta=16'hab89;
33213: douta=16'hab89;
33214: douta=16'ha388;
33215: douta=16'ha388;
33216: douta=16'ha515;
33217: douta=16'h94d6;
33218: douta=16'h94f7;
33219: douta=16'h8454;
33220: douta=16'h2924;
33221: douta=16'h28e3;
33222: douta=16'h28e3;
33223: douta=16'h28e3;
33224: douta=16'h28e3;
33225: douta=16'h28e3;
33226: douta=16'h28e3;
33227: douta=16'h28e3;
33228: douta=16'h20c3;
33229: douta=16'h20e3;
33230: douta=16'h20e3;
33231: douta=16'h2904;
33232: douta=16'h20a2;
33233: douta=16'h20c2;
33234: douta=16'h20c2;
33235: douta=16'h28c3;
33236: douta=16'h28e3;
33237: douta=16'h28e2;
33238: douta=16'h2903;
33239: douta=16'h28e3;
33240: douta=16'h3103;
33241: douta=16'h3123;
33242: douta=16'h3123;
33243: douta=16'h4144;
33244: douta=16'h4143;
33245: douta=16'h4963;
33246: douta=16'h4964;
33247: douta=16'h528a;
33248: douta=16'h0884;
33249: douta=16'h59c4;
33250: douta=16'h59c4;
33251: douta=16'h59c4;
33252: douta=16'h61e4;
33253: douta=16'h61e4;
33254: douta=16'h6a24;
33255: douta=16'h6a04;
33256: douta=16'h7266;
33257: douta=16'h9cd1;
33258: douta=16'h7244;
33259: douta=16'h7a85;
33260: douta=16'h7a85;
33261: douta=16'h7a85;
33262: douta=16'h82a5;
33263: douta=16'h82c6;
33264: douta=16'h8ae6;
33265: douta=16'h8ac6;
33266: douta=16'h8ae6;
33267: douta=16'h8ae7;
33268: douta=16'h9307;
33269: douta=16'h9306;
33270: douta=16'h9b27;
33271: douta=16'h9b28;
33272: douta=16'h8aa5;
33273: douta=16'hd6b7;
33274: douta=16'h0000;
33275: douta=16'h0000;
33276: douta=16'h934a;
33277: douta=16'h59c4;
33278: douta=16'hb3c7;
33279: douta=16'hb3c7;
33280: douta=16'hb3e7;
33281: douta=16'hb3e7;
33282: douta=16'hb3e8;
33283: douta=16'hbbe7;
33284: douta=16'hbc07;
33285: douta=16'hbc08;
33286: douta=16'hc407;
33287: douta=16'hc428;
33288: douta=16'hc428;
33289: douta=16'hc428;
33290: douta=16'hc428;
33291: douta=16'hc428;
33292: douta=16'hc448;
33293: douta=16'hc448;
33294: douta=16'hc448;
33295: douta=16'hcc49;
33296: douta=16'hcc49;
33297: douta=16'hcc49;
33298: douta=16'hc448;
33299: douta=16'hcc68;
33300: douta=16'hcc68;
33301: douta=16'hcc68;
33302: douta=16'hcc68;
33303: douta=16'hcc68;
33304: douta=16'hcc68;
33305: douta=16'hcc68;
33306: douta=16'hcc68;
33307: douta=16'hcc68;
33308: douta=16'hcc68;
33309: douta=16'hcc68;
33310: douta=16'hcc69;
33311: douta=16'hcc69;
33312: douta=16'hcc89;
33313: douta=16'hcc89;
33314: douta=16'hcc89;
33315: douta=16'hcc89;
33316: douta=16'hcc69;
33317: douta=16'hcc8a;
33318: douta=16'hcc69;
33319: douta=16'hcc69;
33320: douta=16'hcc89;
33321: douta=16'hcc89;
33322: douta=16'hcc69;
33323: douta=16'hcc89;
33324: douta=16'hcc89;
33325: douta=16'hcc89;
33326: douta=16'hcc8a;
33327: douta=16'hcc69;
33328: douta=16'hcc8a;
33329: douta=16'hcc89;
33330: douta=16'hcc89;
33331: douta=16'hcc69;
33332: douta=16'hcc89;
33333: douta=16'hcc69;
33334: douta=16'hcc89;
33335: douta=16'hcc89;
33336: douta=16'hcc89;
33337: douta=16'hd488;
33338: douta=16'hb594;
33339: douta=16'he696;
33340: douta=16'hcc69;
33341: douta=16'hcc69;
33342: douta=16'hcc89;
33343: douta=16'hcc69;
33344: douta=16'hcc69;
33345: douta=16'hcc69;
33346: douta=16'hcc69;
33347: douta=16'hcc89;
33348: douta=16'hcc69;
33349: douta=16'hcc69;
33350: douta=16'hcc69;
33351: douta=16'hcc69;
33352: douta=16'hcc69;
33353: douta=16'hcc69;
33354: douta=16'hcc49;
33355: douta=16'hcc49;
33356: douta=16'hcc69;
33357: douta=16'hcc49;
33358: douta=16'hcc69;
33359: douta=16'hcc49;
33360: douta=16'hc449;
33361: douta=16'hc449;
33362: douta=16'hc449;
33363: douta=16'hc449;
33364: douta=16'hc429;
33365: douta=16'hc429;
33366: douta=16'hc429;
33367: douta=16'hc449;
33368: douta=16'hc449;
33369: douta=16'hc449;
33370: douta=16'hbc29;
33371: douta=16'hc429;
33372: douta=16'hbc09;
33373: douta=16'hbc29;
33374: douta=16'hbc29;
33375: douta=16'hbc09;
33376: douta=16'hbc09;
33377: douta=16'hbc09;
33378: douta=16'hbc09;
33379: douta=16'hbc09;
33380: douta=16'hbc09;
33381: douta=16'hbbe9;
33382: douta=16'hbc0a;
33383: douta=16'hb3e9;
33384: douta=16'hbbe9;
33385: douta=16'hb3c9;
33386: douta=16'hbc09;
33387: douta=16'hb3e9;
33388: douta=16'hb3c9;
33389: douta=16'hb3e9;
33390: douta=16'hb3c9;
33391: douta=16'hb3c9;
33392: douta=16'hb3c9;
33393: douta=16'hb3c9;
33394: douta=16'habc9;
33395: douta=16'haba9;
33396: douta=16'habc9;
33397: douta=16'habc9;
33398: douta=16'haba9;
33399: douta=16'haba9;
33400: douta=16'hab89;
33401: douta=16'haba8;
33402: douta=16'haba8;
33403: douta=16'hab89;
33404: douta=16'haba9;
33405: douta=16'ha389;
33406: douta=16'hab89;
33407: douta=16'ha389;
33408: douta=16'h9cd5;
33409: douta=16'h94d6;
33410: douta=16'h94b6;
33411: douta=16'h638f;
33412: douta=16'h2903;
33413: douta=16'h2904;
33414: douta=16'h28e4;
33415: douta=16'h28e3;
33416: douta=16'h28e3;
33417: douta=16'h28e3;
33418: douta=16'h28e3;
33419: douta=16'h28e3;
33420: douta=16'h20e3;
33421: douta=16'h20e3;
33422: douta=16'h20e3;
33423: douta=16'h2904;
33424: douta=16'h20c2;
33425: douta=16'h20c2;
33426: douta=16'h20c2;
33427: douta=16'h28e3;
33428: douta=16'h28c3;
33429: douta=16'h28e3;
33430: douta=16'h28e3;
33431: douta=16'h3103;
33432: douta=16'h3103;
33433: douta=16'h3923;
33434: douta=16'h3923;
33435: douta=16'h3943;
33436: douta=16'h4143;
33437: douta=16'h4964;
33438: douta=16'h4964;
33439: douta=16'h4a6a;
33440: douta=16'h0885;
33441: douta=16'h59c4;
33442: douta=16'h59c4;
33443: douta=16'h59e4;
33444: douta=16'h61e4;
33445: douta=16'h61e4;
33446: douta=16'h6a24;
33447: douta=16'h6a25;
33448: douta=16'h72a8;
33449: douta=16'ha513;
33450: douta=16'h7204;
33451: douta=16'h7a85;
33452: douta=16'h82a5;
33453: douta=16'h7a85;
33454: douta=16'h82c6;
33455: douta=16'h82c6;
33456: douta=16'h8ac6;
33457: douta=16'h8ac6;
33458: douta=16'h8ac6;
33459: douta=16'h8b06;
33460: douta=16'h9307;
33461: douta=16'h9326;
33462: douta=16'h9b27;
33463: douta=16'h9b27;
33464: douta=16'h92c4;
33465: douta=16'hf71a;
33466: douta=16'h4a28;
33467: douta=16'h0000;
33468: douta=16'h8b4a;
33469: douta=16'h59c3;
33470: douta=16'hb3a8;
33471: douta=16'hb3c7;
33472: douta=16'hb3e7;
33473: douta=16'hb3c7;
33474: douta=16'hbbe8;
33475: douta=16'hbc07;
33476: douta=16'hbc07;
33477: douta=16'hbc07;
33478: douta=16'hbc07;
33479: douta=16'hc428;
33480: douta=16'hc428;
33481: douta=16'hc428;
33482: douta=16'hc428;
33483: douta=16'hc448;
33484: douta=16'hc448;
33485: douta=16'hc448;
33486: douta=16'hc448;
33487: douta=16'hcc49;
33488: douta=16'hcc49;
33489: douta=16'hcc49;
33490: douta=16'hcc68;
33491: douta=16'hc448;
33492: douta=16'hcc68;
33493: douta=16'hcc68;
33494: douta=16'hcc67;
33495: douta=16'hcc68;
33496: douta=16'hcc68;
33497: douta=16'hcc48;
33498: douta=16'hcc69;
33499: douta=16'hcc68;
33500: douta=16'hcc68;
33501: douta=16'hcc68;
33502: douta=16'hcc69;
33503: douta=16'hcc69;
33504: douta=16'hcc69;
33505: douta=16'hcc69;
33506: douta=16'hcc69;
33507: douta=16'hcc69;
33508: douta=16'hcc89;
33509: douta=16'hcc69;
33510: douta=16'hcc89;
33511: douta=16'hcc89;
33512: douta=16'hcc8a;
33513: douta=16'hcc69;
33514: douta=16'hcc69;
33515: douta=16'hcc89;
33516: douta=16'hcc89;
33517: douta=16'hcc89;
33518: douta=16'hcc89;
33519: douta=16'hcc89;
33520: douta=16'hcc89;
33521: douta=16'hcc8a;
33522: douta=16'hcc89;
33523: douta=16'hcc89;
33524: douta=16'hcc89;
33525: douta=16'hcc69;
33526: douta=16'hcc69;
33527: douta=16'hcc89;
33528: douta=16'hcc89;
33529: douta=16'hd488;
33530: douta=16'had74;
33531: douta=16'he696;
33532: douta=16'hcc69;
33533: douta=16'hcc69;
33534: douta=16'hcc89;
33535: douta=16'hcc69;
33536: douta=16'hcc69;
33537: douta=16'hcc69;
33538: douta=16'hcc49;
33539: douta=16'hcc69;
33540: douta=16'hcc69;
33541: douta=16'hcc69;
33542: douta=16'hcc69;
33543: douta=16'hcc69;
33544: douta=16'hcc69;
33545: douta=16'hcc69;
33546: douta=16'hcc69;
33547: douta=16'hcc49;
33548: douta=16'hcc49;
33549: douta=16'hcc49;
33550: douta=16'hcc49;
33551: douta=16'hcc69;
33552: douta=16'hc449;
33553: douta=16'hc449;
33554: douta=16'hc449;
33555: douta=16'hc449;
33556: douta=16'hc449;
33557: douta=16'hc449;
33558: douta=16'hc429;
33559: douta=16'hc429;
33560: douta=16'hc449;
33561: douta=16'hc429;
33562: douta=16'hc449;
33563: douta=16'hc429;
33564: douta=16'hbc29;
33565: douta=16'hc429;
33566: douta=16'hbc29;
33567: douta=16'hbc29;
33568: douta=16'hbc09;
33569: douta=16'hbc09;
33570: douta=16'hbc29;
33571: douta=16'hbc09;
33572: douta=16'hbbe9;
33573: douta=16'hbc09;
33574: douta=16'hbc09;
33575: douta=16'hbbe9;
33576: douta=16'hbc09;
33577: douta=16'hb3e9;
33578: douta=16'hb3e9;
33579: douta=16'hb3c9;
33580: douta=16'hb3c9;
33581: douta=16'hb3e9;
33582: douta=16'hb3e9;
33583: douta=16'hb3e9;
33584: douta=16'hb3c9;
33585: douta=16'hb3c9;
33586: douta=16'hb3a9;
33587: douta=16'habc9;
33588: douta=16'haba9;
33589: douta=16'hb3c9;
33590: douta=16'haba9;
33591: douta=16'haba9;
33592: douta=16'haba9;
33593: douta=16'haba9;
33594: douta=16'habc9;
33595: douta=16'hab89;
33596: douta=16'haba9;
33597: douta=16'ha389;
33598: douta=16'ha389;
33599: douta=16'ha388;
33600: douta=16'h8c54;
33601: douta=16'h94b6;
33602: douta=16'h8cf7;
33603: douta=16'h20e3;
33604: douta=16'h2904;
33605: douta=16'h28e3;
33606: douta=16'h28e3;
33607: douta=16'h28e3;
33608: douta=16'h28e3;
33609: douta=16'h28e3;
33610: douta=16'h20e3;
33611: douta=16'h20e3;
33612: douta=16'h20e3;
33613: douta=16'h20e3;
33614: douta=16'h20e3;
33615: douta=16'h20e3;
33616: douta=16'h20a2;
33617: douta=16'h20c2;
33618: douta=16'h20c3;
33619: douta=16'h28c3;
33620: douta=16'h28e3;
33621: douta=16'h28e3;
33622: douta=16'h30e3;
33623: douta=16'h3103;
33624: douta=16'h3103;
33625: douta=16'h3923;
33626: douta=16'h3923;
33627: douta=16'h4124;
33628: douta=16'h4143;
33629: douta=16'h4964;
33630: douta=16'h4964;
33631: douta=16'h39c8;
33632: douta=16'h18a4;
33633: douta=16'h59c4;
33634: douta=16'h59e4;
33635: douta=16'h59c4;
33636: douta=16'h61e4;
33637: douta=16'h6a04;
33638: douta=16'h6a24;
33639: douta=16'h6a24;
33640: douta=16'h83ee;
33641: douta=16'hb573;
33642: douta=16'h7203;
33643: douta=16'h7a85;
33644: douta=16'h7a85;
33645: douta=16'h7a85;
33646: douta=16'h82c6;
33647: douta=16'h82c6;
33648: douta=16'h8ac6;
33649: douta=16'h8ae6;
33650: douta=16'h8ae6;
33651: douta=16'h8ae7;
33652: douta=16'h9307;
33653: douta=16'h9b27;
33654: douta=16'h9b47;
33655: douta=16'h9306;
33656: douta=16'ha387;
33657: douta=16'hde37;
33658: douta=16'h5269;
33659: douta=16'hde96;
33660: douta=16'hde55;
33661: douta=16'h79e2;
33662: douta=16'hb3c8;
33663: douta=16'haba7;
33664: douta=16'hb3e8;
33665: douta=16'hb3e7;
33666: douta=16'hbbe8;
33667: douta=16'hbc07;
33668: douta=16'hbc07;
33669: douta=16'hbc08;
33670: douta=16'hc407;
33671: douta=16'hc407;
33672: douta=16'hbc07;
33673: douta=16'hc448;
33674: douta=16'hc428;
33675: douta=16'hc448;
33676: douta=16'hc448;
33677: douta=16'hc448;
33678: douta=16'hc448;
33679: douta=16'hc448;
33680: douta=16'hc449;
33681: douta=16'hcc49;
33682: douta=16'hc448;
33683: douta=16'hc448;
33684: douta=16'hcc68;
33685: douta=16'hcc68;
33686: douta=16'hcc68;
33687: douta=16'hcc68;
33688: douta=16'hcc69;
33689: douta=16'hcc68;
33690: douta=16'hcc69;
33691: douta=16'hcc68;
33692: douta=16'hcc69;
33693: douta=16'hcc69;
33694: douta=16'hcc69;
33695: douta=16'hcc68;
33696: douta=16'hcc69;
33697: douta=16'hcc69;
33698: douta=16'hcc69;
33699: douta=16'hcc69;
33700: douta=16'hcc89;
33701: douta=16'hcc69;
33702: douta=16'hcc89;
33703: douta=16'hcc89;
33704: douta=16'hcc89;
33705: douta=16'hcc89;
33706: douta=16'hcc69;
33707: douta=16'hcc89;
33708: douta=16'hcc89;
33709: douta=16'hcc89;
33710: douta=16'hcc89;
33711: douta=16'hcc8a;
33712: douta=16'hcc89;
33713: douta=16'hcc89;
33714: douta=16'hcc89;
33715: douta=16'hcc69;
33716: douta=16'hcc69;
33717: douta=16'hcc89;
33718: douta=16'hcc69;
33719: douta=16'hcc69;
33720: douta=16'hcc69;
33721: douta=16'hd488;
33722: douta=16'hb594;
33723: douta=16'hde76;
33724: douta=16'hcc69;
33725: douta=16'hcc69;
33726: douta=16'hcc69;
33727: douta=16'hcc69;
33728: douta=16'hcc69;
33729: douta=16'hcc69;
33730: douta=16'hcc69;
33731: douta=16'hcc69;
33732: douta=16'hcc69;
33733: douta=16'hcc69;
33734: douta=16'hcc69;
33735: douta=16'hcc69;
33736: douta=16'hcc6a;
33737: douta=16'hcc69;
33738: douta=16'hcc69;
33739: douta=16'hcc69;
33740: douta=16'hc449;
33741: douta=16'hc449;
33742: douta=16'hc449;
33743: douta=16'hc448;
33744: douta=16'hc449;
33745: douta=16'hcc49;
33746: douta=16'hc449;
33747: douta=16'hc449;
33748: douta=16'hc429;
33749: douta=16'hc429;
33750: douta=16'hc429;
33751: douta=16'hc429;
33752: douta=16'hc429;
33753: douta=16'hc449;
33754: douta=16'hc429;
33755: douta=16'hc429;
33756: douta=16'hc429;
33757: douta=16'hbc09;
33758: douta=16'hbc09;
33759: douta=16'hbc09;
33760: douta=16'hc429;
33761: douta=16'hbc09;
33762: douta=16'hbc09;
33763: douta=16'hbc09;
33764: douta=16'hbc09;
33765: douta=16'hbc09;
33766: douta=16'hbc09;
33767: douta=16'hbbe9;
33768: douta=16'hbbe9;
33769: douta=16'hb3e9;
33770: douta=16'hbbe9;
33771: douta=16'hb3e9;
33772: douta=16'hb3e9;
33773: douta=16'hb3c9;
33774: douta=16'hbbe9;
33775: douta=16'hb3e9;
33776: douta=16'hb3c9;
33777: douta=16'hb3c8;
33778: douta=16'hb3a9;
33779: douta=16'hb3ca;
33780: douta=16'haba9;
33781: douta=16'haba9;
33782: douta=16'haba9;
33783: douta=16'hb3c9;
33784: douta=16'haba9;
33785: douta=16'haba9;
33786: douta=16'haba9;
33787: douta=16'ha388;
33788: douta=16'ha389;
33789: douta=16'ha389;
33790: douta=16'ha389;
33791: douta=16'ha389;
33792: douta=16'h8c95;
33793: douta=16'h94b6;
33794: douta=16'h9518;
33795: douta=16'h2061;
33796: douta=16'h3104;
33797: douta=16'h28e3;
33798: douta=16'h28e3;
33799: douta=16'h20e3;
33800: douta=16'h28e3;
33801: douta=16'h28e3;
33802: douta=16'h20e3;
33803: douta=16'h20e3;
33804: douta=16'h28e3;
33805: douta=16'h20c3;
33806: douta=16'h28e3;
33807: douta=16'h18a2;
33808: douta=16'h20a2;
33809: douta=16'h20c3;
33810: douta=16'h20c2;
33811: douta=16'h28c3;
33812: douta=16'h28e3;
33813: douta=16'h28e3;
33814: douta=16'h3103;
33815: douta=16'h3103;
33816: douta=16'h3123;
33817: douta=16'h3943;
33818: douta=16'h3923;
33819: douta=16'h4144;
33820: douta=16'h4163;
33821: douta=16'h4964;
33822: douta=16'h4964;
33823: douta=16'h2967;
33824: douta=16'h3104;
33825: douta=16'h59c4;
33826: douta=16'h59e4;
33827: douta=16'h61e4;
33828: douta=16'h61e4;
33829: douta=16'h6a24;
33830: douta=16'h7245;
33831: douta=16'h7224;
33832: douta=16'h9cf2;
33833: douta=16'hacf0;
33834: douta=16'h7a64;
33835: douta=16'h7a85;
33836: douta=16'h7a85;
33837: douta=16'h82a5;
33838: douta=16'h82c6;
33839: douta=16'h82c6;
33840: douta=16'h8ac6;
33841: douta=16'h8ac6;
33842: douta=16'h8ae6;
33843: douta=16'h92e6;
33844: douta=16'h9307;
33845: douta=16'h9b27;
33846: douta=16'h9b47;
33847: douta=16'h92c6;
33848: douta=16'hac4b;
33849: douta=16'he6d7;
33850: douta=16'h29e7;
33851: douta=16'hb44e;
33852: douta=16'heef8;
33853: douta=16'h9ae4;
33854: douta=16'haba7;
33855: douta=16'haba7;
33856: douta=16'hb3e7;
33857: douta=16'hbbe8;
33858: douta=16'hb3e7;
33859: douta=16'hbc07;
33860: douta=16'hbc08;
33861: douta=16'hbc08;
33862: douta=16'hc407;
33863: douta=16'hc407;
33864: douta=16'hc428;
33865: douta=16'hc428;
33866: douta=16'hc448;
33867: douta=16'hc428;
33868: douta=16'hc448;
33869: douta=16'hcc49;
33870: douta=16'hc448;
33871: douta=16'hc448;
33872: douta=16'hc449;
33873: douta=16'hc448;
33874: douta=16'hc448;
33875: douta=16'hc448;
33876: douta=16'hc448;
33877: douta=16'hcc68;
33878: douta=16'hcc68;
33879: douta=16'hcc68;
33880: douta=16'hcc68;
33881: douta=16'hcc68;
33882: douta=16'hcc68;
33883: douta=16'hcc69;
33884: douta=16'hcc69;
33885: douta=16'hcc69;
33886: douta=16'hcc69;
33887: douta=16'hcc69;
33888: douta=16'hcc69;
33889: douta=16'hcc69;
33890: douta=16'hcc69;
33891: douta=16'hcc69;
33892: douta=16'hcc69;
33893: douta=16'hcc89;
33894: douta=16'hcc69;
33895: douta=16'hcc89;
33896: douta=16'hcc89;
33897: douta=16'hcc89;
33898: douta=16'hcc89;
33899: douta=16'hcc89;
33900: douta=16'hcc89;
33901: douta=16'hcc89;
33902: douta=16'hcc69;
33903: douta=16'hcc89;
33904: douta=16'hcc89;
33905: douta=16'hcc89;
33906: douta=16'hcc69;
33907: douta=16'hcc89;
33908: douta=16'hcc69;
33909: douta=16'hcc89;
33910: douta=16'hcc69;
33911: douta=16'hcc69;
33912: douta=16'hcc69;
33913: douta=16'hcc68;
33914: douta=16'hb594;
33915: douta=16'he696;
33916: douta=16'hcc89;
33917: douta=16'hcc69;
33918: douta=16'hcc69;
33919: douta=16'hcc69;
33920: douta=16'hcc69;
33921: douta=16'hcc69;
33922: douta=16'hcc69;
33923: douta=16'hcc69;
33924: douta=16'hcc69;
33925: douta=16'hcc69;
33926: douta=16'hcc69;
33927: douta=16'hcc69;
33928: douta=16'hcc69;
33929: douta=16'hcc69;
33930: douta=16'hcc69;
33931: douta=16'hcc69;
33932: douta=16'hcc69;
33933: douta=16'hcc49;
33934: douta=16'hcc69;
33935: douta=16'hc449;
33936: douta=16'hcc69;
33937: douta=16'hc449;
33938: douta=16'hc449;
33939: douta=16'hc449;
33940: douta=16'hc429;
33941: douta=16'hc429;
33942: douta=16'hc449;
33943: douta=16'hc429;
33944: douta=16'hc429;
33945: douta=16'hc429;
33946: douta=16'hc429;
33947: douta=16'hc429;
33948: douta=16'hc429;
33949: douta=16'hbc09;
33950: douta=16'hbc29;
33951: douta=16'hbc29;
33952: douta=16'hbc09;
33953: douta=16'hbc09;
33954: douta=16'hbc09;
33955: douta=16'hbc09;
33956: douta=16'hbc09;
33957: douta=16'hbc09;
33958: douta=16'hbbe9;
33959: douta=16'hbc09;
33960: douta=16'hbc09;
33961: douta=16'hbbe9;
33962: douta=16'hbbe9;
33963: douta=16'hbbe9;
33964: douta=16'hb3e9;
33965: douta=16'hb3e9;
33966: douta=16'hb3e9;
33967: douta=16'hb3c9;
33968: douta=16'hb3c9;
33969: douta=16'hb3c9;
33970: douta=16'haba9;
33971: douta=16'haba9;
33972: douta=16'habc9;
33973: douta=16'haba9;
33974: douta=16'haba9;
33975: douta=16'haba9;
33976: douta=16'habc9;
33977: douta=16'haba9;
33978: douta=16'haba9;
33979: douta=16'haba9;
33980: douta=16'haba9;
33981: douta=16'ha389;
33982: douta=16'ha389;
33983: douta=16'ha389;
33984: douta=16'h8c95;
33985: douta=16'h8c96;
33986: douta=16'h8495;
33987: douta=16'h20a2;
33988: douta=16'h2904;
33989: douta=16'h20e3;
33990: douta=16'h2904;
33991: douta=16'h28e3;
33992: douta=16'h28e3;
33993: douta=16'h28e3;
33994: douta=16'h20e3;
33995: douta=16'h20e3;
33996: douta=16'h20e3;
33997: douta=16'h20c3;
33998: douta=16'h28e3;
33999: douta=16'h18a2;
34000: douta=16'h20a2;
34001: douta=16'h20c2;
34002: douta=16'h28c3;
34003: douta=16'h28e3;
34004: douta=16'h28e3;
34005: douta=16'h28e3;
34006: douta=16'h30e3;
34007: douta=16'h3103;
34008: douta=16'h3103;
34009: douta=16'h3923;
34010: douta=16'h3943;
34011: douta=16'h4164;
34012: douta=16'h4163;
34013: douta=16'h4964;
34014: douta=16'h4144;
34015: douta=16'h2967;
34016: douta=16'h3924;
34017: douta=16'h59c4;
34018: douta=16'h59e4;
34019: douta=16'h61e4;
34020: douta=16'h61e4;
34021: douta=16'h6a24;
34022: douta=16'h6a25;
34023: douta=16'h7245;
34024: douta=16'ha553;
34025: douta=16'ha4af;
34026: douta=16'h7a64;
34027: douta=16'h7a85;
34028: douta=16'h82a5;
34029: douta=16'h82a5;
34030: douta=16'h82c6;
34031: douta=16'h82c6;
34032: douta=16'h8ac6;
34033: douta=16'h8ae7;
34034: douta=16'h8ae7;
34035: douta=16'h9307;
34036: douta=16'h9307;
34037: douta=16'h9326;
34038: douta=16'h9b27;
34039: douta=16'h92c5;
34040: douta=16'hbc8e;
34041: douta=16'hc5d4;
34042: douta=16'h41e6;
34043: douta=16'h8aea;
34044: douta=16'hf739;
34045: douta=16'ha325;
34046: douta=16'hb3c8;
34047: douta=16'hb3c7;
34048: douta=16'hbc08;
34049: douta=16'hbc08;
34050: douta=16'hbc08;
34051: douta=16'hbc07;
34052: douta=16'hbc07;
34053: douta=16'hbc08;
34054: douta=16'hc428;
34055: douta=16'hc428;
34056: douta=16'hc428;
34057: douta=16'hc428;
34058: douta=16'hc448;
34059: douta=16'hc448;
34060: douta=16'hc448;
34061: douta=16'hc448;
34062: douta=16'hc428;
34063: douta=16'hc448;
34064: douta=16'hc448;
34065: douta=16'hc448;
34066: douta=16'hcc68;
34067: douta=16'hcc68;
34068: douta=16'hc448;
34069: douta=16'hcc68;
34070: douta=16'hcc68;
34071: douta=16'hcc68;
34072: douta=16'hcc68;
34073: douta=16'hcc68;
34074: douta=16'hcc69;
34075: douta=16'hcc69;
34076: douta=16'hcc69;
34077: douta=16'hcc68;
34078: douta=16'hcc69;
34079: douta=16'hcc69;
34080: douta=16'hcc69;
34081: douta=16'hcc69;
34082: douta=16'hcc69;
34083: douta=16'hcc69;
34084: douta=16'hcc89;
34085: douta=16'hcc69;
34086: douta=16'hcc89;
34087: douta=16'hcc89;
34088: douta=16'hcc89;
34089: douta=16'hcc89;
34090: douta=16'hcc89;
34091: douta=16'hcc89;
34092: douta=16'hcc89;
34093: douta=16'hcc89;
34094: douta=16'hcc89;
34095: douta=16'hcc89;
34096: douta=16'hcc89;
34097: douta=16'hcc89;
34098: douta=16'hcc89;
34099: douta=16'hcc89;
34100: douta=16'hcc69;
34101: douta=16'hcc69;
34102: douta=16'hcc89;
34103: douta=16'hcc89;
34104: douta=16'hcc69;
34105: douta=16'hcc88;
34106: douta=16'hb594;
34107: douta=16'he696;
34108: douta=16'hcc69;
34109: douta=16'hcc89;
34110: douta=16'hcc68;
34111: douta=16'hcc89;
34112: douta=16'hcc69;
34113: douta=16'hcc69;
34114: douta=16'hcc69;
34115: douta=16'hcc69;
34116: douta=16'hcc69;
34117: douta=16'hcc6a;
34118: douta=16'hcc69;
34119: douta=16'hcc69;
34120: douta=16'hcc69;
34121: douta=16'hcc69;
34122: douta=16'hcc69;
34123: douta=16'hcc69;
34124: douta=16'hc449;
34125: douta=16'hcc49;
34126: douta=16'hcc6a;
34127: douta=16'hc449;
34128: douta=16'hc449;
34129: douta=16'hc449;
34130: douta=16'hc449;
34131: douta=16'hc449;
34132: douta=16'hc429;
34133: douta=16'hc449;
34134: douta=16'hc449;
34135: douta=16'hc429;
34136: douta=16'hc429;
34137: douta=16'hc429;
34138: douta=16'hc44a;
34139: douta=16'hc429;
34140: douta=16'hc429;
34141: douta=16'hc429;
34142: douta=16'hc429;
34143: douta=16'hc429;
34144: douta=16'hbc09;
34145: douta=16'hbc09;
34146: douta=16'hbc09;
34147: douta=16'hbc09;
34148: douta=16'hbbe9;
34149: douta=16'hbc09;
34150: douta=16'hbc09;
34151: douta=16'hb3e9;
34152: douta=16'hb3e9;
34153: douta=16'hbc09;
34154: douta=16'hb3e9;
34155: douta=16'hbbe9;
34156: douta=16'hbbe9;
34157: douta=16'hb3e9;
34158: douta=16'hb3e9;
34159: douta=16'hb3c9;
34160: douta=16'hb3c9;
34161: douta=16'hb3c9;
34162: douta=16'hb3ea;
34163: douta=16'hb3ca;
34164: douta=16'hb3ca;
34165: douta=16'haba9;
34166: douta=16'haba9;
34167: douta=16'haba9;
34168: douta=16'haba9;
34169: douta=16'habc9;
34170: douta=16'haba9;
34171: douta=16'ha388;
34172: douta=16'haba8;
34173: douta=16'ha389;
34174: douta=16'ha389;
34175: douta=16'ha389;
34176: douta=16'h9495;
34177: douta=16'h84b7;
34178: douta=16'h3166;
34179: douta=16'h2904;
34180: douta=16'h2904;
34181: douta=16'h28e3;
34182: douta=16'h28e3;
34183: douta=16'h28e3;
34184: douta=16'h2904;
34185: douta=16'h2904;
34186: douta=16'h20e4;
34187: douta=16'h20e3;
34188: douta=16'h2904;
34189: douta=16'h20e3;
34190: douta=16'h20a2;
34191: douta=16'h20a2;
34192: douta=16'h20c3;
34193: douta=16'h20c2;
34194: douta=16'h28e2;
34195: douta=16'h28e3;
34196: douta=16'h28e3;
34197: douta=16'h28e3;
34198: douta=16'h3103;
34199: douta=16'h3103;
34200: douta=16'h3103;
34201: douta=16'h3944;
34202: douta=16'h3923;
34203: douta=16'h4144;
34204: douta=16'h4163;
34205: douta=16'h4943;
34206: douta=16'h49c6;
34207: douta=16'h10c4;
34208: douta=16'h51a5;
34209: douta=16'h59c4;
34210: douta=16'h6205;
34211: douta=16'h6204;
34212: douta=16'h6205;
34213: douta=16'h6a44;
34214: douta=16'h7245;
34215: douta=16'h7244;
34216: douta=16'hb572;
34217: douta=16'h8b49;
34218: douta=16'h7a85;
34219: douta=16'h7a85;
34220: douta=16'h82a5;
34221: douta=16'h82c6;
34222: douta=16'h82c6;
34223: douta=16'h8ac6;
34224: douta=16'h8ae7;
34225: douta=16'h8b07;
34226: douta=16'h9307;
34227: douta=16'h9307;
34228: douta=16'h9307;
34229: douta=16'h9b27;
34230: douta=16'h9b47;
34231: douta=16'h9b26;
34232: douta=16'hd5b3;
34233: douta=16'hbdd3;
34234: douta=16'h1861;
34235: douta=16'he6d8;
34236: douta=16'heed8;
34237: douta=16'hbbe8;
34238: douta=16'habc7;
34239: douta=16'hb3c7;
34240: douta=16'hb3c8;
34241: douta=16'hb3e7;
34242: douta=16'hbbe8;
34243: douta=16'hbbe8;
34244: douta=16'hbc08;
34245: douta=16'hbc08;
34246: douta=16'hc428;
34247: douta=16'hc408;
34248: douta=16'hc428;
34249: douta=16'hc448;
34250: douta=16'hc428;
34251: douta=16'hc449;
34252: douta=16'hc448;
34253: douta=16'hc448;
34254: douta=16'hc448;
34255: douta=16'hc449;
34256: douta=16'hc448;
34257: douta=16'hcc49;
34258: douta=16'hc449;
34259: douta=16'hcc69;
34260: douta=16'hcc69;
34261: douta=16'hcc69;
34262: douta=16'hcc69;
34263: douta=16'hcc68;
34264: douta=16'hcc69;
34265: douta=16'hcc68;
34266: douta=16'hcc68;
34267: douta=16'hcc69;
34268: douta=16'hcc69;
34269: douta=16'hcc69;
34270: douta=16'hcc69;
34271: douta=16'hcc89;
34272: douta=16'hcc69;
34273: douta=16'hcc69;
34274: douta=16'hcc89;
34275: douta=16'hcc69;
34276: douta=16'hcc89;
34277: douta=16'hcc89;
34278: douta=16'hcc89;
34279: douta=16'hcc89;
34280: douta=16'hcc89;
34281: douta=16'hcc89;
34282: douta=16'hcc89;
34283: douta=16'hcc89;
34284: douta=16'hcc8a;
34285: douta=16'hcc89;
34286: douta=16'hcc69;
34287: douta=16'hcc69;
34288: douta=16'hcc69;
34289: douta=16'hcc89;
34290: douta=16'hcc89;
34291: douta=16'hcc69;
34292: douta=16'hcc69;
34293: douta=16'hcc89;
34294: douta=16'hcc69;
34295: douta=16'hcc89;
34296: douta=16'hcc69;
34297: douta=16'hcc69;
34298: douta=16'hb5b5;
34299: douta=16'he696;
34300: douta=16'hcc6a;
34301: douta=16'hcc69;
34302: douta=16'hcc49;
34303: douta=16'hcc89;
34304: douta=16'hcc69;
34305: douta=16'hcc69;
34306: douta=16'hcc69;
34307: douta=16'hcc69;
34308: douta=16'hcc69;
34309: douta=16'hcc69;
34310: douta=16'hcc69;
34311: douta=16'hcc49;
34312: douta=16'hcc69;
34313: douta=16'hcc49;
34314: douta=16'hcc69;
34315: douta=16'hcc69;
34316: douta=16'hc449;
34317: douta=16'hc449;
34318: douta=16'hc449;
34319: douta=16'hcc49;
34320: douta=16'hc449;
34321: douta=16'hc449;
34322: douta=16'hc429;
34323: douta=16'hc449;
34324: douta=16'hc449;
34325: douta=16'hc429;
34326: douta=16'hc429;
34327: douta=16'hc429;
34328: douta=16'hc429;
34329: douta=16'hc429;
34330: douta=16'hc429;
34331: douta=16'hc44a;
34332: douta=16'hbc09;
34333: douta=16'hbc09;
34334: douta=16'hc429;
34335: douta=16'hc40a;
34336: douta=16'hbc09;
34337: douta=16'hbc09;
34338: douta=16'hbc09;
34339: douta=16'hbc09;
34340: douta=16'hbc09;
34341: douta=16'hbc09;
34342: douta=16'hbc09;
34343: douta=16'hbc09;
34344: douta=16'hbbe9;
34345: douta=16'hbbe9;
34346: douta=16'hbbe9;
34347: douta=16'hbc09;
34348: douta=16'hbbe9;
34349: douta=16'hbbe9;
34350: douta=16'hb3e9;
34351: douta=16'hb3e9;
34352: douta=16'hb3ca;
34353: douta=16'hb3ca;
34354: douta=16'hb3c9;
34355: douta=16'hb3c9;
34356: douta=16'habc9;
34357: douta=16'habc9;
34358: douta=16'haba9;
34359: douta=16'haba9;
34360: douta=16'habc9;
34361: douta=16'haba9;
34362: douta=16'haba8;
34363: douta=16'haba9;
34364: douta=16'ha389;
34365: douta=16'ha389;
34366: douta=16'ha389;
34367: douta=16'ha389;
34368: douta=16'h8c95;
34369: douta=16'h9d5a;
34370: douta=16'h1861;
34371: douta=16'h2904;
34372: douta=16'h2904;
34373: douta=16'h20e3;
34374: douta=16'h2904;
34375: douta=16'h28e3;
34376: douta=16'h2904;
34377: douta=16'h2904;
34378: douta=16'h20e3;
34379: douta=16'h20e3;
34380: douta=16'h20e3;
34381: douta=16'h28e3;
34382: douta=16'h20a3;
34383: douta=16'h20a3;
34384: douta=16'h20c2;
34385: douta=16'h20c2;
34386: douta=16'h28e3;
34387: douta=16'h28e3;
34388: douta=16'h28e3;
34389: douta=16'h28e3;
34390: douta=16'h3103;
34391: douta=16'h3103;
34392: douta=16'h3103;
34393: douta=16'h3923;
34394: douta=16'h3944;
34395: douta=16'h4164;
34396: douta=16'h4164;
34397: douta=16'h4964;
34398: douta=16'h4a28;
34399: douta=16'h0885;
34400: douta=16'h6204;
34401: douta=16'h59c4;
34402: douta=16'h59e4;
34403: douta=16'h6204;
34404: douta=16'h6204;
34405: douta=16'h6a24;
34406: douta=16'h6a44;
34407: douta=16'h6a44;
34408: douta=16'had10;
34409: douta=16'h7a85;
34410: douta=16'h7a85;
34411: douta=16'h8286;
34412: douta=16'h82a5;
34413: douta=16'h82a6;
34414: douta=16'h82c6;
34415: douta=16'h82c6;
34416: douta=16'h8ac6;
34417: douta=16'h8ae7;
34418: douta=16'h8b07;
34419: douta=16'h9307;
34420: douta=16'h9327;
34421: douta=16'h9b47;
34422: douta=16'h9b47;
34423: douta=16'hb3eb;
34424: douta=16'hde77;
34425: douta=16'hd636;
34426: douta=16'he6b7;
34427: douta=16'hde76;
34428: douta=16'hde98;
34429: douta=16'hb3e8;
34430: douta=16'habc8;
34431: douta=16'hb3c7;
34432: douta=16'hb3e8;
34433: douta=16'hb3e8;
34434: douta=16'hbbe8;
34435: douta=16'hbc08;
34436: douta=16'hbc08;
34437: douta=16'hbc08;
34438: douta=16'hbc08;
34439: douta=16'hc428;
34440: douta=16'hc428;
34441: douta=16'hc448;
34442: douta=16'hc448;
34443: douta=16'hc449;
34444: douta=16'hc448;
34445: douta=16'hc448;
34446: douta=16'hc448;
34447: douta=16'hc448;
34448: douta=16'hc448;
34449: douta=16'hc449;
34450: douta=16'hc468;
34451: douta=16'hc448;
34452: douta=16'hcc69;
34453: douta=16'hcc49;
34454: douta=16'hcc69;
34455: douta=16'hcc69;
34456: douta=16'hcc68;
34457: douta=16'hcc68;
34458: douta=16'hcc68;
34459: douta=16'hcc68;
34460: douta=16'hcc89;
34461: douta=16'hcc69;
34462: douta=16'hcc89;
34463: douta=16'hcc69;
34464: douta=16'hcc69;
34465: douta=16'hcc69;
34466: douta=16'hcc69;
34467: douta=16'hcc89;
34468: douta=16'hcc69;
34469: douta=16'hcc69;
34470: douta=16'hcc89;
34471: douta=16'hcc69;
34472: douta=16'hcc69;
34473: douta=16'hcc8a;
34474: douta=16'hcc89;
34475: douta=16'hcc89;
34476: douta=16'hcc89;
34477: douta=16'hcc89;
34478: douta=16'hcc89;
34479: douta=16'hcc89;
34480: douta=16'hcc89;
34481: douta=16'hcc89;
34482: douta=16'hcc69;
34483: douta=16'hcc89;
34484: douta=16'hcc69;
34485: douta=16'hcc69;
34486: douta=16'hcc69;
34487: douta=16'hcc89;
34488: douta=16'hcc89;
34489: douta=16'hcc89;
34490: douta=16'hb595;
34491: douta=16'he675;
34492: douta=16'hcc69;
34493: douta=16'hcc6a;
34494: douta=16'hcc69;
34495: douta=16'hcc69;
34496: douta=16'hcc6a;
34497: douta=16'hcc6a;
34498: douta=16'hcc6a;
34499: douta=16'hcc69;
34500: douta=16'hcc69;
34501: douta=16'hcc6a;
34502: douta=16'hcc49;
34503: douta=16'hcc69;
34504: douta=16'hcc49;
34505: douta=16'hc449;
34506: douta=16'hcc49;
34507: douta=16'hcc49;
34508: douta=16'hcc49;
34509: douta=16'hc449;
34510: douta=16'hcc49;
34511: douta=16'hc449;
34512: douta=16'hc449;
34513: douta=16'hc449;
34514: douta=16'hc449;
34515: douta=16'hc469;
34516: douta=16'hc449;
34517: douta=16'hc449;
34518: douta=16'hc44a;
34519: douta=16'hc429;
34520: douta=16'hc429;
34521: douta=16'hc44a;
34522: douta=16'hbc29;
34523: douta=16'hc429;
34524: douta=16'hc429;
34525: douta=16'hc42a;
34526: douta=16'hc40a;
34527: douta=16'hbc09;
34528: douta=16'hbc2a;
34529: douta=16'hbc2a;
34530: douta=16'hbc09;
34531: douta=16'hbc09;
34532: douta=16'hbc09;
34533: douta=16'hbc09;
34534: douta=16'hbc09;
34535: douta=16'hbc09;
34536: douta=16'hbc09;
34537: douta=16'hbc09;
34538: douta=16'hb3e9;
34539: douta=16'hb3e9;
34540: douta=16'hb3e9;
34541: douta=16'hb3e9;
34542: douta=16'hb3e9;
34543: douta=16'hb3e9;
34544: douta=16'hb3c9;
34545: douta=16'hb3e9;
34546: douta=16'hb3ca;
34547: douta=16'habc9;
34548: douta=16'habc9;
34549: douta=16'hb3ca;
34550: douta=16'habc9;
34551: douta=16'habc9;
34552: douta=16'haba9;
34553: douta=16'habc9;
34554: douta=16'haba9;
34555: douta=16'haba9;
34556: douta=16'haba9;
34557: douta=16'haba9;
34558: douta=16'ha389;
34559: douta=16'ha389;
34560: douta=16'h8c96;
34561: douta=16'h84b7;
34562: douta=16'h20a2;
34563: douta=16'h2904;
34564: douta=16'h2904;
34565: douta=16'h28e3;
34566: douta=16'h28e3;
34567: douta=16'h2904;
34568: douta=16'h2904;
34569: douta=16'h2904;
34570: douta=16'h20e4;
34571: douta=16'h20e3;
34572: douta=16'h20e3;
34573: douta=16'h2904;
34574: douta=16'h20a2;
34575: douta=16'h20a3;
34576: douta=16'h20c2;
34577: douta=16'h20c2;
34578: douta=16'h28c3;
34579: douta=16'h28e3;
34580: douta=16'h28e3;
34581: douta=16'h28e3;
34582: douta=16'h3103;
34583: douta=16'h3103;
34584: douta=16'h3903;
34585: douta=16'h3944;
34586: douta=16'h3944;
34587: douta=16'h4164;
34588: douta=16'h4964;
34589: douta=16'h4985;
34590: douta=16'h4a29;
34591: douta=16'h0885;
34592: douta=16'h61c4;
34593: douta=16'h59e4;
34594: douta=16'h61e4;
34595: douta=16'h6204;
34596: douta=16'h6205;
34597: douta=16'h6a44;
34598: douta=16'h6a44;
34599: douta=16'h7245;
34600: douta=16'haccf;
34601: douta=16'h7244;
34602: douta=16'h7a85;
34603: douta=16'h7a85;
34604: douta=16'h82a5;
34605: douta=16'h82c6;
34606: douta=16'h82c6;
34607: douta=16'h82c6;
34608: douta=16'h8ae7;
34609: douta=16'h8ae7;
34610: douta=16'h8b07;
34611: douta=16'h8b07;
34612: douta=16'h9327;
34613: douta=16'h9b47;
34614: douta=16'h9b47;
34615: douta=16'hc48f;
34616: douta=16'heef9;
34617: douta=16'hdeb8;
34618: douta=16'he6d9;
34619: douta=16'hef3b;
34620: douta=16'hce78;
34621: douta=16'hb3e8;
34622: douta=16'hb3c8;
34623: douta=16'hb3c7;
34624: douta=16'hb3e8;
34625: douta=16'hb3e8;
34626: douta=16'hbc08;
34627: douta=16'hbc08;
34628: douta=16'hbc08;
34629: douta=16'hbc08;
34630: douta=16'hbc08;
34631: douta=16'hc428;
34632: douta=16'hc428;
34633: douta=16'hc428;
34634: douta=16'hc428;
34635: douta=16'hc449;
34636: douta=16'hc449;
34637: douta=16'hc448;
34638: douta=16'hc448;
34639: douta=16'hc448;
34640: douta=16'hc448;
34641: douta=16'hc448;
34642: douta=16'hcc69;
34643: douta=16'hc468;
34644: douta=16'hcc69;
34645: douta=16'hcc49;
34646: douta=16'hcc69;
34647: douta=16'hcc69;
34648: douta=16'hcc69;
34649: douta=16'hcc69;
34650: douta=16'hcc69;
34651: douta=16'hcc69;
34652: douta=16'hcc89;
34653: douta=16'hcc69;
34654: douta=16'hcc89;
34655: douta=16'hcc89;
34656: douta=16'hcc69;
34657: douta=16'hcc89;
34658: douta=16'hcc69;
34659: douta=16'hcc69;
34660: douta=16'hcc69;
34661: douta=16'hcc89;
34662: douta=16'hcc69;
34663: douta=16'hcc89;
34664: douta=16'hcc69;
34665: douta=16'hcc89;
34666: douta=16'hcc89;
34667: douta=16'hcc89;
34668: douta=16'hcc69;
34669: douta=16'hcc89;
34670: douta=16'hcc89;
34671: douta=16'hcc89;
34672: douta=16'hcc89;
34673: douta=16'hcc69;
34674: douta=16'hcc69;
34675: douta=16'hcc89;
34676: douta=16'hcc69;
34677: douta=16'hcc89;
34678: douta=16'hcc89;
34679: douta=16'hcc89;
34680: douta=16'hcc89;
34681: douta=16'hcc69;
34682: douta=16'hb5b5;
34683: douta=16'he675;
34684: douta=16'hcc6a;
34685: douta=16'hcc6a;
34686: douta=16'hcc69;
34687: douta=16'hcc69;
34688: douta=16'hcc6a;
34689: douta=16'hcc69;
34690: douta=16'hcc69;
34691: douta=16'hcc49;
34692: douta=16'hcc69;
34693: douta=16'hcc69;
34694: douta=16'hcc69;
34695: douta=16'hcc69;
34696: douta=16'hcc69;
34697: douta=16'hcc69;
34698: douta=16'hcc69;
34699: douta=16'hcc69;
34700: douta=16'hc449;
34701: douta=16'hcc69;
34702: douta=16'hc449;
34703: douta=16'hc449;
34704: douta=16'hc449;
34705: douta=16'hc449;
34706: douta=16'hc449;
34707: douta=16'hc449;
34708: douta=16'hc469;
34709: douta=16'hc449;
34710: douta=16'hc44a;
34711: douta=16'hc44a;
34712: douta=16'hc429;
34713: douta=16'hc429;
34714: douta=16'hc429;
34715: douta=16'hc429;
34716: douta=16'hbc29;
34717: douta=16'hbc09;
34718: douta=16'hc40a;
34719: douta=16'hc40a;
34720: douta=16'hbc09;
34721: douta=16'hbc09;
34722: douta=16'hbc2a;
34723: douta=16'hbc09;
34724: douta=16'hbc09;
34725: douta=16'hbc09;
34726: douta=16'hbc09;
34727: douta=16'hbc09;
34728: douta=16'hbc09;
34729: douta=16'hbc09;
34730: douta=16'hbbe9;
34731: douta=16'hbbe9;
34732: douta=16'hbbe9;
34733: douta=16'hb3e9;
34734: douta=16'hbbe9;
34735: douta=16'hb3e9;
34736: douta=16'hb3c9;
34737: douta=16'hb3e9;
34738: douta=16'hb3ca;
34739: douta=16'hb3c9;
34740: douta=16'habc9;
34741: douta=16'hb3ca;
34742: douta=16'habc9;
34743: douta=16'habc9;
34744: douta=16'haba9;
34745: douta=16'haba9;
34746: douta=16'haba9;
34747: douta=16'hab89;
34748: douta=16'haba9;
34749: douta=16'ha389;
34750: douta=16'ha389;
34751: douta=16'ha369;
34752: douta=16'h8496;
34753: douta=16'h3186;
34754: douta=16'h2924;
34755: douta=16'h3124;
34756: douta=16'h2904;
34757: douta=16'h2904;
34758: douta=16'h2904;
34759: douta=16'h2924;
34760: douta=16'h2904;
34761: douta=16'h2904;
34762: douta=16'h20e4;
34763: douta=16'h20e3;
34764: douta=16'h2103;
34765: douta=16'h2904;
34766: douta=16'h20c2;
34767: douta=16'h20e3;
34768: douta=16'h28e3;
34769: douta=16'h28e3;
34770: douta=16'h28e3;
34771: douta=16'h28e3;
34772: douta=16'h28e3;
34773: douta=16'h2903;
34774: douta=16'h3103;
34775: douta=16'h3103;
34776: douta=16'h3103;
34777: douta=16'h4144;
34778: douta=16'h4144;
34779: douta=16'h4964;
34780: douta=16'h4964;
34781: douta=16'h49e7;
34782: douta=16'h5acd;
34783: douta=16'h20e5;
34784: douta=16'h59e4;
34785: douta=16'h59c4;
34786: douta=16'h61e4;
34787: douta=16'h6204;
34788: douta=16'h6a25;
34789: douta=16'h7245;
34790: douta=16'h7245;
34791: douta=16'h7244;
34792: douta=16'h938a;
34793: douta=16'h7a24;
34794: douta=16'h7a85;
34795: douta=16'h8285;
34796: douta=16'h82a5;
34797: douta=16'h82c6;
34798: douta=16'h82c6;
34799: douta=16'h82c6;
34800: douta=16'h8ae7;
34801: douta=16'h8ae7;
34802: douta=16'h8b07;
34803: douta=16'h9307;
34804: douta=16'h9327;
34805: douta=16'h9b47;
34806: douta=16'h9b47;
34807: douta=16'h9b46;
34808: douta=16'h9b05;
34809: douta=16'h9b46;
34810: douta=16'ha367;
34811: douta=16'ha388;
34812: douta=16'ha387;
34813: douta=16'hb3a8;
34814: douta=16'hb3c8;
34815: douta=16'hb3c8;
34816: douta=16'hb3e8;
34817: douta=16'hb3e8;
34818: douta=16'hb3e8;
34819: douta=16'hbc08;
34820: douta=16'hbc08;
34821: douta=16'hbc29;
34822: douta=16'hbc28;
34823: douta=16'hbc28;
34824: douta=16'hc428;
34825: douta=16'hc449;
34826: douta=16'hc449;
34827: douta=16'hc449;
34828: douta=16'hc449;
34829: douta=16'hc449;
34830: douta=16'hc448;
34831: douta=16'hc448;
34832: douta=16'hc448;
34833: douta=16'hc468;
34834: douta=16'hcc69;
34835: douta=16'hc468;
34836: douta=16'hcc69;
34837: douta=16'hcc69;
34838: douta=16'hcc69;
34839: douta=16'hcc69;
34840: douta=16'hcc69;
34841: douta=16'hcc69;
34842: douta=16'hcc69;
34843: douta=16'hcc69;
34844: douta=16'hcc69;
34845: douta=16'hcc89;
34846: douta=16'hcc89;
34847: douta=16'hcc89;
34848: douta=16'hcc89;
34849: douta=16'hcc89;
34850: douta=16'hcc89;
34851: douta=16'hcc89;
34852: douta=16'hcc69;
34853: douta=16'hcc69;
34854: douta=16'hcc69;
34855: douta=16'hcc69;
34856: douta=16'hcc69;
34857: douta=16'hcc89;
34858: douta=16'hcc89;
34859: douta=16'hcc89;
34860: douta=16'hcc89;
34861: douta=16'hcc89;
34862: douta=16'hcc89;
34863: douta=16'hcc69;
34864: douta=16'hcc89;
34865: douta=16'hcc69;
34866: douta=16'hcc69;
34867: douta=16'hcc89;
34868: douta=16'hcc69;
34869: douta=16'hcc89;
34870: douta=16'hcc89;
34871: douta=16'hcc89;
34872: douta=16'hc489;
34873: douta=16'hcc68;
34874: douta=16'hb5d5;
34875: douta=16'he655;
34876: douta=16'hcc6a;
34877: douta=16'hcc6a;
34878: douta=16'hcc89;
34879: douta=16'hcc89;
34880: douta=16'hcc69;
34881: douta=16'hcc6a;
34882: douta=16'hcc69;
34883: douta=16'hcc49;
34884: douta=16'hcc49;
34885: douta=16'hcc69;
34886: douta=16'hcc69;
34887: douta=16'hcc69;
34888: douta=16'hcc69;
34889: douta=16'hcc49;
34890: douta=16'hc44a;
34891: douta=16'hcc6a;
34892: douta=16'hc44a;
34893: douta=16'hc449;
34894: douta=16'hc449;
34895: douta=16'hc469;
34896: douta=16'hc449;
34897: douta=16'hc449;
34898: douta=16'hc449;
34899: douta=16'hc449;
34900: douta=16'hc449;
34901: douta=16'hc429;
34902: douta=16'hc44a;
34903: douta=16'hc429;
34904: douta=16'hc44a;
34905: douta=16'hc429;
34906: douta=16'hc429;
34907: douta=16'hc429;
34908: douta=16'hbc29;
34909: douta=16'hc40a;
34910: douta=16'hbc2a;
34911: douta=16'hbc09;
34912: douta=16'hbc2a;
34913: douta=16'hbc2a;
34914: douta=16'hbc2a;
34915: douta=16'hbc2a;
34916: douta=16'hbc09;
34917: douta=16'hbc09;
34918: douta=16'hbc09;
34919: douta=16'hbc09;
34920: douta=16'hbc09;
34921: douta=16'hbc09;
34922: douta=16'hbbe9;
34923: douta=16'hb3e9;
34924: douta=16'hbbe9;
34925: douta=16'hb3e9;
34926: douta=16'hb3e9;
34927: douta=16'hb3e9;
34928: douta=16'hb3e9;
34929: douta=16'hb3c9;
34930: douta=16'hb3c9;
34931: douta=16'hb3ca;
34932: douta=16'habc9;
34933: douta=16'hb3c9;
34934: douta=16'habc9;
34935: douta=16'haba9;
34936: douta=16'haba9;
34937: douta=16'haba9;
34938: douta=16'haba9;
34939: douta=16'haba9;
34940: douta=16'ha389;
34941: douta=16'habaa;
34942: douta=16'ha389;
34943: douta=16'ha389;
34944: douta=16'h8cb7;
34945: douta=16'h1861;
34946: douta=16'h2904;
34947: douta=16'h2924;
34948: douta=16'h3124;
34949: douta=16'h2904;
34950: douta=16'h2904;
34951: douta=16'h2924;
34952: douta=16'h2904;
34953: douta=16'h2904;
34954: douta=16'h20e3;
34955: douta=16'h20e3;
34956: douta=16'h2103;
34957: douta=16'h28e3;
34958: douta=16'h20c2;
34959: douta=16'h20e3;
34960: douta=16'h20e3;
34961: douta=16'h28e3;
34962: douta=16'h28e3;
34963: douta=16'h28e3;
34964: douta=16'h2903;
34965: douta=16'h2903;
34966: douta=16'h3124;
34967: douta=16'h3903;
34968: douta=16'h3923;
34969: douta=16'h3923;
34970: douta=16'h4144;
34971: douta=16'h4964;
34972: douta=16'h4984;
34973: douta=16'h4a28;
34974: douta=16'h528b;
34975: douta=16'h3124;
34976: douta=16'h59c4;
34977: douta=16'h61e4;
34978: douta=16'h6a05;
34979: douta=16'h6204;
34980: douta=16'h6a24;
34981: douta=16'h7244;
34982: douta=16'h7245;
34983: douta=16'h7224;
34984: douta=16'h7aa5;
34985: douta=16'h7244;
34986: douta=16'h82a5;
34987: douta=16'h8285;
34988: douta=16'h82a6;
34989: douta=16'h8ac6;
34990: douta=16'h8ac6;
34991: douta=16'h8ae6;
34992: douta=16'h9307;
34993: douta=16'h8ae7;
34994: douta=16'h9307;
34995: douta=16'h9307;
34996: douta=16'h9327;
34997: douta=16'h9b47;
34998: douta=16'h9b47;
34999: douta=16'ha368;
35000: douta=16'ha368;
35001: douta=16'h9b67;
35002: douta=16'ha368;
35003: douta=16'ha388;
35004: douta=16'ha388;
35005: douta=16'haba8;
35006: douta=16'hb3c8;
35007: douta=16'hb3c8;
35008: douta=16'hb3e8;
35009: douta=16'hb3e8;
35010: douta=16'hbbe8;
35011: douta=16'hbc08;
35012: douta=16'hbc08;
35013: douta=16'hbc29;
35014: douta=16'hbc29;
35015: douta=16'hbc28;
35016: douta=16'hbc29;
35017: douta=16'hc449;
35018: douta=16'hc449;
35019: douta=16'hc449;
35020: douta=16'hc449;
35021: douta=16'hc449;
35022: douta=16'hc449;
35023: douta=16'hc448;
35024: douta=16'hc468;
35025: douta=16'hcc49;
35026: douta=16'hcc69;
35027: douta=16'hcc69;
35028: douta=16'hcc69;
35029: douta=16'hcc69;
35030: douta=16'hcc69;
35031: douta=16'hcc69;
35032: douta=16'hcc69;
35033: douta=16'hcc69;
35034: douta=16'hcc69;
35035: douta=16'hcc69;
35036: douta=16'hcc89;
35037: douta=16'hcc69;
35038: douta=16'hcc89;
35039: douta=16'hcc69;
35040: douta=16'hcc89;
35041: douta=16'hcc69;
35042: douta=16'hcc89;
35043: douta=16'hcc69;
35044: douta=16'hcc89;
35045: douta=16'hcc69;
35046: douta=16'hcc69;
35047: douta=16'hcc89;
35048: douta=16'hcc89;
35049: douta=16'hcc89;
35050: douta=16'hcc89;
35051: douta=16'hcc69;
35052: douta=16'hcc89;
35053: douta=16'hcc89;
35054: douta=16'hcc89;
35055: douta=16'hcc89;
35056: douta=16'hcc69;
35057: douta=16'hcc69;
35058: douta=16'hcc89;
35059: douta=16'hcc69;
35060: douta=16'hcc69;
35061: douta=16'hcc69;
35062: douta=16'hcc89;
35063: douta=16'hc489;
35064: douta=16'hcc6a;
35065: douta=16'hcc69;
35066: douta=16'hb5d5;
35067: douta=16'he675;
35068: douta=16'hc469;
35069: douta=16'hcc69;
35070: douta=16'hcc69;
35071: douta=16'hcc69;
35072: douta=16'hcc69;
35073: douta=16'hcc6a;
35074: douta=16'hcc6a;
35075: douta=16'hcc69;
35076: douta=16'hcc49;
35077: douta=16'hcc6a;
35078: douta=16'hcc6a;
35079: douta=16'hcc69;
35080: douta=16'hcc49;
35081: douta=16'hcc6a;
35082: douta=16'hcc6a;
35083: douta=16'hc449;
35084: douta=16'hc449;
35085: douta=16'hc46a;
35086: douta=16'hc469;
35087: douta=16'hc449;
35088: douta=16'hc469;
35089: douta=16'hc449;
35090: douta=16'hc449;
35091: douta=16'hc44a;
35092: douta=16'hc44a;
35093: douta=16'hc44a;
35094: douta=16'hc44a;
35095: douta=16'hc429;
35096: douta=16'hc42a;
35097: douta=16'hc42a;
35098: douta=16'hbc2a;
35099: douta=16'hbc29;
35100: douta=16'hbc09;
35101: douta=16'hbc0a;
35102: douta=16'hbc0a;
35103: douta=16'hbc2a;
35104: douta=16'hbc09;
35105: douta=16'hbc2a;
35106: douta=16'hbc09;
35107: douta=16'hbc09;
35108: douta=16'hbc09;
35109: douta=16'hbc09;
35110: douta=16'hbc09;
35111: douta=16'hbc09;
35112: douta=16'hbc09;
35113: douta=16'hbc09;
35114: douta=16'hbc09;
35115: douta=16'hbbe9;
35116: douta=16'hb3e9;
35117: douta=16'hb3e9;
35118: douta=16'hb3e9;
35119: douta=16'hb3e9;
35120: douta=16'hb3c9;
35121: douta=16'hb3c9;
35122: douta=16'hb3ca;
35123: douta=16'haba9;
35124: douta=16'hb3ca;
35125: douta=16'habc9;
35126: douta=16'habc9;
35127: douta=16'habc9;
35128: douta=16'haba9;
35129: douta=16'haba9;
35130: douta=16'haba9;
35131: douta=16'haba9;
35132: douta=16'ha389;
35133: douta=16'hab89;
35134: douta=16'hab8a;
35135: douta=16'ha389;
35136: douta=16'h9519;
35137: douta=16'h28e3;
35138: douta=16'h2904;
35139: douta=16'h2924;
35140: douta=16'h2904;
35141: douta=16'h3124;
35142: douta=16'h2904;
35143: douta=16'h2904;
35144: douta=16'h2904;
35145: douta=16'h28e4;
35146: douta=16'h20e3;
35147: douta=16'h2103;
35148: douta=16'h20e3;
35149: douta=16'h20e3;
35150: douta=16'h20c3;
35151: douta=16'h20c3;
35152: douta=16'h28e3;
35153: douta=16'h28e3;
35154: douta=16'h28e3;
35155: douta=16'h2903;
35156: douta=16'h3123;
35157: douta=16'h3103;
35158: douta=16'h3103;
35159: douta=16'h3903;
35160: douta=16'h3923;
35161: douta=16'h3944;
35162: douta=16'h4144;
35163: douta=16'h4964;
35164: douta=16'h51a5;
35165: douta=16'h4a49;
35166: douta=16'h4a2a;
35167: douta=16'h3945;
35168: douta=16'h59c4;
35169: douta=16'h59e4;
35170: douta=16'h6a05;
35171: douta=16'h6a05;
35172: douta=16'h6a24;
35173: douta=16'h6a24;
35174: douta=16'h7245;
35175: douta=16'h7224;
35176: douta=16'h7244;
35177: douta=16'h7a64;
35178: douta=16'h7a85;
35179: douta=16'h82a6;
35180: douta=16'h82a6;
35181: douta=16'h82c6;
35182: douta=16'h82a6;
35183: douta=16'h82c6;
35184: douta=16'h8ae7;
35185: douta=16'h8ae7;
35186: douta=16'h8b07;
35187: douta=16'h9307;
35188: douta=16'h9327;
35189: douta=16'h9327;
35190: douta=16'h9b47;
35191: douta=16'ha368;
35192: douta=16'h9b67;
35193: douta=16'ha368;
35194: douta=16'ha388;
35195: douta=16'hab88;
35196: douta=16'ha388;
35197: douta=16'haba8;
35198: douta=16'hb3c8;
35199: douta=16'hb3e8;
35200: douta=16'hb3e8;
35201: douta=16'hbbe8;
35202: douta=16'hb3e8;
35203: douta=16'hbc08;
35204: douta=16'hbc08;
35205: douta=16'hbc08;
35206: douta=16'hbc29;
35207: douta=16'hc428;
35208: douta=16'hc429;
35209: douta=16'hc449;
35210: douta=16'hc449;
35211: douta=16'hc449;
35212: douta=16'hc449;
35213: douta=16'hc449;
35214: douta=16'hc449;
35215: douta=16'hc468;
35216: douta=16'hc448;
35217: douta=16'hcc49;
35218: douta=16'hcc69;
35219: douta=16'hcc69;
35220: douta=16'hcc69;
35221: douta=16'hcc6a;
35222: douta=16'hcc69;
35223: douta=16'hcc69;
35224: douta=16'hcc69;
35225: douta=16'hcc69;
35226: douta=16'hcc69;
35227: douta=16'hcc69;
35228: douta=16'hcc89;
35229: douta=16'hcc89;
35230: douta=16'hcc8a;
35231: douta=16'hcc6a;
35232: douta=16'hcc89;
35233: douta=16'hcc89;
35234: douta=16'hcc89;
35235: douta=16'hcc89;
35236: douta=16'hcc69;
35237: douta=16'hcc69;
35238: douta=16'hcc89;
35239: douta=16'hcc89;
35240: douta=16'hcc89;
35241: douta=16'hcc89;
35242: douta=16'hcc89;
35243: douta=16'hcc69;
35244: douta=16'hcc6a;
35245: douta=16'hcc89;
35246: douta=16'hcc69;
35247: douta=16'hcc89;
35248: douta=16'hcc69;
35249: douta=16'hcc69;
35250: douta=16'hcc69;
35251: douta=16'hcc69;
35252: douta=16'hcc89;
35253: douta=16'hcc89;
35254: douta=16'hcc69;
35255: douta=16'hc489;
35256: douta=16'hcc6a;
35257: douta=16'hcc69;
35258: douta=16'hb5b5;
35259: douta=16'he655;
35260: douta=16'hc469;
35261: douta=16'hc469;
35262: douta=16'hcc69;
35263: douta=16'hcc69;
35264: douta=16'hcc69;
35265: douta=16'hcc8a;
35266: douta=16'hcc6a;
35267: douta=16'hcc49;
35268: douta=16'hcc69;
35269: douta=16'hcc6a;
35270: douta=16'hcc6a;
35271: douta=16'hcc49;
35272: douta=16'hcc69;
35273: douta=16'hc44a;
35274: douta=16'hc44a;
35275: douta=16'hc44a;
35276: douta=16'hc46a;
35277: douta=16'hc469;
35278: douta=16'hc449;
35279: douta=16'hc46a;
35280: douta=16'hc469;
35281: douta=16'hc449;
35282: douta=16'hc449;
35283: douta=16'hc44a;
35284: douta=16'hc44a;
35285: douta=16'hc44a;
35286: douta=16'hc429;
35287: douta=16'hc429;
35288: douta=16'hc42a;
35289: douta=16'hc42a;
35290: douta=16'hc42a;
35291: douta=16'hbc29;
35292: douta=16'hbc29;
35293: douta=16'hbc09;
35294: douta=16'hbc09;
35295: douta=16'hbc2a;
35296: douta=16'hbc2a;
35297: douta=16'hbc09;
35298: douta=16'hbc09;
35299: douta=16'hbc09;
35300: douta=16'hbc2a;
35301: douta=16'hbc0a;
35302: douta=16'hbc09;
35303: douta=16'hbc09;
35304: douta=16'hbc09;
35305: douta=16'hbbe9;
35306: douta=16'hbbe9;
35307: douta=16'hbbe9;
35308: douta=16'hb3e9;
35309: douta=16'hb3e9;
35310: douta=16'hb3e9;
35311: douta=16'hb3c9;
35312: douta=16'hb3e9;
35313: douta=16'hb3c9;
35314: douta=16'hb3ca;
35315: douta=16'habc9;
35316: douta=16'hb3c9;
35317: douta=16'habc9;
35318: douta=16'habc9;
35319: douta=16'haba9;
35320: douta=16'haba9;
35321: douta=16'haba9;
35322: douta=16'hab89;
35323: douta=16'hab89;
35324: douta=16'ha389;
35325: douta=16'hab89;
35326: douta=16'ha38a;
35327: douta=16'ha389;
35328: douta=16'h7c55;
35329: douta=16'h3145;
35330: douta=16'h2925;
35331: douta=16'h3124;
35332: douta=16'h3124;
35333: douta=16'h3124;
35334: douta=16'h2904;
35335: douta=16'h2904;
35336: douta=16'h2904;
35337: douta=16'h28e4;
35338: douta=16'h20e3;
35339: douta=16'h28e3;
35340: douta=16'h2904;
35341: douta=16'h20a2;
35342: douta=16'h20e3;
35343: douta=16'h20e3;
35344: douta=16'h28e3;
35345: douta=16'h2903;
35346: douta=16'h2903;
35347: douta=16'h2903;
35348: douta=16'h28e3;
35349: douta=16'h3103;
35350: douta=16'h3123;
35351: douta=16'h3923;
35352: douta=16'h3923;
35353: douta=16'h3943;
35354: douta=16'h4144;
35355: douta=16'h4964;
35356: douta=16'h4984;
35357: douta=16'h5a8b;
35358: douta=16'h3987;
35359: douta=16'h59c5;
35360: douta=16'h59e4;
35361: douta=16'h59c4;
35362: douta=16'h6204;
35363: douta=16'h6204;
35364: douta=16'h6a25;
35365: douta=16'h7245;
35366: douta=16'h7225;
35367: douta=16'h7224;
35368: douta=16'h7224;
35369: douta=16'h7a84;
35370: douta=16'h7a85;
35371: douta=16'h82a6;
35372: douta=16'h82c6;
35373: douta=16'h82c6;
35374: douta=16'h82c6;
35375: douta=16'h8ae7;
35376: douta=16'h8b07;
35377: douta=16'h9307;
35378: douta=16'h9307;
35379: douta=16'h9327;
35380: douta=16'h9328;
35381: douta=16'h9b47;
35382: douta=16'h9b68;
35383: douta=16'h9b67;
35384: douta=16'h9b67;
35385: douta=16'ha368;
35386: douta=16'ha388;
35387: douta=16'ha388;
35388: douta=16'ha388;
35389: douta=16'haba8;
35390: douta=16'hb3c8;
35391: douta=16'hb3e7;
35392: douta=16'hbc08;
35393: douta=16'hbbe8;
35394: douta=16'hbc09;
35395: douta=16'hbc09;
35396: douta=16'hbc08;
35397: douta=16'hbc29;
35398: douta=16'hbc29;
35399: douta=16'hc429;
35400: douta=16'hc449;
35401: douta=16'hc449;
35402: douta=16'hc449;
35403: douta=16'hc449;
35404: douta=16'hc429;
35405: douta=16'hc449;
35406: douta=16'hc428;
35407: douta=16'hcc49;
35408: douta=16'hc449;
35409: douta=16'hc469;
35410: douta=16'hc449;
35411: douta=16'hc449;
35412: douta=16'hc469;
35413: douta=16'hcc69;
35414: douta=16'hcc69;
35415: douta=16'hcc69;
35416: douta=16'hcc49;
35417: douta=16'hcc69;
35418: douta=16'hcc69;
35419: douta=16'hcc6a;
35420: douta=16'hcc6a;
35421: douta=16'hcc6a;
35422: douta=16'hcc6a;
35423: douta=16'hcc69;
35424: douta=16'hcc8a;
35425: douta=16'hcc89;
35426: douta=16'hcc69;
35427: douta=16'hcc69;
35428: douta=16'hcc69;
35429: douta=16'hcc89;
35430: douta=16'hcc69;
35431: douta=16'hcc69;
35432: douta=16'hcc89;
35433: douta=16'hcc69;
35434: douta=16'hcc6a;
35435: douta=16'hcc69;
35436: douta=16'hcc6a;
35437: douta=16'hcc69;
35438: douta=16'hcc89;
35439: douta=16'hcc89;
35440: douta=16'hcc89;
35441: douta=16'hcc6a;
35442: douta=16'hcc6a;
35443: douta=16'hcc89;
35444: douta=16'hcc89;
35445: douta=16'hcc6a;
35446: douta=16'hcc8a;
35447: douta=16'hc469;
35448: douta=16'hcc6a;
35449: douta=16'hcc69;
35450: douta=16'hb5b5;
35451: douta=16'he655;
35452: douta=16'hc469;
35453: douta=16'hc469;
35454: douta=16'hcc6a;
35455: douta=16'hcc6a;
35456: douta=16'hcc69;
35457: douta=16'hcc69;
35458: douta=16'hcc6a;
35459: douta=16'hcc49;
35460: douta=16'hc449;
35461: douta=16'hcc6a;
35462: douta=16'hc44a;
35463: douta=16'hcc69;
35464: douta=16'hc449;
35465: douta=16'hcc6a;
35466: douta=16'hc44a;
35467: douta=16'hc469;
35468: douta=16'hc46a;
35469: douta=16'hc449;
35470: douta=16'hc449;
35471: douta=16'hc449;
35472: douta=16'hc449;
35473: douta=16'hc449;
35474: douta=16'hc429;
35475: douta=16'hc429;
35476: douta=16'hc429;
35477: douta=16'hc44a;
35478: douta=16'hc44a;
35479: douta=16'hc44a;
35480: douta=16'hc42a;
35481: douta=16'hc42a;
35482: douta=16'hbc2a;
35483: douta=16'hc42a;
35484: douta=16'hbc09;
35485: douta=16'hbc09;
35486: douta=16'hbc09;
35487: douta=16'hbc2a;
35488: douta=16'hbc2a;
35489: douta=16'hbc09;
35490: douta=16'hbc09;
35491: douta=16'hbc09;
35492: douta=16'hbc0a;
35493: douta=16'hbc09;
35494: douta=16'hbc09;
35495: douta=16'hbbe9;
35496: douta=16'hbc09;
35497: douta=16'hbc09;
35498: douta=16'hbbe9;
35499: douta=16'hb3c9;
35500: douta=16'hb3e9;
35501: douta=16'hb3e9;
35502: douta=16'hb3e9;
35503: douta=16'hb3c9;
35504: douta=16'hb3ea;
35505: douta=16'hb3ca;
35506: douta=16'habc9;
35507: douta=16'habc9;
35508: douta=16'habc9;
35509: douta=16'habc9;
35510: douta=16'habca;
35511: douta=16'haba9;
35512: douta=16'haba9;
35513: douta=16'haba9;
35514: douta=16'haba9;
35515: douta=16'haba9;
35516: douta=16'ha389;
35517: douta=16'ha389;
35518: douta=16'ha369;
35519: douta=16'ha389;
35520: douta=16'h4229;
35521: douta=16'h3145;
35522: douta=16'h3125;
35523: douta=16'h3124;
35524: douta=16'h3124;
35525: douta=16'h2924;
35526: douta=16'h2904;
35527: douta=16'h2904;
35528: douta=16'h2904;
35529: douta=16'h28e4;
35530: douta=16'h2104;
35531: douta=16'h2103;
35532: douta=16'h2904;
35533: douta=16'h20a2;
35534: douta=16'h20e3;
35535: douta=16'h28e3;
35536: douta=16'h28e3;
35537: douta=16'h2903;
35538: douta=16'h28e3;
35539: douta=16'h28e3;
35540: douta=16'h28e3;
35541: douta=16'h3103;
35542: douta=16'h3123;
35543: douta=16'h3923;
35544: douta=16'h3923;
35545: douta=16'h4144;
35546: douta=16'h4143;
35547: douta=16'h4984;
35548: douta=16'h49a5;
35549: douta=16'h4a4a;
35550: douta=16'h2105;
35551: douta=16'h61e4;
35552: douta=16'h59e4;
35553: douta=16'h59e4;
35554: douta=16'h6225;
35555: douta=16'h6a25;
35556: douta=16'h6a45;
35557: douta=16'h6a25;
35558: douta=16'h7224;
35559: douta=16'h72a8;
35560: douta=16'h7a44;
35561: douta=16'h7a85;
35562: douta=16'h82a5;
35563: douta=16'h82a6;
35564: douta=16'h82c6;
35565: douta=16'h82c6;
35566: douta=16'h8ac7;
35567: douta=16'h8ae7;
35568: douta=16'h8b07;
35569: douta=16'h9307;
35570: douta=16'h9327;
35571: douta=16'h9327;
35572: douta=16'h9327;
35573: douta=16'h9b47;
35574: douta=16'h9b47;
35575: douta=16'h9b68;
35576: douta=16'h9b68;
35577: douta=16'ha368;
35578: douta=16'ha388;
35579: douta=16'ha387;
35580: douta=16'ha388;
35581: douta=16'haba8;
35582: douta=16'hb3c8;
35583: douta=16'hb3e8;
35584: douta=16'hb408;
35585: douta=16'hb408;
35586: douta=16'hb3e8;
35587: douta=16'hbc09;
35588: douta=16'hbc09;
35589: douta=16'hbc09;
35590: douta=16'hbc29;
35591: douta=16'hbc29;
35592: douta=16'hbc49;
35593: douta=16'hc449;
35594: douta=16'hc449;
35595: douta=16'hc449;
35596: douta=16'hc449;
35597: douta=16'hc449;
35598: douta=16'hc469;
35599: douta=16'hc449;
35600: douta=16'hc469;
35601: douta=16'hc46a;
35602: douta=16'hc469;
35603: douta=16'hcc8a;
35604: douta=16'hcc6a;
35605: douta=16'hc469;
35606: douta=16'hcc6a;
35607: douta=16'hcc6a;
35608: douta=16'hcc6a;
35609: douta=16'hcc69;
35610: douta=16'hcc6a;
35611: douta=16'hcc8a;
35612: douta=16'hcc69;
35613: douta=16'hcc6a;
35614: douta=16'hcc6a;
35615: douta=16'hcc6a;
35616: douta=16'hcc8a;
35617: douta=16'hcc89;
35618: douta=16'hcc69;
35619: douta=16'hcc69;
35620: douta=16'hcc69;
35621: douta=16'hcc89;
35622: douta=16'hcc69;
35623: douta=16'hcc69;
35624: douta=16'hcc69;
35625: douta=16'hcc69;
35626: douta=16'hcc69;
35627: douta=16'hcc69;
35628: douta=16'hcc69;
35629: douta=16'hcc69;
35630: douta=16'hcc69;
35631: douta=16'hc489;
35632: douta=16'hcc6a;
35633: douta=16'hcc6a;
35634: douta=16'hcc69;
35635: douta=16'hcc6a;
35636: douta=16'hcc69;
35637: douta=16'hcc6a;
35638: douta=16'hcc8a;
35639: douta=16'hcc6a;
35640: douta=16'hcc6a;
35641: douta=16'hcc6a;
35642: douta=16'hb5d5;
35643: douta=16'he654;
35644: douta=16'hcc6a;
35645: douta=16'hcc6a;
35646: douta=16'hc469;
35647: douta=16'hcc69;
35648: douta=16'hcc69;
35649: douta=16'hcc69;
35650: douta=16'hcc69;
35651: douta=16'hcc69;
35652: douta=16'hcc49;
35653: douta=16'hc44a;
35654: douta=16'hc46a;
35655: douta=16'hcc69;
35656: douta=16'hc46a;
35657: douta=16'hc469;
35658: douta=16'hc46a;
35659: douta=16'hc449;
35660: douta=16'hc449;
35661: douta=16'hc46a;
35662: douta=16'hc44a;
35663: douta=16'hc469;
35664: douta=16'hc469;
35665: douta=16'hc44a;
35666: douta=16'hc44a;
35667: douta=16'hc44a;
35668: douta=16'hc42a;
35669: douta=16'hc44a;
35670: douta=16'hc42a;
35671: douta=16'hbc2a;
35672: douta=16'hc44a;
35673: douta=16'hc42a;
35674: douta=16'hbc2a;
35675: douta=16'hbc2a;
35676: douta=16'hbc2a;
35677: douta=16'hbc29;
35678: douta=16'hbc2a;
35679: douta=16'hbc2a;
35680: douta=16'hbc0a;
35681: douta=16'hbc0a;
35682: douta=16'hbc0a;
35683: douta=16'hbc0a;
35684: douta=16'hbc09;
35685: douta=16'hbc09;
35686: douta=16'hbc09;
35687: douta=16'hbbe9;
35688: douta=16'hbbe9;
35689: douta=16'hb3e9;
35690: douta=16'hbbe9;
35691: douta=16'hbbe9;
35692: douta=16'hb3e9;
35693: douta=16'hb3e9;
35694: douta=16'hb3e9;
35695: douta=16'hb3ca;
35696: douta=16'hb3c9;
35697: douta=16'hb3c9;
35698: douta=16'hb3e9;
35699: douta=16'habc9;
35700: douta=16'habc9;
35701: douta=16'haba9;
35702: douta=16'haba9;
35703: douta=16'haba9;
35704: douta=16'haba9;
35705: douta=16'haba9;
35706: douta=16'haba9;
35707: douta=16'ha389;
35708: douta=16'ha389;
35709: douta=16'ha389;
35710: douta=16'ha369;
35711: douta=16'ha389;
35712: douta=16'h2124;
35713: douta=16'h3145;
35714: douta=16'h3125;
35715: douta=16'h2924;
35716: douta=16'h3124;
35717: douta=16'h2904;
35718: douta=16'h2924;
35719: douta=16'h2904;
35720: douta=16'h2904;
35721: douta=16'h2904;
35722: douta=16'h2104;
35723: douta=16'h2104;
35724: douta=16'h28e3;
35725: douta=16'h20c3;
35726: douta=16'h20c3;
35727: douta=16'h20e3;
35728: douta=16'h28e3;
35729: douta=16'h2903;
35730: douta=16'h2903;
35731: douta=16'h3103;
35732: douta=16'h3103;
35733: douta=16'h3103;
35734: douta=16'h3123;
35735: douta=16'h3923;
35736: douta=16'h3923;
35737: douta=16'h4144;
35738: douta=16'h4143;
35739: douta=16'h4984;
35740: douta=16'h4185;
35741: douta=16'h4229;
35742: douta=16'h18e5;
35743: douta=16'h6205;
35744: douta=16'h59e4;
35745: douta=16'h6205;
35746: douta=16'h6205;
35747: douta=16'h6205;
35748: douta=16'h6a25;
35749: douta=16'h6a25;
35750: douta=16'h7224;
35751: douta=16'h72ea;
35752: douta=16'h8285;
35753: douta=16'h8285;
35754: douta=16'h7a85;
35755: douta=16'h82c6;
35756: douta=16'h82c6;
35757: douta=16'h82c6;
35758: douta=16'h8ac7;
35759: douta=16'h8ac6;
35760: douta=16'h8b07;
35761: douta=16'h9307;
35762: douta=16'h9307;
35763: douta=16'h9307;
35764: douta=16'h9327;
35765: douta=16'h9b47;
35766: douta=16'h9b68;
35767: douta=16'h9b68;
35768: douta=16'h9b68;
35769: douta=16'h9b68;
35770: douta=16'ha368;
35771: douta=16'ha388;
35772: douta=16'ha388;
35773: douta=16'habc8;
35774: douta=16'hb3e8;
35775: douta=16'hb3e8;
35776: douta=16'hbc08;
35777: douta=16'hb3e8;
35778: douta=16'hbc29;
35779: douta=16'hbc09;
35780: douta=16'hbc09;
35781: douta=16'hbc09;
35782: douta=16'hbc09;
35783: douta=16'hbc29;
35784: douta=16'hbc49;
35785: douta=16'hc449;
35786: douta=16'hbc29;
35787: douta=16'hbc49;
35788: douta=16'hc449;
35789: douta=16'hc449;
35790: douta=16'hc469;
35791: douta=16'hc46a;
35792: douta=16'hc46a;
35793: douta=16'hcc6a;
35794: douta=16'hc469;
35795: douta=16'hc469;
35796: douta=16'hc469;
35797: douta=16'hc469;
35798: douta=16'hcc6a;
35799: douta=16'hcc6a;
35800: douta=16'hcc6a;
35801: douta=16'hcc69;
35802: douta=16'hcc8a;
35803: douta=16'hcc8a;
35804: douta=16'hcc8a;
35805: douta=16'hcc69;
35806: douta=16'hcc6a;
35807: douta=16'hcc6a;
35808: douta=16'hcc6a;
35809: douta=16'hcc8a;
35810: douta=16'hcc6a;
35811: douta=16'hcc69;
35812: douta=16'hcc6a;
35813: douta=16'hcc69;
35814: douta=16'hcc69;
35815: douta=16'hcc69;
35816: douta=16'hcc89;
35817: douta=16'hcc89;
35818: douta=16'hcc69;
35819: douta=16'hcc69;
35820: douta=16'hc468;
35821: douta=16'hcc89;
35822: douta=16'hcc89;
35823: douta=16'hcc69;
35824: douta=16'hcc8a;
35825: douta=16'hcc6a;
35826: douta=16'hcc6a;
35827: douta=16'hcc6a;
35828: douta=16'hcc6a;
35829: douta=16'hcc6a;
35830: douta=16'hcc6a;
35831: douta=16'hcc6a;
35832: douta=16'hcc6a;
35833: douta=16'hcc6a;
35834: douta=16'hb5d5;
35835: douta=16'he634;
35836: douta=16'hc469;
35837: douta=16'hcc6a;
35838: douta=16'hcc6a;
35839: douta=16'hcc6a;
35840: douta=16'hcc6a;
35841: douta=16'hcc69;
35842: douta=16'hcc69;
35843: douta=16'hcc69;
35844: douta=16'hcc69;
35845: douta=16'hcc6a;
35846: douta=16'hc449;
35847: douta=16'hc449;
35848: douta=16'hc46a;
35849: douta=16'hc46a;
35850: douta=16'hc44a;
35851: douta=16'hc46a;
35852: douta=16'hc469;
35853: douta=16'hc469;
35854: douta=16'hc44a;
35855: douta=16'hc44a;
35856: douta=16'hc44a;
35857: douta=16'hc44a;
35858: douta=16'hc44a;
35859: douta=16'hc429;
35860: douta=16'hc44a;
35861: douta=16'hc44a;
35862: douta=16'hc42a;
35863: douta=16'hc44a;
35864: douta=16'hc44a;
35865: douta=16'hc44a;
35866: douta=16'hc42a;
35867: douta=16'hbc2a;
35868: douta=16'hc44a;
35869: douta=16'hbc2a;
35870: douta=16'hbc2a;
35871: douta=16'hbc2a;
35872: douta=16'hbc0a;
35873: douta=16'hbc0a;
35874: douta=16'hbc0a;
35875: douta=16'hbc09;
35876: douta=16'hbc09;
35877: douta=16'hbc09;
35878: douta=16'hbc09;
35879: douta=16'hbc09;
35880: douta=16'hb3e9;
35881: douta=16'hb3e9;
35882: douta=16'hbbe9;
35883: douta=16'hb3e9;
35884: douta=16'hb3e9;
35885: douta=16'hb3e9;
35886: douta=16'hb3c9;
35887: douta=16'habc9;
35888: douta=16'hb3c9;
35889: douta=16'hb3ca;
35890: douta=16'habc9;
35891: douta=16'hb3e9;
35892: douta=16'habc9;
35893: douta=16'habca;
35894: douta=16'haba9;
35895: douta=16'haba9;
35896: douta=16'haba9;
35897: douta=16'haba9;
35898: douta=16'haba9;
35899: douta=16'haba9;
35900: douta=16'ha389;
35901: douta=16'haba9;
35902: douta=16'ha389;
35903: douta=16'ha389;
35904: douta=16'h2904;
35905: douta=16'h3125;
35906: douta=16'h2924;
35907: douta=16'h2904;
35908: douta=16'h2924;
35909: douta=16'h2924;
35910: douta=16'h28e3;
35911: douta=16'h2924;
35912: douta=16'h2904;
35913: douta=16'h2904;
35914: douta=16'h2103;
35915: douta=16'h2104;
35916: douta=16'h2924;
35917: douta=16'h20e3;
35918: douta=16'h20e3;
35919: douta=16'h20c3;
35920: douta=16'h2903;
35921: douta=16'h28e3;
35922: douta=16'h2903;
35923: douta=16'h3124;
35924: douta=16'h3104;
35925: douta=16'h3103;
35926: douta=16'h3923;
35927: douta=16'h3923;
35928: douta=16'h3923;
35929: douta=16'h4124;
35930: douta=16'h4144;
35931: douta=16'h4964;
35932: douta=16'h49c7;
35933: douta=16'h3187;
35934: douta=16'h0884;
35935: douta=16'h59c4;
35936: douta=16'h59e4;
35937: douta=16'h6205;
35938: douta=16'h6a25;
35939: douta=16'h6a25;
35940: douta=16'h7266;
35941: douta=16'h7265;
35942: douta=16'h7285;
35943: douta=16'h8430;
35944: douta=16'h7aa6;
35945: douta=16'h7aa5;
35946: douta=16'h82a6;
35947: douta=16'h82c6;
35948: douta=16'h82c6;
35949: douta=16'h82c6;
35950: douta=16'h8ac7;
35951: douta=16'h8ae7;
35952: douta=16'h8b07;
35953: douta=16'h8b07;
35954: douta=16'h8b07;
35955: douta=16'h9327;
35956: douta=16'h9b48;
35957: douta=16'h9b48;
35958: douta=16'h9b48;
35959: douta=16'h9b68;
35960: douta=16'ha388;
35961: douta=16'ha368;
35962: douta=16'ha388;
35963: douta=16'ha388;
35964: douta=16'ha388;
35965: douta=16'habc8;
35966: douta=16'hb3c8;
35967: douta=16'hb3e9;
35968: douta=16'hbc09;
35969: douta=16'hb409;
35970: douta=16'hbc09;
35971: douta=16'hbc09;
35972: douta=16'hbc2a;
35973: douta=16'hbc2a;
35974: douta=16'hbc29;
35975: douta=16'hbc29;
35976: douta=16'hc44a;
35977: douta=16'hbc49;
35978: douta=16'hbc49;
35979: douta=16'hbc49;
35980: douta=16'hc449;
35981: douta=16'hc469;
35982: douta=16'hc469;
35983: douta=16'hc469;
35984: douta=16'hc46a;
35985: douta=16'hc48a;
35986: douta=16'hcc8a;
35987: douta=16'hc469;
35988: douta=16'hc469;
35989: douta=16'hc469;
35990: douta=16'hc48a;
35991: douta=16'hc48a;
35992: douta=16'hcc6a;
35993: douta=16'hc469;
35994: douta=16'hcc6a;
35995: douta=16'hcc6a;
35996: douta=16'hc469;
35997: douta=16'hcc6a;
35998: douta=16'hcc8a;
35999: douta=16'hcc8a;
36000: douta=16'hcc6a;
36001: douta=16'hcc6a;
36002: douta=16'hcc6a;
36003: douta=16'hcc6a;
36004: douta=16'hcc6a;
36005: douta=16'hcc6a;
36006: douta=16'hc469;
36007: douta=16'hcc6a;
36008: douta=16'hcc69;
36009: douta=16'hcc69;
36010: douta=16'hcc69;
36011: douta=16'hcc69;
36012: douta=16'hcc6a;
36013: douta=16'hcc69;
36014: douta=16'hcc89;
36015: douta=16'hcc69;
36016: douta=16'hcc6a;
36017: douta=16'hcc6a;
36018: douta=16'hcc6a;
36019: douta=16'hcc6a;
36020: douta=16'hcc6a;
36021: douta=16'hc469;
36022: douta=16'hcc6a;
36023: douta=16'hcc6a;
36024: douta=16'hcc6a;
36025: douta=16'hcc6a;
36026: douta=16'hbdd6;
36027: douta=16'he634;
36028: douta=16'hcc6a;
36029: douta=16'hcc6a;
36030: douta=16'hcc6a;
36031: douta=16'hc46a;
36032: douta=16'hc46a;
36033: douta=16'hcc6a;
36034: douta=16'hcc69;
36035: douta=16'hcc69;
36036: douta=16'hcc69;
36037: douta=16'hc44a;
36038: douta=16'hc44a;
36039: douta=16'hc469;
36040: douta=16'hc46a;
36041: douta=16'hc449;
36042: douta=16'hc46a;
36043: douta=16'hc449;
36044: douta=16'hc44a;
36045: douta=16'hc44a;
36046: douta=16'hc44a;
36047: douta=16'hc44a;
36048: douta=16'hc44a;
36049: douta=16'hc44a;
36050: douta=16'hc429;
36051: douta=16'hc44a;
36052: douta=16'hc44a;
36053: douta=16'hbc2a;
36054: douta=16'hc42a;
36055: douta=16'hc42a;
36056: douta=16'hbc2a;
36057: douta=16'hbc2a;
36058: douta=16'hbc2a;
36059: douta=16'hbc2a;
36060: douta=16'hbc2a;
36061: douta=16'hbc2a;
36062: douta=16'hbc2a;
36063: douta=16'hbc0a;
36064: douta=16'hbc2a;
36065: douta=16'hbc2a;
36066: douta=16'hbc0a;
36067: douta=16'hbc09;
36068: douta=16'hbc0a;
36069: douta=16'hbc09;
36070: douta=16'hbbe9;
36071: douta=16'hbbe9;
36072: douta=16'hbbe9;
36073: douta=16'hb3e9;
36074: douta=16'hb3ea;
36075: douta=16'hb3e9;
36076: douta=16'hb3e9;
36077: douta=16'hb3e9;
36078: douta=16'hb3e9;
36079: douta=16'hb3ca;
36080: douta=16'habc9;
36081: douta=16'habc9;
36082: douta=16'habca;
36083: douta=16'haba9;
36084: douta=16'haba9;
36085: douta=16'haba9;
36086: douta=16'haba9;
36087: douta=16'haba9;
36088: douta=16'hab89;
36089: douta=16'habaa;
36090: douta=16'ha389;
36091: douta=16'ha369;
36092: douta=16'ha369;
36093: douta=16'ha389;
36094: douta=16'ha38a;
36095: douta=16'ha389;
36096: douta=16'h3146;
36097: douta=16'h2945;
36098: douta=16'h2924;
36099: douta=16'h2904;
36100: douta=16'h2924;
36101: douta=16'h2904;
36102: douta=16'h2904;
36103: douta=16'h2924;
36104: douta=16'h2904;
36105: douta=16'h2904;
36106: douta=16'h2104;
36107: douta=16'h2104;
36108: douta=16'h2924;
36109: douta=16'h20e3;
36110: douta=16'h20e3;
36111: douta=16'h20e3;
36112: douta=16'h2903;
36113: douta=16'h28e3;
36114: douta=16'h2904;
36115: douta=16'h3123;
36116: douta=16'h3103;
36117: douta=16'h3124;
36118: douta=16'h3923;
36119: douta=16'h3923;
36120: douta=16'h3944;
36121: douta=16'h4164;
36122: douta=16'h4164;
36123: douta=16'h4964;
36124: douta=16'h526a;
36125: douta=16'h1906;
36126: douta=16'h0884;
36127: douta=16'h59c4;
36128: douta=16'h59e5;
36129: douta=16'h59e4;
36130: douta=16'h6a25;
36131: douta=16'h6a25;
36132: douta=16'h7246;
36133: douta=16'h7286;
36134: douta=16'h7ae9;
36135: douta=16'h9d14;
36136: douta=16'h7a86;
36137: douta=16'h82a6;
36138: douta=16'h82a6;
36139: douta=16'h82c6;
36140: douta=16'h82c6;
36141: douta=16'h8ae6;
36142: douta=16'h8ae7;
36143: douta=16'h8ae7;
36144: douta=16'h8b07;
36145: douta=16'h8ae7;
36146: douta=16'h8b07;
36147: douta=16'h9327;
36148: douta=16'h9b48;
36149: douta=16'h9b28;
36150: douta=16'h9b48;
36151: douta=16'ha388;
36152: douta=16'ha388;
36153: douta=16'h9b67;
36154: douta=16'ha388;
36155: douta=16'ha387;
36156: douta=16'hab88;
36157: douta=16'habc8;
36158: douta=16'hb3e8;
36159: douta=16'hb3e9;
36160: douta=16'hb3e9;
36161: douta=16'hb409;
36162: douta=16'hbc09;
36163: douta=16'hbc2a;
36164: douta=16'hbc2a;
36165: douta=16'hbc2a;
36166: douta=16'hc42a;
36167: douta=16'hbc29;
36168: douta=16'hbc29;
36169: douta=16'hbc29;
36170: douta=16'hc449;
36171: douta=16'hc449;
36172: douta=16'hc449;
36173: douta=16'hc469;
36174: douta=16'hc449;
36175: douta=16'hc46a;
36176: douta=16'hc46a;
36177: douta=16'hcc6a;
36178: douta=16'hc46a;
36179: douta=16'hc46a;
36180: douta=16'hc46a;
36181: douta=16'hc46a;
36182: douta=16'hc48a;
36183: douta=16'hc48a;
36184: douta=16'hc469;
36185: douta=16'hcc89;
36186: douta=16'hcc8a;
36187: douta=16'hcc6a;
36188: douta=16'hcc6a;
36189: douta=16'hcc6a;
36190: douta=16'hcc6a;
36191: douta=16'hc469;
36192: douta=16'hcc8a;
36193: douta=16'hcc69;
36194: douta=16'hcc89;
36195: douta=16'hcc69;
36196: douta=16'hc469;
36197: douta=16'hcc6a;
36198: douta=16'hcc6a;
36199: douta=16'hcc69;
36200: douta=16'hcc6a;
36201: douta=16'hcc69;
36202: douta=16'hcc69;
36203: douta=16'hcc6a;
36204: douta=16'hcc69;
36205: douta=16'hcc6a;
36206: douta=16'hcc6a;
36207: douta=16'hcc69;
36208: douta=16'hcc69;
36209: douta=16'hcc6a;
36210: douta=16'hc469;
36211: douta=16'hcc69;
36212: douta=16'hcc6a;
36213: douta=16'hcc6a;
36214: douta=16'hcc6a;
36215: douta=16'hcc8a;
36216: douta=16'hcc6a;
36217: douta=16'hc46a;
36218: douta=16'hbdd6;
36219: douta=16'he634;
36220: douta=16'hcc6a;
36221: douta=16'hcc6a;
36222: douta=16'hc46a;
36223: douta=16'hc46a;
36224: douta=16'hc46a;
36225: douta=16'hc46a;
36226: douta=16'hc469;
36227: douta=16'hc449;
36228: douta=16'hc449;
36229: douta=16'hc469;
36230: douta=16'hc44a;
36231: douta=16'hc469;
36232: douta=16'hc469;
36233: douta=16'hc469;
36234: douta=16'hc469;
36235: douta=16'hc429;
36236: douta=16'hc44a;
36237: douta=16'hc44a;
36238: douta=16'hc44a;
36239: douta=16'hc44a;
36240: douta=16'hc44a;
36241: douta=16'hc44a;
36242: douta=16'hc44a;
36243: douta=16'hc429;
36244: douta=16'hbc2a;
36245: douta=16'hc44a;
36246: douta=16'hc42a;
36247: douta=16'hc44a;
36248: douta=16'hbc2a;
36249: douta=16'hc42a;
36250: douta=16'hbc2a;
36251: douta=16'hbc2a;
36252: douta=16'hbc2a;
36253: douta=16'hbc2a;
36254: douta=16'hbc2a;
36255: douta=16'hbc2a;
36256: douta=16'hbc2a;
36257: douta=16'hbc09;
36258: douta=16'hbc09;
36259: douta=16'hbc09;
36260: douta=16'hbc09;
36261: douta=16'hbc09;
36262: douta=16'hbbe9;
36263: douta=16'hb3ea;
36264: douta=16'hb40a;
36265: douta=16'hb3ea;
36266: douta=16'hb3e9;
36267: douta=16'hb3e9;
36268: douta=16'hb3ea;
36269: douta=16'hb3ca;
36270: douta=16'hb3ca;
36271: douta=16'hb3ca;
36272: douta=16'hb3e9;
36273: douta=16'hb3e9;
36274: douta=16'habca;
36275: douta=16'haba9;
36276: douta=16'haba9;
36277: douta=16'haba9;
36278: douta=16'haba9;
36279: douta=16'haba9;
36280: douta=16'habaa;
36281: douta=16'ha389;
36282: douta=16'habaa;
36283: douta=16'hab89;
36284: douta=16'ha369;
36285: douta=16'hab89;
36286: douta=16'ha369;
36287: douta=16'ha389;
36288: douta=16'h3145;
36289: douta=16'h2925;
36290: douta=16'h2924;
36291: douta=16'h2904;
36292: douta=16'h2904;
36293: douta=16'h2904;
36294: douta=16'h2904;
36295: douta=16'h2924;
36296: douta=16'h2904;
36297: douta=16'h2904;
36298: douta=16'h2104;
36299: douta=16'h2104;
36300: douta=16'h2104;
36301: douta=16'h20e3;
36302: douta=16'h20e3;
36303: douta=16'h20e3;
36304: douta=16'h2903;
36305: douta=16'h2903;
36306: douta=16'h28e3;
36307: douta=16'h3103;
36308: douta=16'h3103;
36309: douta=16'h3123;
36310: douta=16'h3924;
36311: douta=16'h3923;
36312: douta=16'h3944;
36313: douta=16'h4964;
36314: douta=16'h4164;
36315: douta=16'h4985;
36316: douta=16'h5aab;
36317: douta=16'h18e5;
36318: douta=16'h1084;
36319: douta=16'h51c4;
36320: douta=16'h6205;
36321: douta=16'h59e5;
36322: douta=16'h6a25;
36323: douta=16'h6a45;
36324: douta=16'h7246;
36325: douta=16'h7265;
36326: douta=16'h732b;
36327: douta=16'ha576;
36328: douta=16'h82c7;
36329: douta=16'h82a6;
36330: douta=16'h82a6;
36331: douta=16'h82c6;
36332: douta=16'h8ae7;
36333: douta=16'h8ae7;
36334: douta=16'h8ac7;
36335: douta=16'h8b07;
36336: douta=16'h8b07;
36337: douta=16'h8b07;
36338: douta=16'h9308;
36339: douta=16'h9327;
36340: douta=16'h9b48;
36341: douta=16'h9b48;
36342: douta=16'h9b48;
36343: douta=16'ha368;
36344: douta=16'ha388;
36345: douta=16'h9b67;
36346: douta=16'ha388;
36347: douta=16'ha387;
36348: douta=16'ha387;
36349: douta=16'habc8;
36350: douta=16'hb3c9;
36351: douta=16'hb409;
36352: douta=16'hb409;
36353: douta=16'hb409;
36354: douta=16'hb409;
36355: douta=16'hbc2a;
36356: douta=16'hc42a;
36357: douta=16'hc42a;
36358: douta=16'hbc2a;
36359: douta=16'hc44a;
36360: douta=16'hbc29;
36361: douta=16'hbc29;
36362: douta=16'hc44a;
36363: douta=16'hbc49;
36364: douta=16'hc44a;
36365: douta=16'hc469;
36366: douta=16'hc449;
36367: douta=16'hcc6a;
36368: douta=16'hc46a;
36369: douta=16'hcc6a;
36370: douta=16'hc46a;
36371: douta=16'hc46a;
36372: douta=16'hc46a;
36373: douta=16'hc46a;
36374: douta=16'hc48a;
36375: douta=16'hc48a;
36376: douta=16'hcc6a;
36377: douta=16'hcc6a;
36378: douta=16'hcc8a;
36379: douta=16'hcc6a;
36380: douta=16'hcc8a;
36381: douta=16'hcc8a;
36382: douta=16'hcc6a;
36383: douta=16'hcc6a;
36384: douta=16'hcc6a;
36385: douta=16'hcc69;
36386: douta=16'hc489;
36387: douta=16'hc489;
36388: douta=16'hcc6a;
36389: douta=16'hcc6a;
36390: douta=16'hcc69;
36391: douta=16'hcc69;
36392: douta=16'hcc69;
36393: douta=16'hcc49;
36394: douta=16'hcc69;
36395: douta=16'hcc69;
36396: douta=16'hcc6a;
36397: douta=16'hcc69;
36398: douta=16'hcc69;
36399: douta=16'hcc69;
36400: douta=16'hcc6a;
36401: douta=16'hcc6a;
36402: douta=16'hc469;
36403: douta=16'hcc6a;
36404: douta=16'hcc6a;
36405: douta=16'hcc8a;
36406: douta=16'hc469;
36407: douta=16'hcc8a;
36408: douta=16'hcc6a;
36409: douta=16'hc46a;
36410: douta=16'hbdd6;
36411: douta=16'hde33;
36412: douta=16'hc46a;
36413: douta=16'hc46a;
36414: douta=16'hc46a;
36415: douta=16'hc46a;
36416: douta=16'hc46a;
36417: douta=16'hc46a;
36418: douta=16'hc469;
36419: douta=16'hc469;
36420: douta=16'hc469;
36421: douta=16'hc449;
36422: douta=16'hc449;
36423: douta=16'hc469;
36424: douta=16'hc46a;
36425: douta=16'hc469;
36426: douta=16'hc449;
36427: douta=16'hc44a;
36428: douta=16'hc44a;
36429: douta=16'hc44a;
36430: douta=16'hc44a;
36431: douta=16'hc44a;
36432: douta=16'hc44a;
36433: douta=16'hc44a;
36434: douta=16'hc429;
36435: douta=16'hc44a;
36436: douta=16'hc42a;
36437: douta=16'hc42a;
36438: douta=16'hbc2a;
36439: douta=16'hc44a;
36440: douta=16'hbc2a;
36441: douta=16'hbc2a;
36442: douta=16'hbc2a;
36443: douta=16'hbc2a;
36444: douta=16'hbc2a;
36445: douta=16'hbc0a;
36446: douta=16'hbc2a;
36447: douta=16'hbc0a;
36448: douta=16'hbc0a;
36449: douta=16'hbc0a;
36450: douta=16'hbc0a;
36451: douta=16'hbc0a;
36452: douta=16'hbc09;
36453: douta=16'hbc09;
36454: douta=16'hb40a;
36455: douta=16'hb3ea;
36456: douta=16'hb3e9;
36457: douta=16'hb3e9;
36458: douta=16'hb3e9;
36459: douta=16'hb3ea;
36460: douta=16'hb3ca;
36461: douta=16'hb3ca;
36462: douta=16'hb3ca;
36463: douta=16'hb3c9;
36464: douta=16'habc9;
36465: douta=16'habc9;
36466: douta=16'habca;
36467: douta=16'habca;
36468: douta=16'haba9;
36469: douta=16'haba9;
36470: douta=16'haba9;
36471: douta=16'hab89;
36472: douta=16'hab89;
36473: douta=16'ha389;
36474: douta=16'ha389;
36475: douta=16'ha389;
36476: douta=16'ha369;
36477: douta=16'ha389;
36478: douta=16'hab89;
36479: douta=16'ha369;
36480: douta=16'h2945;
36481: douta=16'h2924;
36482: douta=16'h2924;
36483: douta=16'h2104;
36484: douta=16'h2924;
36485: douta=16'h2104;
36486: douta=16'h2104;
36487: douta=16'h2904;
36488: douta=16'h2104;
36489: douta=16'h2104;
36490: douta=16'h2104;
36491: douta=16'h2104;
36492: douta=16'h20e3;
36493: douta=16'h20c3;
36494: douta=16'h28e3;
36495: douta=16'h28e3;
36496: douta=16'h2903;
36497: douta=16'h2904;
36498: douta=16'h3104;
36499: douta=16'h3124;
36500: douta=16'h3124;
36501: douta=16'h3124;
36502: douta=16'h3944;
36503: douta=16'h3944;
36504: douta=16'h3944;
36505: douta=16'h4164;
36506: douta=16'h4985;
36507: douta=16'h4985;
36508: douta=16'h5aaa;
36509: douta=16'h0884;
36510: douta=16'h28e3;
36511: douta=16'h59c4;
36512: douta=16'h59e4;
36513: douta=16'h6205;
36514: douta=16'h6a25;
36515: douta=16'h6a45;
36516: douta=16'h7266;
36517: douta=16'h7266;
36518: douta=16'h8430;
36519: douta=16'hbe17;
36520: douta=16'h82a6;
36521: douta=16'h82c7;
36522: douta=16'h82c7;
36523: douta=16'h82c6;
36524: douta=16'h8ae6;
36525: douta=16'h8ae7;
36526: douta=16'h8ae7;
36527: douta=16'h8b07;
36528: douta=16'h8b07;
36529: douta=16'h8b07;
36530: douta=16'h8b07;
36531: douta=16'h9308;
36532: douta=16'h9348;
36533: douta=16'h9b48;
36534: douta=16'h9b48;
36535: douta=16'h9b68;
36536: douta=16'h9b68;
36537: douta=16'h9b68;
36538: douta=16'ha388;
36539: douta=16'ha388;
36540: douta=16'ha388;
36541: douta=16'habc8;
36542: douta=16'habe9;
36543: douta=16'hb3e9;
36544: douta=16'hb409;
36545: douta=16'hb409;
36546: douta=16'hb409;
36547: douta=16'hbc2a;
36548: douta=16'hbc2a;
36549: douta=16'hbc2a;
36550: douta=16'hc42a;
36551: douta=16'hc44a;
36552: douta=16'hbc49;
36553: douta=16'hbc29;
36554: douta=16'hbc29;
36555: douta=16'hc44a;
36556: douta=16'hbc49;
36557: douta=16'hc44a;
36558: douta=16'hc44a;
36559: douta=16'hc46a;
36560: douta=16'hc46a;
36561: douta=16'hc46a;
36562: douta=16'hc44a;
36563: douta=16'hcc6a;
36564: douta=16'hc46a;
36565: douta=16'hc46a;
36566: douta=16'hcc6a;
36567: douta=16'hc48a;
36568: douta=16'hcc6a;
36569: douta=16'hc46a;
36570: douta=16'hc469;
36571: douta=16'hc48a;
36572: douta=16'hc48a;
36573: douta=16'hc48a;
36574: douta=16'hcc8a;
36575: douta=16'hcc6a;
36576: douta=16'hcc6a;
36577: douta=16'hc469;
36578: douta=16'hc489;
36579: douta=16'hcc69;
36580: douta=16'hc469;
36581: douta=16'hcc6a;
36582: douta=16'hc469;
36583: douta=16'hcc6a;
36584: douta=16'hc469;
36585: douta=16'hcc6a;
36586: douta=16'hcc69;
36587: douta=16'hcc69;
36588: douta=16'hc469;
36589: douta=16'hcc69;
36590: douta=16'hcc6a;
36591: douta=16'hcc6a;
36592: douta=16'hcc6a;
36593: douta=16'hcc6a;
36594: douta=16'hcc6a;
36595: douta=16'hc46a;
36596: douta=16'hcc6a;
36597: douta=16'hcc6a;
36598: douta=16'hcc6a;
36599: douta=16'hcc6a;
36600: douta=16'hcc6a;
36601: douta=16'hc46a;
36602: douta=16'hbe16;
36603: douta=16'hde34;
36604: douta=16'hc46a;
36605: douta=16'hcc6a;
36606: douta=16'hc46a;
36607: douta=16'hc46a;
36608: douta=16'hc46a;
36609: douta=16'hc469;
36610: douta=16'hc46a;
36611: douta=16'hc46a;
36612: douta=16'hc469;
36613: douta=16'hc46a;
36614: douta=16'hc46a;
36615: douta=16'hc469;
36616: douta=16'hc44a;
36617: douta=16'hc44a;
36618: douta=16'hc44a;
36619: douta=16'hc429;
36620: douta=16'hc44a;
36621: douta=16'hbc29;
36622: douta=16'hc44a;
36623: douta=16'hc44a;
36624: douta=16'hbc29;
36625: douta=16'hc42a;
36626: douta=16'hc42a;
36627: douta=16'hc42a;
36628: douta=16'hc42a;
36629: douta=16'hc42a;
36630: douta=16'hbc2a;
36631: douta=16'hbc2a;
36632: douta=16'hc42a;
36633: douta=16'hbc2a;
36634: douta=16'hbc2a;
36635: douta=16'hbc2a;
36636: douta=16'hbc0a;
36637: douta=16'hbc0a;
36638: douta=16'hbc0a;
36639: douta=16'hbc0a;
36640: douta=16'hbc0a;
36641: douta=16'hbc0a;
36642: douta=16'hbc0a;
36643: douta=16'hb40a;
36644: douta=16'hb40a;
36645: douta=16'hb3ea;
36646: douta=16'hb40a;
36647: douta=16'hb40a;
36648: douta=16'hb40a;
36649: douta=16'hb3ea;
36650: douta=16'hb40a;
36651: douta=16'habc9;
36652: douta=16'hb3ea;
36653: douta=16'hb3e9;
36654: douta=16'hb3e9;
36655: douta=16'habc9;
36656: douta=16'habc9;
36657: douta=16'habc9;
36658: douta=16'haba9;
36659: douta=16'haba9;
36660: douta=16'haba9;
36661: douta=16'habaa;
36662: douta=16'habaa;
36663: douta=16'ha389;
36664: douta=16'ha389;
36665: douta=16'hab89;
36666: douta=16'habaa;
36667: douta=16'ha389;
36668: douta=16'ha389;
36669: douta=16'ha389;
36670: douta=16'ha389;
36671: douta=16'ha38a;
36672: douta=16'h3145;
36673: douta=16'h2924;
36674: douta=16'h2924;
36675: douta=16'h2924;
36676: douta=16'h2104;
36677: douta=16'h2104;
36678: douta=16'h2104;
36679: douta=16'h2924;
36680: douta=16'h2104;
36681: douta=16'h2104;
36682: douta=16'h2924;
36683: douta=16'h2924;
36684: douta=16'h20e3;
36685: douta=16'h20e3;
36686: douta=16'h20e3;
36687: douta=16'h28e3;
36688: douta=16'h2903;
36689: douta=16'h28e3;
36690: douta=16'h3103;
36691: douta=16'h3123;
36692: douta=16'h3124;
36693: douta=16'h3944;
36694: douta=16'h3944;
36695: douta=16'h4144;
36696: douta=16'h4164;
36697: douta=16'h4165;
36698: douta=16'h4185;
36699: douta=16'h4985;
36700: douta=16'h4228;
36701: douta=16'h1084;
36702: douta=16'h3944;
36703: douta=16'h59e4;
36704: douta=16'h59e4;
36705: douta=16'h59e4;
36706: douta=16'h6a25;
36707: douta=16'h6a25;
36708: douta=16'h7266;
36709: douta=16'h7244;
36710: douta=16'h94f4;
36711: douta=16'hb5b4;
36712: douta=16'h7aa6;
36713: douta=16'h82a7;
36714: douta=16'h82a7;
36715: douta=16'h8ac7;
36716: douta=16'h82c6;
36717: douta=16'h8ae6;
36718: douta=16'h8ae7;
36719: douta=16'h8b07;
36720: douta=16'h9308;
36721: douta=16'h9328;
36722: douta=16'h9328;
36723: douta=16'h9328;
36724: douta=16'h9348;
36725: douta=16'h9b48;
36726: douta=16'h9b69;
36727: douta=16'h9b68;
36728: douta=16'h9b48;
36729: douta=16'ha369;
36730: douta=16'ha388;
36731: douta=16'ha388;
36732: douta=16'ha3a8;
36733: douta=16'haba8;
36734: douta=16'hb3e9;
36735: douta=16'hb3e9;
36736: douta=16'hb409;
36737: douta=16'hb409;
36738: douta=16'hb409;
36739: douta=16'hbc2a;
36740: douta=16'hbc2a;
36741: douta=16'hbc2a;
36742: douta=16'hbc2a;
36743: douta=16'hbc2a;
36744: douta=16'hc42a;
36745: douta=16'hbc2a;
36746: douta=16'hc44a;
36747: douta=16'hc44a;
36748: douta=16'hc44a;
36749: douta=16'hc44a;
36750: douta=16'hc46b;
36751: douta=16'hc46a;
36752: douta=16'hc46a;
36753: douta=16'hc46a;
36754: douta=16'hc46a;
36755: douta=16'hc48a;
36756: douta=16'hcc6a;
36757: douta=16'hcc6a;
36758: douta=16'hc46a;
36759: douta=16'hc46a;
36760: douta=16'hcc8a;
36761: douta=16'hcc8a;
36762: douta=16'hcc8a;
36763: douta=16'hcc8a;
36764: douta=16'hc46a;
36765: douta=16'hc469;
36766: douta=16'hc469;
36767: douta=16'hcc6a;
36768: douta=16'hc469;
36769: douta=16'hcc8a;
36770: douta=16'hcc6a;
36771: douta=16'hc469;
36772: douta=16'hcc6a;
36773: douta=16'hcc6a;
36774: douta=16'hcc6a;
36775: douta=16'hc469;
36776: douta=16'hc469;
36777: douta=16'hcc6a;
36778: douta=16'hc469;
36779: douta=16'hcc6a;
36780: douta=16'hcc6a;
36781: douta=16'hcc6a;
36782: douta=16'hc46a;
36783: douta=16'hc46a;
36784: douta=16'hcc6a;
36785: douta=16'hcc6a;
36786: douta=16'hcc6a;
36787: douta=16'hcc6a;
36788: douta=16'hcc6a;
36789: douta=16'hcc6a;
36790: douta=16'hc469;
36791: douta=16'hc46a;
36792: douta=16'hcc6a;
36793: douta=16'hc46a;
36794: douta=16'hbe16;
36795: douta=16'hde13;
36796: douta=16'hc46a;
36797: douta=16'hc469;
36798: douta=16'hc46a;
36799: douta=16'hc469;
36800: douta=16'hc469;
36801: douta=16'hc46a;
36802: douta=16'hc46a;
36803: douta=16'hc469;
36804: douta=16'hc469;
36805: douta=16'hcc6a;
36806: douta=16'hc46a;
36807: douta=16'hc469;
36808: douta=16'hc44a;
36809: douta=16'hc44a;
36810: douta=16'hc44a;
36811: douta=16'hc44a;
36812: douta=16'hc44a;
36813: douta=16'hc44a;
36814: douta=16'hc44a;
36815: douta=16'hc44a;
36816: douta=16'hc44a;
36817: douta=16'hbc2a;
36818: douta=16'hc44a;
36819: douta=16'hc44a;
36820: douta=16'hbc2a;
36821: douta=16'hc42a;
36822: douta=16'hc42a;
36823: douta=16'hbc2a;
36824: douta=16'hbc2a;
36825: douta=16'hbc0a;
36826: douta=16'hbc2a;
36827: douta=16'hbc2a;
36828: douta=16'hbc0a;
36829: douta=16'hbc0a;
36830: douta=16'hbc0a;
36831: douta=16'hbc0a;
36832: douta=16'hbc09;
36833: douta=16'hbc09;
36834: douta=16'hbc0a;
36835: douta=16'hbc0a;
36836: douta=16'hb40a;
36837: douta=16'hb3ea;
36838: douta=16'hb40a;
36839: douta=16'hb3ea;
36840: douta=16'hb40a;
36841: douta=16'hb3ea;
36842: douta=16'hb3ea;
36843: douta=16'hb3e9;
36844: douta=16'hb3ca;
36845: douta=16'habca;
36846: douta=16'habca;
36847: douta=16'hb3ca;
36848: douta=16'habca;
36849: douta=16'haba9;
36850: douta=16'haba9;
36851: douta=16'haba9;
36852: douta=16'habaa;
36853: douta=16'habaa;
36854: douta=16'habaa;
36855: douta=16'habaa;
36856: douta=16'habaa;
36857: douta=16'hab89;
36858: douta=16'ha389;
36859: douta=16'ha389;
36860: douta=16'ha389;
36861: douta=16'ha38a;
36862: douta=16'ha38a;
36863: douta=16'ha369;

default :douta  =	16'h	0000;
endcase
end


endmodule 
