
module bufferram (
  input [15:0] addra,      
  output reg [15:0] douta 
);

always@(*) begin
  case(addra)
0: douta=16'h328f;
1: douta=16'h5373;
2: douta=16'h5bb4;
3: douta=16'h53f6;
4: douta=16'h4af0;
5: douta=16'h8cd7;
6: douta=16'h9d79;
7: douta=16'h8d18;
8: douta=16'h2127;
9: douta=16'h8494;
10: douta=16'hadb8;
11: douta=16'hded9;
12: douta=16'hdeba;
13: douta=16'ha537;
14: douta=16'h5b52;
15: douta=16'h8cb6;
16: douta=16'hdeba;
17: douta=16'hd6ba;
18: douta=16'ha557;
19: douta=16'h3a4c;
20: douta=16'h7bf3;
21: douta=16'he6da;
22: douta=16'he6da;
23: douta=16'h8434;
24: douta=16'h7c95;
25: douta=16'ha536;
26: douta=16'hb5f9;
27: douta=16'h7436;
28: douta=16'hb597;
29: douta=16'hbdf8;
30: douta=16'he6da;
31: douta=16'hc5f8;
32: douta=16'h63b4;
33: douta=16'h9559;
34: douta=16'h9535;
35: douta=16'had75;
36: douta=16'he6ba;
37: douta=16'h8c97;
38: douta=16'h53b3;
39: douta=16'h6c15;
40: douta=16'h6bf2;
41: douta=16'h84b5;
42: douta=16'hd67a;
43: douta=16'h5373;
44: douta=16'h3b12;
45: douta=16'h6c55;
46: douta=16'hbe7b;
47: douta=16'hd69b;
48: douta=16'h4b52;
49: douta=16'h19ee;
50: douta=16'h74b8;
51: douta=16'ha5ba;
52: douta=16'hceba;
53: douta=16'had98;
54: douta=16'h9558;
55: douta=16'h7c55;
56: douta=16'h7c98;
57: douta=16'hb67c;
58: douta=16'h4b53;
59: douta=16'h7c12;
60: douta=16'h94d4;
61: douta=16'h9d16;
62: douta=16'hd6bb;
63: douta=16'h8cd6;
64: douta=16'h7454;
65: douta=16'h8c93;
66: douta=16'ha514;
67: douta=16'hce16;
68: douta=16'hbd96;
69: douta=16'h524a;
70: douta=16'h9d13;
71: douta=16'h8c72;
72: douta=16'h8473;
73: douta=16'h1989;
74: douta=16'h8430;
75: douta=16'hce56;
76: douta=16'h83cf;
77: douta=16'h52ac;
78: douta=16'h6bd1;
79: douta=16'h52ed;
80: douta=16'h322a;
81: douta=16'hef3a;
82: douta=16'ha4d4;
83: douta=16'h5b2f;
84: douta=16'h3a0a;
85: douta=16'h6b8f;
86: douta=16'h8c92;
87: douta=16'h9c92;
88: douta=16'h4b0f;
89: douta=16'h5371;
90: douta=16'h4aef;
91: douta=16'h4aae;
92: douta=16'hd677;
93: douta=16'h2145;
94: douta=16'h10e5;
95: douta=16'h320b;
96: douta=16'h00a6;
97: douta=16'h6370;
98: douta=16'h738f;
99: douta=16'h5b31;
100: douta=16'h94d4;
101: douta=16'h73f2;
102: douta=16'h63f3;
103: douta=16'had57;
104: douta=16'h5393;
105: douta=16'h6bd1;
106: douta=16'hce79;
107: douta=16'h7455;
108: douta=16'h6415;
109: douta=16'h3af0;
110: douta=16'h2a6f;
111: douta=16'had98;
112: douta=16'h8cb5;
113: douta=16'h220e;
114: douta=16'h32b0;
115: douta=16'h5393;
116: douta=16'h7476;
117: douta=16'h6436;
118: douta=16'h3b12;
119: douta=16'h3b12;
120: douta=16'h84b8;
121: douta=16'h326f;
122: douta=16'h5416;
123: douta=16'h6478;
124: douta=16'h6435;
125: douta=16'h4395;
126: douta=16'h32d1;
127: douta=16'h6c77;
128: douta=16'h2a8f;
129: douta=16'h6457;
130: douta=16'h4b73;
131: douta=16'h53f5;
132: douta=16'h7c55;
133: douta=16'h9517;
134: douta=16'h8cb5;
135: douta=16'h5311;
136: douta=16'h5351;
137: douta=16'had98;
138: douta=16'h9d78;
139: douta=16'h8455;
140: douta=16'had78;
141: douta=16'h8c95;
142: douta=16'h9cd6;
143: douta=16'h84d7;
144: douta=16'he6da;
145: douta=16'hbdd8;
146: douta=16'h8c94;
147: douta=16'ha598;
148: douta=16'hb597;
149: douta=16'hbdb6;
150: douta=16'had76;
151: douta=16'h73f2;
152: douta=16'hce58;
153: douta=16'h73b2;
154: douta=16'h7c76;
155: douta=16'h4333;
156: douta=16'hd678;
157: douta=16'hbe7a;
158: douta=16'hc5d7;
159: douta=16'h9d36;
160: douta=16'h5331;
161: douta=16'hd658;
162: douta=16'h9d37;
163: douta=16'hd6b9;
164: douta=16'hce5a;
165: douta=16'h3b11;
166: douta=16'h8cd5;
167: douta=16'hc5f8;
168: douta=16'hf79c;
169: douta=16'hc67a;
170: douta=16'h7c33;
171: douta=16'h2af0;
172: douta=16'h9d36;
173: douta=16'h9d58;
174: douta=16'h7476;
175: douta=16'h8c95;
176: douta=16'h42d0;
177: douta=16'h84d6;
178: douta=16'h7d3a;
179: douta=16'h8538;
180: douta=16'h5bf4;
181: douta=16'h9599;
182: douta=16'ha5b9;
183: douta=16'hbe39;
184: douta=16'h9cd7;
185: douta=16'h3b32;
186: douta=16'h6bd3;
187: douta=16'hce59;
188: douta=16'had97;
189: douta=16'ha536;
190: douta=16'h5bb3;
191: douta=16'h21cd;
192: douta=16'hbe59;
193: douta=16'had55;
194: douta=16'h5b0e;
195: douta=16'h2188;
196: douta=16'h73f1;
197: douta=16'ha555;
198: douta=16'hd5f6;
199: douta=16'h5aee;
200: douta=16'h6b2e;
201: douta=16'h9cd3;
202: douta=16'heed8;
203: douta=16'h8c51;
204: douta=16'h2967;
205: douta=16'h634e;
206: douta=16'h4aad;
207: douta=16'hbdb5;
208: douta=16'h630d;
209: douta=16'h8c71;
210: douta=16'h21a9;
211: douta=16'h636f;
212: douta=16'hb554;
213: douta=16'h73d0;
214: douta=16'h42f0;
215: douta=16'h6391;
216: douta=16'h3a6c;
217: douta=16'h2989;
218: douta=16'h8c72;
219: douta=16'h9cf3;
220: douta=16'h2a4e;
221: douta=16'h2105;
222: douta=16'h10c4;
223: douta=16'h3a4c;
224: douta=16'hb594;
225: douta=16'h52ce;
226: douta=16'h6371;
227: douta=16'h7bf1;
228: douta=16'h94b3;
229: douta=16'h9d37;
230: douta=16'h530f;
231: douta=16'h2a2d;
232: douta=16'h7c32;
233: douta=16'hbdb7;
234: douta=16'h6c56;
235: douta=16'h4b31;
236: douta=16'h9538;
237: douta=16'h6c34;
238: douta=16'h8cf9;
239: douta=16'h19ee;
240: douta=16'h2a90;
241: douta=16'h4b31;
242: douta=16'h8d17;
243: douta=16'h8d18;
244: douta=16'h7c76;
245: douta=16'h21ce;
246: douta=16'h4374;
247: douta=16'h8d18;
248: douta=16'h63f5;
249: douta=16'h6435;
250: douta=16'hae1c;
251: douta=16'h5c15;
252: douta=16'h32d2;
253: douta=16'h53d5;
254: douta=16'h74d9;
255: douta=16'h5bf7;
256: douta=16'h3b12;
257: douta=16'h3b12;
258: douta=16'h32b0;
259: douta=16'h5bd5;
260: douta=16'h6bf3;
261: douta=16'h6bf4;
262: douta=16'h5372;
263: douta=16'h6392;
264: douta=16'hbdf9;
265: douta=16'hb5d9;
266: douta=16'ha5ba;
267: douta=16'h94b6;
268: douta=16'ha557;
269: douta=16'h94b4;
270: douta=16'hb5d9;
271: douta=16'h7476;
272: douta=16'h94d5;
273: douta=16'h7413;
274: douta=16'hadb8;
275: douta=16'hde79;
276: douta=16'h8cd6;
277: douta=16'h94d4;
278: douta=16'hde99;
279: douta=16'hbdf8;
280: douta=16'hde79;
281: douta=16'h6371;
282: douta=16'h6370;
283: douta=16'h7413;
284: douta=16'hff7b;
285: douta=16'hc6bb;
286: douta=16'hb596;
287: douta=16'h8c94;
288: douta=16'h9d56;
289: douta=16'he73c;
290: douta=16'h6c54;
291: douta=16'hc619;
292: douta=16'h9d58;
293: douta=16'hb5b8;
294: douta=16'hce18;
295: douta=16'hce17;
296: douta=16'hdefa;
297: douta=16'h63b3;
298: douta=16'h7c33;
299: douta=16'hc638;
300: douta=16'hce39;
301: douta=16'hd65b;
302: douta=16'h3aaf;
303: douta=16'ha5b8;
304: douta=16'hce7a;
305: douta=16'hadb9;
306: douta=16'h63d4;
307: douta=16'h2a6f;
308: douta=16'h63f4;
309: douta=16'h9579;
310: douta=16'hce7b;
311: douta=16'hbe3a;
312: douta=16'hbdb8;
313: douta=16'h5b93;
314: douta=16'h5bb2;
315: douta=16'hb65a;
316: douta=16'h3aae;
317: douta=16'h9515;
318: douta=16'h8cb6;
319: douta=16'h7c95;
320: douta=16'hb619;
321: douta=16'h7c13;
322: douta=16'h634f;
323: douta=16'h63af;
324: douta=16'ha533;
325: douta=16'h73d0;
326: douta=16'h3a2c;
327: douta=16'h6b90;
328: douta=16'hbd95;
329: douta=16'h8bf0;
330: douta=16'h4a8c;
331: douta=16'h636e;
332: douta=16'hadb5;
333: douta=16'had35;
334: douta=16'h9c0f;
335: douta=16'h1905;
336: douta=16'h422a;
337: douta=16'h94d4;
338: douta=16'h8c94;
339: douta=16'h6b90;
340: douta=16'h3a2b;
341: douta=16'h31ca;
342: douta=16'h5b6f;
343: douta=16'h8473;
344: douta=16'hce78;
345: douta=16'he658;
346: douta=16'h3a0b;
347: douta=16'h326c;
348: douta=16'h5b2e;
349: douta=16'h18a3;
350: douta=16'h10c4;
351: douta=16'h94b4;
352: douta=16'h29ca;
353: douta=16'h8453;
354: douta=16'h636f;
355: douta=16'h8452;
356: douta=16'h73f3;
357: douta=16'h21aa;
358: douta=16'h8493;
359: douta=16'h7c34;
360: douta=16'hce59;
361: douta=16'h7414;
362: douta=16'h2a2d;
363: douta=16'ha578;
364: douta=16'h6456;
365: douta=16'h63f4;
366: douta=16'h4b72;
367: douta=16'h6412;
368: douta=16'h9d57;
369: douta=16'h7414;
370: douta=16'h7498;
371: douta=16'h2250;
372: douta=16'h6c35;
373: douta=16'ha59a;
374: douta=16'h6435;
375: douta=16'h2a2e;
376: douta=16'h19ed;
377: douta=16'h8d18;
378: douta=16'h6499;
379: douta=16'h5c16;
380: douta=16'h6c77;
381: douta=16'h6c35;
382: douta=16'h53d6;
383: douta=16'h1a2e;
384: douta=16'h4bd6;
385: douta=16'h4bf6;
386: douta=16'h4b53;
387: douta=16'h7cd8;
388: douta=16'h6bd3;
389: douta=16'h5351;
390: douta=16'h6bd3;
391: douta=16'had98;
392: douta=16'hd6bd;
393: douta=16'h5bd3;
394: douta=16'h4332;
395: douta=16'h6bf1;
396: douta=16'he6da;
397: douta=16'h9d78;
398: douta=16'h9d79;
399: douta=16'h5372;
400: douta=16'h73f2;
401: douta=16'he6da;
402: douta=16'heefa;
403: douta=16'h9495;
404: douta=16'h6bf3;
405: douta=16'had97;
406: douta=16'heefa;
407: douta=16'hbdd8;
408: douta=16'h8433;
409: douta=16'h7c53;
410: douta=16'had56;
411: douta=16'ha4f5;
412: douta=16'hbdf7;
413: douta=16'h6415;
414: douta=16'hded9;
415: douta=16'he73a;
416: douta=16'h7c55;
417: douta=16'h5c36;
418: douta=16'h220d;
419: douta=16'h9515;
420: douta=16'hce59;
421: douta=16'hce7a;
422: douta=16'h5b73;
423: douta=16'h63f3;
424: douta=16'h84f9;
425: douta=16'ha557;
426: douta=16'hce9a;
427: douta=16'heed9;
428: douta=16'h4b11;
429: douta=16'h84f7;
430: douta=16'h7cb6;
431: douta=16'h8d38;
432: douta=16'hbe7c;
433: douta=16'h7c14;
434: douta=16'h7c54;
435: douta=16'h7454;
436: douta=16'hadb8;
437: douta=16'h6c98;
438: douta=16'hdf3e;
439: douta=16'h7434;
440: douta=16'h8d59;
441: douta=16'h9577;
442: douta=16'hb5f9;
443: douta=16'h5331;
444: douta=16'h29aa;
445: douta=16'h9536;
446: douta=16'h9d77;
447: douta=16'had76;
448: douta=16'h29cc;
449: douta=16'h3a4c;
450: douta=16'ha597;
451: douta=16'hef3a;
452: douta=16'h8bf0;
453: douta=16'h0885;
454: douta=16'hb595;
455: douta=16'h738f;
456: douta=16'h526b;
457: douta=16'hce14;
458: douta=16'h424a;
459: douta=16'ha512;
460: douta=16'h9431;
461: douta=16'h31ec;
462: douta=16'h428c;
463: douta=16'had75;
464: douta=16'h9c71;
465: douta=16'h8433;
466: douta=16'h1169;
467: douta=16'h0063;
468: douta=16'h7c32;
469: douta=16'ha575;
470: douta=16'hbd54;
471: douta=16'h21cb;
472: douta=16'h3a2c;
473: douta=16'h63f2;
474: douta=16'h7411;
475: douta=16'h8473;
476: douta=16'h9471;
477: douta=16'h18a3;
478: douta=16'h10a4;
479: douta=16'h2189;
480: douta=16'ha514;
481: douta=16'h7c12;
482: douta=16'h3a2b;
483: douta=16'h52cd;
484: douta=16'h428c;
485: douta=16'hff58;
486: douta=16'h9c93;
487: douta=16'h3a4c;
488: douta=16'h0129;
489: douta=16'h9d57;
490: douta=16'hb598;
491: douta=16'h9539;
492: douta=16'h63d3;
493: douta=16'h3aaf;
494: douta=16'h42cf;
495: douta=16'h5bf5;
496: douta=16'h53b4;
497: douta=16'h3af0;
498: douta=16'h5bf5;
499: douta=16'hc639;
500: douta=16'h53b4;
501: douta=16'h32d2;
502: douta=16'h4b53;
503: douta=16'h8d19;
504: douta=16'h9539;
505: douta=16'h63f5;
506: douta=16'h220d;
507: douta=16'h7497;
508: douta=16'h53f6;
509: douta=16'h5438;
510: douta=16'h2ab0;
511: douta=16'ha5da;
512: douta=16'h53d5;
513: douta=16'h5436;
514: douta=16'h53b4;
515: douta=16'h84f8;
516: douta=16'h3aaf;
517: douta=16'h6391;
518: douta=16'h7c56;
519: douta=16'hadfb;
520: douta=16'hadda;
521: douta=16'h6b92;
522: douta=16'ha578;
523: douta=16'hce59;
524: douta=16'hc618;
525: douta=16'h63d3;
526: douta=16'ha536;
527: douta=16'ha516;
528: douta=16'hd679;
529: douta=16'hbdb7;
530: douta=16'hb577;
531: douta=16'h7c95;
532: douta=16'hce18;
533: douta=16'hce38;
534: douta=16'hd698;
535: douta=16'h8c93;
536: douta=16'h8c73;
537: douta=16'he6d9;
538: douta=16'hce58;
539: douta=16'h7433;
540: douta=16'hadd7;
541: douta=16'h8c93;
542: douta=16'hf77a;
543: douta=16'hce17;
544: douta=16'h3ab0;
545: douta=16'h7474;
546: douta=16'h9d37;
547: douta=16'had97;
548: douta=16'hb619;
549: douta=16'ha576;
550: douta=16'h94d4;
551: douta=16'hd69a;
552: douta=16'h9d79;
553: douta=16'h6436;
554: douta=16'h8d58;
555: douta=16'h94f6;
556: douta=16'h9db8;
557: douta=16'hc69b;
558: douta=16'hadd9;
559: douta=16'h5416;
560: douta=16'h7498;
561: douta=16'h4aaf;
562: douta=16'h4352;
563: douta=16'ha597;
564: douta=16'hde99;
565: douta=16'h6bd4;
566: douta=16'h5bb4;
567: douta=16'ha599;
568: douta=16'h9dba;
569: douta=16'hadfa;
570: douta=16'h8c33;
571: douta=16'h1169;
572: douta=16'h9493;
573: douta=16'h8474;
574: douta=16'h6391;
575: douta=16'h52ef;
576: douta=16'h428d;
577: douta=16'h6bd2;
578: douta=16'h8474;
579: douta=16'h6bb1;
580: douta=16'h320a;
581: douta=16'h2987;
582: douta=16'h20a2;
583: douta=16'h0862;
584: douta=16'h2127;
585: douta=16'h21a9;
586: douta=16'h6baf;
587: douta=16'h8c94;
588: douta=16'h8c94;
589: douta=16'h9cb3;
590: douta=16'h6b4f;
591: douta=16'h73d1;
592: douta=16'h530f;
593: douta=16'had76;
594: douta=16'h4aad;
595: douta=16'h8452;
596: douta=16'h6b90;
597: douta=16'h8c94;
598: douta=16'h42cf;
599: douta=16'hb596;
600: douta=16'hb535;
601: douta=16'h428e;
602: douta=16'h2a2b;
603: douta=16'h6bb1;
604: douta=16'h3aae;
605: douta=16'h18a3;
606: douta=16'h10c4;
607: douta=16'h7412;
608: douta=16'h7c75;
609: douta=16'h29c9;
610: douta=16'h5b0f;
611: douta=16'h8c52;
612: douta=16'h8495;
613: douta=16'h5b51;
614: douta=16'h21ca;
615: douta=16'h7c73;
616: douta=16'hbdd7;
617: douta=16'h5bd3;
618: douta=16'h5b92;
619: douta=16'h7c95;
620: douta=16'h9536;
621: douta=16'h9517;
622: douta=16'h9538;
623: douta=16'h5373;
624: douta=16'h5bd4;
625: douta=16'hb5fa;
626: douta=16'h5c17;
627: douta=16'h6c99;
628: douta=16'h4bb5;
629: douta=16'h84b5;
630: douta=16'h8d5a;
631: douta=16'h5b94;
632: douta=16'h19ce;
633: douta=16'h326f;
634: douta=16'h7456;
635: douta=16'h7d1c;
636: douta=16'h2ad1;
637: douta=16'h5c15;
638: douta=16'hce59;
639: douta=16'h857b;
640: douta=16'h4bb5;
641: douta=16'h53f6;
642: douta=16'h5352;
643: douta=16'h6436;
644: douta=16'h42d0;
645: douta=16'h7414;
646: douta=16'h84d7;
647: douta=16'hadfb;
648: douta=16'h7c75;
649: douta=16'h8452;
650: douta=16'had77;
651: douta=16'hce59;
652: douta=16'h7350;
653: douta=16'h5352;
654: douta=16'hb577;
655: douta=16'had56;
656: douta=16'h9d37;
657: douta=16'h8474;
658: douta=16'ha515;
659: douta=16'hb598;
660: douta=16'had98;
661: douta=16'h7413;
662: douta=16'hb576;
663: douta=16'h83f2;
664: douta=16'hd678;
665: douta=16'he6ba;
666: douta=16'hbd76;
667: douta=16'h4aee;
668: douta=16'hb5d6;
669: douta=16'hbd95;
670: douta=16'hde98;
671: douta=16'had75;
672: douta=16'h7bf2;
673: douta=16'h6370;
674: douta=16'h9cd5;
675: douta=16'hb5b7;
676: douta=16'h4b94;
677: douta=16'hbe18;
678: douta=16'hbe17;
679: douta=16'hbdf9;
680: douta=16'h8cd8;
681: douta=16'h1a0e;
682: douta=16'h9d78;
683: douta=16'ha5b9;
684: douta=16'he71c;
685: douta=16'h95ba;
686: douta=16'h94d7;
687: douta=16'h4b51;
688: douta=16'h9557;
689: douta=16'had97;
690: douta=16'h7496;
691: douta=16'h6c96;
692: douta=16'h8d99;
693: douta=16'h9d78;
694: douta=16'h7c75;
695: douta=16'hb619;
696: douta=16'h84d8;
697: douta=16'h4b74;
698: douta=16'h7434;
699: douta=16'h9d36;
700: douta=16'ha4f4;
701: douta=16'h6bd1;
702: douta=16'h530f;
703: douta=16'h7c53;
704: douta=16'h8473;
705: douta=16'hb5b8;
706: douta=16'ha576;
707: douta=16'h530e;
708: douta=16'h422b;
709: douta=16'h424a;
710: douta=16'h2104;
711: douta=16'h18e3;
712: douta=16'h31c8;
713: douta=16'h29a8;
714: douta=16'h5aed;
715: douta=16'ha4f4;
716: douta=16'h2967;
717: douta=16'h320b;
718: douta=16'h8c93;
719: douta=16'hbd33;
720: douta=16'h7412;
721: douta=16'h7c31;
722: douta=16'h6b8f;
723: douta=16'hce37;
724: douta=16'h7baf;
725: douta=16'h3a2c;
726: douta=16'h7bf1;
727: douta=16'ha536;
728: douta=16'h42d0;
729: douta=16'h5b70;
730: douta=16'hc638;
731: douta=16'hbdd7;
732: douta=16'ha4d5;
733: douta=16'h1083;
734: douta=16'h08c4;
735: douta=16'h7413;
736: douta=16'h7413;
737: douta=16'h73f3;
738: douta=16'h7bf1;
739: douta=16'h5350;
740: douta=16'h2a0b;
741: douta=16'h94d4;
742: douta=16'h7413;
743: douta=16'h328f;
744: douta=16'h00c8;
745: douta=16'h42ad;
746: douta=16'h63b1;
747: douta=16'h9517;
748: douta=16'hadb9;
749: douta=16'h6392;
750: douta=16'h3ad1;
751: douta=16'h7436;
752: douta=16'h84d8;
753: douta=16'h7cda;
754: douta=16'h9559;
755: douta=16'h2a2d;
756: douta=16'h5373;
757: douta=16'h84f9;
758: douta=16'h116a;
759: douta=16'h5b93;
760: douta=16'h9558;
761: douta=16'h5b52;
762: douta=16'h6436;
763: douta=16'h118b;
764: douta=16'h8d19;
765: douta=16'h5bb5;
766: douta=16'h5c38;
767: douta=16'h3b33;
768: douta=16'h6c77;
769: douta=16'h7d1a;
770: douta=16'h42d0;
771: douta=16'h5393;
772: douta=16'h3aaf;
773: douta=16'h7434;
774: douta=16'h9538;
775: douta=16'h9d37;
776: douta=16'h6bd2;
777: douta=16'h8453;
778: douta=16'he6fb;
779: douta=16'h8c94;
780: douta=16'h5352;
781: douta=16'h324e;
782: douta=16'ha536;
783: douta=16'h9d15;
784: douta=16'h9cf6;
785: douta=16'h7413;
786: douta=16'ha555;
787: douta=16'hde98;
788: douta=16'hce38;
789: douta=16'h9493;
790: douta=16'ha576;
791: douta=16'hbdd7;
792: douta=16'hde98;
793: douta=16'hbd96;
794: douta=16'h83f1;
795: douta=16'h5aee;
796: douta=16'hc616;
797: douta=16'h8c93;
798: douta=16'h9d35;
799: douta=16'h8c93;
800: douta=16'hc5f7;
801: douta=16'h9d15;
802: douta=16'h94f6;
803: douta=16'h8cb4;
804: douta=16'ha577;
805: douta=16'hdeba;
806: douta=16'he6fb;
807: douta=16'he71c;
808: douta=16'h39c9;
809: douta=16'h8cf7;
810: douta=16'hadf9;
811: douta=16'h8538;
812: douta=16'hceba;
813: douta=16'h3af0;
814: douta=16'h73f2;
815: douta=16'h8c94;
816: douta=16'hb5b9;
817: douta=16'hb69c;
818: douta=16'h42f1;
819: douta=16'h3af0;
820: douta=16'h5373;
821: douta=16'ha5b8;
822: douta=16'ha578;
823: douta=16'hd69b;
824: douta=16'h7c75;
825: douta=16'h63f4;
826: douta=16'h3a2c;
827: douta=16'h6c12;
828: douta=16'hadb7;
829: douta=16'h5350;
830: douta=16'h5b2f;
831: douta=16'h7c53;
832: douta=16'h8c74;
833: douta=16'h324b;
834: douta=16'h430e;
835: douta=16'h4aef;
836: douta=16'hde98;
837: douta=16'h8c32;
838: douta=16'h528a;
839: douta=16'h2104;
840: douta=16'h5b0c;
841: douta=16'h73d0;
842: douta=16'hc637;
843: douta=16'h29ca;
844: douta=16'h5b2d;
845: douta=16'h73d1;
846: douta=16'h9c92;
847: douta=16'h31ea;
848: douta=16'h52ed;
849: douta=16'h5b4e;
850: douta=16'h73d1;
851: douta=16'h8c11;
852: douta=16'h0928;
853: douta=16'h6bd2;
854: douta=16'hbe77;
855: douta=16'h8cb3;
856: douta=16'h4aac;
857: douta=16'h428c;
858: douta=16'h328c;
859: douta=16'h08e6;
860: douta=16'h08e6;
861: douta=16'h10a3;
862: douta=16'h10a3;
863: douta=16'h8cf4;
864: douta=16'h84d5;
865: douta=16'h63b1;
866: douta=16'h8493;
867: douta=16'h5b70;
868: douta=16'h9cb2;
869: douta=16'h2a4d;
870: douta=16'h4aef;
871: douta=16'h7474;
872: douta=16'h7434;
873: douta=16'h8474;
874: douta=16'h29ec;
875: douta=16'h29ed;
876: douta=16'h5bd5;
877: douta=16'h5bd4;
878: douta=16'h9d78;
879: douta=16'ha5da;
880: douta=16'h6c35;
881: douta=16'h4b31;
882: douta=16'h5373;
883: douta=16'h8519;
884: douta=16'h53b5;
885: douta=16'h118c;
886: douta=16'h7455;
887: douta=16'h84d7;
888: douta=16'h3aaf;
889: douta=16'h5bd3;
890: douta=16'h6414;
891: douta=16'h4353;
892: douta=16'h4bf7;
893: douta=16'h4373;
894: douta=16'h8d5b;
895: douta=16'h9ddc;
896: douta=16'h5b93;
897: douta=16'h6498;
898: douta=16'h5bf5;
899: douta=16'h4352;
900: douta=16'h63d3;
901: douta=16'h8518;
902: douta=16'h4b31;
903: douta=16'h426e;
904: douta=16'h6392;
905: douta=16'hc5d7;
906: douta=16'had55;
907: douta=16'h8cb4;
908: douta=16'h5352;
909: douta=16'h6bd2;
910: douta=16'hbe39;
911: douta=16'hbe38;
912: douta=16'h8c95;
913: douta=16'h5b30;
914: douta=16'hbdf7;
915: douta=16'hf75a;
916: douta=16'h84b5;
917: douta=16'h9493;
918: douta=16'hce78;
919: douta=16'hdeb9;
920: douta=16'he6dc;
921: douta=16'h8c11;
922: douta=16'h4acd;
923: douta=16'h8c30;
924: douta=16'hbd95;
925: douta=16'h83f2;
926: douta=16'h9d15;
927: douta=16'h8451;
928: douta=16'hf75a;
929: douta=16'hd657;
930: douta=16'h4a8e;
931: douta=16'h4350;
932: douta=16'had77;
933: douta=16'h9d98;
934: douta=16'hc619;
935: douta=16'h9517;
936: douta=16'h8432;
937: douta=16'hd67a;
938: douta=16'h9cd6;
939: douta=16'h32f3;
940: douta=16'hbe5a;
941: douta=16'h84d7;
942: douta=16'had98;
943: douta=16'hce7b;
944: douta=16'h8475;
945: douta=16'h6c77;
946: douta=16'h4b32;
947: douta=16'h8495;
948: douta=16'h6c98;
949: douta=16'hbe9c;
950: douta=16'h7497;
951: douta=16'hbe5b;
952: douta=16'h326f;
953: douta=16'hc639;
954: douta=16'h8c52;
955: douta=16'h6bd2;
956: douta=16'h4aef;
957: douta=16'h6391;
958: douta=16'hdeda;
959: douta=16'hd5f8;
960: douta=16'h52ce;
961: douta=16'h8473;
962: douta=16'h9d15;
963: douta=16'h5b70;
964: douta=16'h8c93;
965: douta=16'h1926;
966: douta=16'ha576;
967: douta=16'h2124;
968: douta=16'h1082;
969: douta=16'h5b0e;
970: douta=16'h4aac;
971: douta=16'h634e;
972: douta=16'h8451;
973: douta=16'h9492;
974: douta=16'hb533;
975: douta=16'h8cb3;
976: douta=16'h6b6f;
977: douta=16'h6370;
978: douta=16'h1148;
979: douta=16'h1127;
980: douta=16'h0022;
981: douta=16'h0863;
982: douta=16'h0884;
983: douta=16'h08a4;
984: douta=16'h08a4;
985: douta=16'h10c4;
986: douta=16'h08a4;
987: douta=16'h0884;
988: douta=16'h0884;
989: douta=16'h0883;
990: douta=16'h0883;
991: douta=16'h0863;
992: douta=16'h0883;
993: douta=16'h0062;
994: douta=16'h0062;
995: douta=16'h0001;
996: douta=16'h0022;
997: douta=16'h42ad;
998: douta=16'h9517;
999: douta=16'h6436;
1000: douta=16'h5bb3;
1001: douta=16'h2a2d;
1002: douta=16'h5b51;
1003: douta=16'hd67a;
1004: douta=16'h84b6;
1005: douta=16'h3af2;
1006: douta=16'h222e;
1007: douta=16'h222e;
1008: douta=16'h4b53;
1009: douta=16'h7476;
1010: douta=16'h7c55;
1011: douta=16'h5351;
1012: douta=16'h3af1;
1013: douta=16'h9517;
1014: douta=16'h6415;
1015: douta=16'h32f1;
1016: douta=16'h11ac;
1017: douta=16'h6416;
1018: douta=16'h6457;
1019: douta=16'h3b13;
1020: douta=16'h5bf6;
1021: douta=16'h959c;
1022: douta=16'h6c78;
1023: douta=16'h2ad2;
1024: douta=16'h6c98;
1025: douta=16'h4b33;
1026: douta=16'h4332;
1027: douta=16'h6c15;
1028: douta=16'h5bb4;
1029: douta=16'h8495;
1030: douta=16'h63d3;
1031: douta=16'h6bd2;
1032: douta=16'h9d36;
1033: douta=16'h9d36;
1034: douta=16'h9cd4;
1035: douta=16'h6bf4;
1036: douta=16'had56;
1037: douta=16'h9d16;
1038: douta=16'hce59;
1039: douta=16'hbe19;
1040: douta=16'h94f5;
1041: douta=16'h63d2;
1042: douta=16'hd699;
1043: douta=16'hf77c;
1044: douta=16'h9cd4;
1045: douta=16'ha515;
1046: douta=16'hd6b9;
1047: douta=16'hef3b;
1048: douta=16'h94d4;
1049: douta=16'hcdf6;
1050: douta=16'hd657;
1051: douta=16'hcdf6;
1052: douta=16'h7c32;
1053: douta=16'h7bb0;
1054: douta=16'h8492;
1055: douta=16'hb595;
1056: douta=16'hef3a;
1057: douta=16'h83d0;
1058: douta=16'h6b6f;
1059: douta=16'h9472;
1060: douta=16'h7413;
1061: douta=16'h6c35;
1062: douta=16'h7c94;
1063: douta=16'h8cf5;
1064: douta=16'hc698;
1065: douta=16'hd67a;
1066: douta=16'h8cd6;
1067: douta=16'h5c36;
1068: douta=16'h7c95;
1069: douta=16'h7435;
1070: douta=16'hcedd;
1071: douta=16'h6c55;
1072: douta=16'h94d5;
1073: douta=16'h428e;
1074: douta=16'hadfa;
1075: douta=16'hd6bb;
1076: douta=16'h5b73;
1077: douta=16'h7435;
1078: douta=16'h4353;
1079: douta=16'h8d39;
1080: douta=16'h53d5;
1081: douta=16'hdeba;
1082: douta=16'h6b91;
1083: douta=16'h420a;
1084: douta=16'h7433;
1085: douta=16'h7433;
1086: douta=16'hadda;
1087: douta=16'h8474;
1088: douta=16'h73b1;
1089: douta=16'hb619;
1090: douta=16'ha4d4;
1091: douta=16'h7b6e;
1092: douta=16'h426d;
1093: douta=16'h6391;
1094: douta=16'h428d;
1095: douta=16'h18c3;
1096: douta=16'h18c4;
1097: douta=16'h2988;
1098: douta=16'h4a8b;
1099: douta=16'h8c51;
1100: douta=16'h8c10;
1101: douta=16'h3a6b;
1102: douta=16'h0083;
1103: douta=16'h0062;
1104: douta=16'h08a3;
1105: douta=16'h08a5;
1106: douta=16'h08a4;
1107: douta=16'h08c4;
1108: douta=16'h10c5;
1109: douta=16'h10c5;
1110: douta=16'h0063;
1111: douta=16'h0042;
1112: douta=16'h0022;
1113: douta=16'h0883;
1114: douta=16'h10c5;
1115: douta=16'h1906;
1116: douta=16'h1906;
1117: douta=16'h1906;
1118: douta=16'h08a4;
1119: douta=16'h0862;
1120: douta=16'h0001;
1121: douta=16'h0041;
1122: douta=16'h0883;
1123: douta=16'h0884;
1124: douta=16'h10a4;
1125: douta=16'h0884;
1126: douta=16'h0883;
1127: douta=16'h0862;
1128: douta=16'h0043;
1129: douta=16'h326c;
1130: douta=16'h8495;
1131: douta=16'h09ac;
1132: douta=16'h4b74;
1133: douta=16'h5393;
1134: douta=16'h6c56;
1135: douta=16'h7497;
1136: douta=16'h9559;
1137: douta=16'h4b31;
1138: douta=16'h21cc;
1139: douta=16'h324d;
1140: douta=16'h63f4;
1141: douta=16'h5bd3;
1142: douta=16'h4332;
1143: douta=16'h7cb6;
1144: douta=16'hb5f8;
1145: douta=16'h7cd9;
1146: douta=16'h224f;
1147: douta=16'h5bb4;
1148: douta=16'h7cb9;
1149: douta=16'h53d6;
1150: douta=16'h1a4f;
1151: douta=16'h5c37;
1152: douta=16'h326f;
1153: douta=16'h3af1;
1154: douta=16'h2a4f;
1155: douta=16'h84f9;
1156: douta=16'h7435;
1157: douta=16'h5331;
1158: douta=16'h63b2;
1159: douta=16'h6350;
1160: douta=16'ha578;
1161: douta=16'ha555;
1162: douta=16'h8433;
1163: douta=16'h7413;
1164: douta=16'h9d15;
1165: douta=16'ha576;
1166: douta=16'hbe1a;
1167: douta=16'h9516;
1168: douta=16'h9d35;
1169: douta=16'h9cf3;
1170: douta=16'he6da;
1171: douta=16'hd699;
1172: douta=16'hbd96;
1173: douta=16'ha514;
1174: douta=16'hde99;
1175: douta=16'hded9;
1176: douta=16'h6bf1;
1177: douta=16'hce16;
1178: douta=16'heed7;
1179: douta=16'h8411;
1180: douta=16'h9d14;
1181: douta=16'hc5d4;
1182: douta=16'hbd73;
1183: douta=16'h8431;
1184: douta=16'h7432;
1185: douta=16'h94b2;
1186: douta=16'hbd95;
1187: douta=16'hbd75;
1188: douta=16'h6370;
1189: douta=16'h4b50;
1190: douta=16'h9515;
1191: douta=16'ha5b8;
1192: douta=16'hce78;
1193: douta=16'hb577;
1194: douta=16'h7c74;
1195: douta=16'hb63b;
1196: douta=16'h5bd5;
1197: douta=16'h7497;
1198: douta=16'h5c15;
1199: douta=16'h32b0;
1200: douta=16'h9d78;
1201: douta=16'h9578;
1202: douta=16'hc67b;
1203: douta=16'ha61b;
1204: douta=16'h6c35;
1205: douta=16'h7c96;
1206: douta=16'h7476;
1207: douta=16'h8518;
1208: douta=16'h3b33;
1209: douta=16'hadfa;
1210: douta=16'h9d56;
1211: douta=16'h9cd3;
1212: douta=16'h5b92;
1213: douta=16'h8d37;
1214: douta=16'h7c95;
1215: douta=16'h5330;
1216: douta=16'h8473;
1217: douta=16'h8d77;
1218: douta=16'hb595;
1219: douta=16'h7cb5;
1220: douta=16'h6bf2;
1221: douta=16'h5b72;
1222: douta=16'h8474;
1223: douta=16'h6b4d;
1224: douta=16'h20e4;
1225: douta=16'h5b0d;
1226: douta=16'hce58;
1227: douta=16'h4aac;
1228: douta=16'h08c3;
1229: douta=16'h10e4;
1230: douta=16'h10e4;
1231: douta=16'h10e5;
1232: douta=16'h08a4;
1233: douta=16'h0862;
1234: douta=16'h2967;
1235: douta=16'h3a2b;
1236: douta=16'h6331;
1237: douta=16'h5b72;
1238: douta=16'h5bb4;
1239: douta=16'h63f6;
1240: douta=16'h6437;
1241: douta=16'h6c57;
1242: douta=16'h6c78;
1243: douta=16'h6c98;
1244: douta=16'h853b;
1245: douta=16'h7cf9;
1246: douta=16'h74b9;
1247: douta=16'h6c57;
1248: douta=16'h6c36;
1249: douta=16'h5b93;
1250: douta=16'h4b10;
1251: douta=16'h322d;
1252: douta=16'h2a0b;
1253: douta=16'h10e5;
1254: douta=16'h0062;
1255: douta=16'h0883;
1256: douta=16'h0884;
1257: douta=16'h08c4;
1258: douta=16'h0022;
1259: douta=16'h29e9;
1260: douta=16'h6c76;
1261: douta=16'h6c54;
1262: douta=16'h6416;
1263: douta=16'h1128;
1264: douta=16'h2a4e;
1265: douta=16'h63f3;
1266: douta=16'ha536;
1267: douta=16'h5b72;
1268: douta=16'h3a8e;
1269: douta=16'h116a;
1270: douta=16'h63d3;
1271: douta=16'h7455;
1272: douta=16'h224f;
1273: douta=16'h5b92;
1274: douta=16'h53b4;
1275: douta=16'h5c58;
1276: douta=16'h3355;
1277: douta=16'h6cb9;
1278: douta=16'h7d19;
1279: douta=16'h959b;
1280: douta=16'h4b74;
1281: douta=16'h6436;
1282: douta=16'h6c98;
1283: douta=16'h8498;
1284: douta=16'h7477;
1285: douta=16'h6b91;
1286: douta=16'h8434;
1287: douta=16'hbdf8;
1288: douta=16'h9d37;
1289: douta=16'h4aac;
1290: douta=16'h6391;
1291: douta=16'hc618;
1292: douta=16'heefa;
1293: douta=16'hdeba;
1294: douta=16'h5b92;
1295: douta=16'h4b72;
1296: douta=16'ha556;
1297: douta=16'hbdd8;
1298: douta=16'had55;
1299: douta=16'hacd3;
1300: douta=16'hb575;
1301: douta=16'hd658;
1302: douta=16'hc618;
1303: douta=16'hce37;
1304: douta=16'h6b90;
1305: douta=16'hded9;
1306: douta=16'heef9;
1307: douta=16'h6b2e;
1308: douta=16'h9451;
1309: douta=16'hbd73;
1310: douta=16'h6baf;
1311: douta=16'h5b6f;
1312: douta=16'hc636;
1313: douta=16'had32;
1314: douta=16'hde57;
1315: douta=16'h62ed;
1316: douta=16'h42ae;
1317: douta=16'h8432;
1318: douta=16'h9d15;
1319: douta=16'h5bf4;
1320: douta=16'h5392;
1321: douta=16'h632f;
1322: douta=16'hc679;
1323: douta=16'had97;
1324: douta=16'h5bb4;
1325: douta=16'h5b92;
1326: douta=16'h322e;
1327: douta=16'h5394;
1328: douta=16'h8d38;
1329: douta=16'h8d38;
1330: douta=16'h8d18;
1331: douta=16'h6c76;
1332: douta=16'h7cb8;
1333: douta=16'h7476;
1334: douta=16'h8518;
1335: douta=16'hc6de;
1336: douta=16'h73f3;
1337: douta=16'h4b31;
1338: douta=16'h21aa;
1339: douta=16'ha555;
1340: douta=16'h7c95;
1341: douta=16'h8474;
1342: douta=16'ha536;
1343: douta=16'h428d;
1344: douta=16'h8454;
1345: douta=16'h63f3;
1346: douta=16'h6bf2;
1347: douta=16'h324e;
1348: douta=16'h9517;
1349: douta=16'hc69a;
1350: douta=16'h9cd4;
1351: douta=16'h8454;
1352: douta=16'h1905;
1353: douta=16'h2167;
1354: douta=16'h18e4;
1355: douta=16'h10c5;
1356: douta=16'h18e5;
1357: douta=16'h0863;
1358: douta=16'h3147;
1359: douta=16'h5aee;
1360: douta=16'h5351;
1361: douta=16'h7499;
1362: douta=16'h855a;
1363: douta=16'h74d9;
1364: douta=16'h74d9;
1365: douta=16'h6457;
1366: douta=16'h7d3a;
1367: douta=16'h6cb8;
1368: douta=16'h74fa;
1369: douta=16'h855a;
1370: douta=16'h7cda;
1371: douta=16'h7d3a;
1372: douta=16'h6c77;
1373: douta=16'h74d9;
1374: douta=16'h6c98;
1375: douta=16'h855c;
1376: douta=16'h7d3b;
1377: douta=16'h74b8;
1378: douta=16'h6cd9;
1379: douta=16'h74fa;
1380: douta=16'h5c37;
1381: douta=16'h7d5b;
1382: douta=16'h6416;
1383: douta=16'h42af;
1384: douta=16'h322c;
1385: douta=16'h10e5;
1386: douta=16'h0883;
1387: douta=16'h10a4;
1388: douta=16'h08a4;
1389: douta=16'h0043;
1390: douta=16'h11aa;
1391: douta=16'h7c54;
1392: douta=16'h8cb6;
1393: douta=16'h5330;
1394: douta=16'h2a4d;
1395: douta=16'h7c75;
1396: douta=16'h9516;
1397: douta=16'h42f0;
1398: douta=16'h2a6f;
1399: douta=16'h2a6f;
1400: douta=16'h53d3;
1401: douta=16'h4b95;
1402: douta=16'h7499;
1403: douta=16'h4bb6;
1404: douta=16'h7cf9;
1405: douta=16'h959c;
1406: douta=16'h7d7b;
1407: douta=16'h7c77;
1408: douta=16'h224f;
1409: douta=16'h6416;
1410: douta=16'h6c78;
1411: douta=16'h42cf;
1412: douta=16'h5372;
1413: douta=16'h6371;
1414: douta=16'h8454;
1415: douta=16'h8c74;
1416: douta=16'h8495;
1417: douta=16'ha536;
1418: douta=16'hce17;
1419: douta=16'hd658;
1420: douta=16'h9d15;
1421: douta=16'h6c34;
1422: douta=16'h8433;
1423: douta=16'h7433;
1424: douta=16'hadb7;
1425: douta=16'hef3a;
1426: douta=16'h8c72;
1427: douta=16'hd678;
1428: douta=16'ha514;
1429: douta=16'hd698;
1430: douta=16'ha515;
1431: douta=16'hce37;
1432: douta=16'ha514;
1433: douta=16'hef5a;
1434: douta=16'hce16;
1435: douta=16'h83ae;
1436: douta=16'had12;
1437: douta=16'he6b8;
1438: douta=16'h632d;
1439: douta=16'h4aad;
1440: douta=16'hce15;
1441: douta=16'hc5d4;
1442: douta=16'ha512;
1443: douta=16'h9450;
1444: douta=16'h94b2;
1445: douta=16'h8431;
1446: douta=16'h6bf2;
1447: douta=16'h5b50;
1448: douta=16'h428d;
1449: douta=16'had96;
1450: douta=16'h9d76;
1451: douta=16'hc658;
1452: douta=16'hd699;
1453: douta=16'h6bd3;
1454: douta=16'h7434;
1455: douta=16'h6477;
1456: douta=16'h8d5a;
1457: douta=16'h5c15;
1458: douta=16'h4b51;
1459: douta=16'h4b73;
1460: douta=16'h6414;
1461: douta=16'h855a;
1462: douta=16'ha5b9;
1463: douta=16'h53d4;
1464: douta=16'hb5f8;
1465: douta=16'h3aaf;
1466: douta=16'h6c76;
1467: douta=16'hbe59;
1468: douta=16'h63f4;
1469: douta=16'hbe3a;
1470: douta=16'hb5b7;
1471: douta=16'h4aad;
1472: douta=16'h7c33;
1473: douta=16'h7c96;
1474: douta=16'h9473;
1475: douta=16'h3a4e;
1476: douta=16'h21ed;
1477: douta=16'h6c35;
1478: douta=16'h7496;
1479: douta=16'h1127;
1480: douta=16'h1906;
1481: douta=16'h1905;
1482: douta=16'h10c5;
1483: douta=16'h39c8;
1484: douta=16'h6b70;
1485: douta=16'h7c55;
1486: douta=16'h7cf9;
1487: douta=16'h855a;
1488: douta=16'h8d5b;
1489: douta=16'ha61c;
1490: douta=16'h7cda;
1491: douta=16'h74d9;
1492: douta=16'h74b9;
1493: douta=16'h6c98;
1494: douta=16'h5c17;
1495: douta=16'h6478;
1496: douta=16'h7d3a;
1497: douta=16'h6458;
1498: douta=16'h7cfa;
1499: douta=16'h6c98;
1500: douta=16'h857b;
1501: douta=16'h74d9;
1502: douta=16'h855b;
1503: douta=16'h74d9;
1504: douta=16'h6cb9;
1505: douta=16'h8d9b;
1506: douta=16'h74fa;
1507: douta=16'h751a;
1508: douta=16'h7d1b;
1509: douta=16'h6498;
1510: douta=16'h6478;
1511: douta=16'h7d3b;
1512: douta=16'h6cfa;
1513: douta=16'h74fa;
1514: douta=16'h5331;
1515: douta=16'h29eb;
1516: douta=16'h0863;
1517: douta=16'h10c5;
1518: douta=16'h10e5;
1519: douta=16'h0064;
1520: douta=16'h63b2;
1521: douta=16'h7c53;
1522: douta=16'h6bb2;
1523: douta=16'h8cb6;
1524: douta=16'h2a4d;
1525: douta=16'h6bd3;
1526: douta=16'had77;
1527: douta=16'h5b72;
1528: douta=16'h4bb5;
1529: douta=16'h3ad0;
1530: douta=16'h5bf5;
1531: douta=16'h6c56;
1532: douta=16'h53f6;
1533: douta=16'h53d5;
1534: douta=16'h2a2f;
1535: douta=16'h53d4;
1536: douta=16'h224f;
1537: douta=16'h6437;
1538: douta=16'h5c37;
1539: douta=16'h6415;
1540: douta=16'h63d4;
1541: douta=16'h7413;
1542: douta=16'h94b6;
1543: douta=16'h8475;
1544: douta=16'h7c96;
1545: douta=16'h8c74;
1546: douta=16'hb5b7;
1547: douta=16'had57;
1548: douta=16'ha598;
1549: douta=16'h7c54;
1550: douta=16'h7c53;
1551: douta=16'hc638;
1552: douta=16'hd678;
1553: douta=16'h94d4;
1554: douta=16'h5b2f;
1555: douta=16'hbdd6;
1556: douta=16'hb5b6;
1557: douta=16'he698;
1558: douta=16'hb5d7;
1559: douta=16'hce37;
1560: douta=16'hb575;
1561: douta=16'hef5a;
1562: douta=16'hbd74;
1563: douta=16'h9430;
1564: douta=16'hc5f5;
1565: douta=16'hd656;
1566: douta=16'h9cd1;
1567: douta=16'h52cc;
1568: douta=16'had53;
1569: douta=16'hef59;
1570: douta=16'h6bce;
1571: douta=16'hc636;
1572: douta=16'hbdf5;
1573: douta=16'hb534;
1574: douta=16'h52f0;
1575: douta=16'h3a4c;
1576: douta=16'h29eb;
1577: douta=16'h9d76;
1578: douta=16'h8cd4;
1579: douta=16'h9db8;
1580: douta=16'h8495;
1581: douta=16'h5b70;
1582: douta=16'h7c52;
1583: douta=16'h4bb4;
1584: douta=16'h3b34;
1585: douta=16'h42d0;
1586: douta=16'h5373;
1587: douta=16'h53b5;
1588: douta=16'h8518;
1589: douta=16'h5416;
1590: douta=16'h9db9;
1591: douta=16'h2a70;
1592: douta=16'h8d17;
1593: douta=16'h7c95;
1594: douta=16'h7c96;
1595: douta=16'h8cf7;
1596: douta=16'h426d;
1597: douta=16'h3aaf;
1598: douta=16'h530f;
1599: douta=16'h5b92;
1600: douta=16'hadd8;
1601: douta=16'had34;
1602: douta=16'h7bd0;
1603: douta=16'h3a8d;
1604: douta=16'h8453;
1605: douta=16'h7c75;
1606: douta=16'h2146;
1607: douta=16'h2126;
1608: douta=16'h1084;
1609: douta=16'h62ab;
1610: douta=16'h73d2;
1611: douta=16'h8d5b;
1612: douta=16'h7d19;
1613: douta=16'h853a;
1614: douta=16'h7cd9;
1615: douta=16'h8d5b;
1616: douta=16'h853a;
1617: douta=16'h853a;
1618: douta=16'h855a;
1619: douta=16'h8d3a;
1620: douta=16'h7d1a;
1621: douta=16'h7d3a;
1622: douta=16'h5bf6;
1623: douta=16'h74b9;
1624: douta=16'h857b;
1625: douta=16'h6478;
1626: douta=16'h7cfa;
1627: douta=16'h74d9;
1628: douta=16'h7d1b;
1629: douta=16'h7d1a;
1630: douta=16'h855b;
1631: douta=16'h7cfa;
1632: douta=16'h7cf9;
1633: douta=16'h6c98;
1634: douta=16'h6c99;
1635: douta=16'h7d7b;
1636: douta=16'h6cb8;
1637: douta=16'h74d9;
1638: douta=16'h7d3a;
1639: douta=16'h7d3b;
1640: douta=16'h751b;
1641: douta=16'h6cfa;
1642: douta=16'h7d3b;
1643: douta=16'h6cb9;
1644: douta=16'h6cb8;
1645: douta=16'h42af;
1646: douta=16'h2147;
1647: douta=16'h10e6;
1648: douta=16'h1106;
1649: douta=16'h0085;
1650: douta=16'h8cb6;
1651: douta=16'h2a6f;
1652: douta=16'h8452;
1653: douta=16'h73f3;
1654: douta=16'h21ec;
1655: douta=16'h32b0;
1656: douta=16'h8d39;
1657: douta=16'h7cd8;
1658: douta=16'h5416;
1659: douta=16'h32d2;
1660: douta=16'h32d2;
1661: douta=16'h7cb8;
1662: douta=16'h8d7b;
1663: douta=16'h7c97;
1664: douta=16'h116c;
1665: douta=16'h6415;
1666: douta=16'h53b5;
1667: douta=16'h6c57;
1668: douta=16'h4311;
1669: douta=16'h6bd4;
1670: douta=16'h9517;
1671: douta=16'h6bf4;
1672: douta=16'hadd9;
1673: douta=16'h5b92;
1674: douta=16'h9cf5;
1675: douta=16'had97;
1676: douta=16'h94f5;
1677: douta=16'hb5b7;
1678: douta=16'hd678;
1679: douta=16'hffdb;
1680: douta=16'he6d9;
1681: douta=16'ha534;
1682: douta=16'hce16;
1683: douta=16'hff7b;
1684: douta=16'h634f;
1685: douta=16'h4acd;
1686: douta=16'h8471;
1687: douta=16'hde98;
1688: douta=16'h94b2;
1689: douta=16'hce57;
1690: douta=16'h94b0;
1691: douta=16'hbd74;
1692: douta=16'hf71a;
1693: douta=16'ha4d0;
1694: douta=16'h4a28;
1695: douta=16'h5b0c;
1696: douta=16'h9470;
1697: douta=16'h840f;
1698: douta=16'h7c10;
1699: douta=16'h94b2;
1700: douta=16'hc636;
1701: douta=16'hde77;
1702: douta=16'h7bf1;
1703: douta=16'h5aaa;
1704: douta=16'h6b2d;
1705: douta=16'h3a2a;
1706: douta=16'ha512;
1707: douta=16'h324d;
1708: douta=16'h32b0;
1709: douta=16'h5bb3;
1710: douta=16'h7496;
1711: douta=16'h5372;
1712: douta=16'h3ad0;
1713: douta=16'h4311;
1714: douta=16'h74b7;
1715: douta=16'h4bd6;
1716: douta=16'h5c37;
1717: douta=16'h5395;
1718: douta=16'h1949;
1719: douta=16'h53d5;
1720: douta=16'h7cb6;
1721: douta=16'h53f5;
1722: douta=16'h7433;
1723: douta=16'h42b0;
1724: douta=16'h2a0c;
1725: douta=16'h4b11;
1726: douta=16'h5b91;
1727: douta=16'ha578;
1728: douta=16'ha5d9;
1729: douta=16'h324e;
1730: douta=16'h42ae;
1731: douta=16'h5b71;
1732: douta=16'h2146;
1733: douta=16'h2966;
1734: douta=16'h18a4;
1735: douta=16'h7b6e;
1736: douta=16'h8cf8;
1737: douta=16'h8519;
1738: douta=16'h8d19;
1739: douta=16'h851a;
1740: douta=16'h8d3a;
1741: douta=16'h851a;
1742: douta=16'h8d3a;
1743: douta=16'h851a;
1744: douta=16'h7cd9;
1745: douta=16'h8d5b;
1746: douta=16'h7cd8;
1747: douta=16'h8d7b;
1748: douta=16'h851a;
1749: douta=16'h8d7b;
1750: douta=16'h7cf9;
1751: douta=16'h6cb9;
1752: douta=16'h5c17;
1753: douta=16'h6c99;
1754: douta=16'h6478;
1755: douta=16'h7d3b;
1756: douta=16'h6478;
1757: douta=16'h7d3a;
1758: douta=16'h859d;
1759: douta=16'h7d3a;
1760: douta=16'h8dbc;
1761: douta=16'h855a;
1762: douta=16'h855b;
1763: douta=16'h6c99;
1764: douta=16'h855a;
1765: douta=16'h7d1a;
1766: douta=16'h751a;
1767: douta=16'h7d1a;
1768: douta=16'h6457;
1769: douta=16'h751a;
1770: douta=16'h74d9;
1771: douta=16'h74d9;
1772: douta=16'h755c;
1773: douta=16'h751a;
1774: douta=16'h74da;
1775: douta=16'h29aa;
1776: douta=16'h10e5;
1777: douta=16'h1107;
1778: douta=16'h1106;
1779: douta=16'h42ee;
1780: douta=16'h73f2;
1781: douta=16'h19ab;
1782: douta=16'h326e;
1783: douta=16'h9d79;
1784: douta=16'h9d37;
1785: douta=16'h5c38;
1786: douta=16'h3b54;
1787: douta=16'h6c97;
1788: douta=16'hadba;
1789: douta=16'h6c57;
1790: douta=16'h2a4f;
1791: douta=16'h3b12;
1792: douta=16'h32d2;
1793: douta=16'h6c37;
1794: douta=16'h6c36;
1795: douta=16'h5bb4;
1796: douta=16'h5b73;
1797: douta=16'h7435;
1798: douta=16'h9517;
1799: douta=16'h7434;
1800: douta=16'h7413;
1801: douta=16'h5b92;
1802: douta=16'hd679;
1803: douta=16'hbdf8;
1804: douta=16'hc5f7;
1805: douta=16'ha515;
1806: douta=16'he6f9;
1807: douta=16'hc658;
1808: douta=16'hc5f7;
1809: douta=16'h8c51;
1810: douta=16'hde98;
1811: douta=16'hf71a;
1812: douta=16'h8452;
1813: douta=16'h8430;
1814: douta=16'hd6b8;
1815: douta=16'hf73a;
1816: douta=16'h638f;
1817: douta=16'h9512;
1818: douta=16'had73;
1819: douta=16'heeb7;
1820: douta=16'hb4b0;
1821: douta=16'hbd72;
1822: douta=16'ha46e;
1823: douta=16'h6b8d;
1824: douta=16'had11;
1825: douta=16'h634d;
1826: douta=16'h52aa;
1827: douta=16'h94b2;
1828: douta=16'hb5b4;
1829: douta=16'he6d7;
1830: douta=16'h738f;
1831: douta=16'h9c91;
1832: douta=16'h8c2e;
1833: douta=16'h18e4;
1834: douta=16'h4a8c;
1835: douta=16'h6bf2;
1836: douta=16'h0841;
1837: douta=16'h3a4d;
1838: douta=16'h29ec;
1839: douta=16'h5bd3;
1840: douta=16'h42af;
1841: douta=16'h2a2d;
1842: douta=16'h84d7;
1843: douta=16'h7c56;
1844: douta=16'h5395;
1845: douta=16'h4333;
1846: douta=16'h4b53;
1847: douta=16'h6456;
1848: douta=16'h6415;
1849: douta=16'h4352;
1850: douta=16'h8cd7;
1851: douta=16'h53b4;
1852: douta=16'h7454;
1853: douta=16'h8495;
1854: douta=16'h4b11;
1855: douta=16'h84b7;
1856: douta=16'h42ef;
1857: douta=16'h4af0;
1858: douta=16'h5b91;
1859: douta=16'h3167;
1860: douta=16'h1946;
1861: douta=16'h72aa;
1862: douta=16'h7c96;
1863: douta=16'h7477;
1864: douta=16'h7497;
1865: douta=16'h84f9;
1866: douta=16'h6415;
1867: douta=16'h957b;
1868: douta=16'h853b;
1869: douta=16'h8d3a;
1870: douta=16'h8d7b;
1871: douta=16'h8d3a;
1872: douta=16'h84f9;
1873: douta=16'h8d3a;
1874: douta=16'h853a;
1875: douta=16'h8d7b;
1876: douta=16'h957b;
1877: douta=16'h853a;
1878: douta=16'h855a;
1879: douta=16'h959b;
1880: douta=16'h957b;
1881: douta=16'h6cb9;
1882: douta=16'h751a;
1883: douta=16'h53f6;
1884: douta=16'h7d1b;
1885: douta=16'h859c;
1886: douta=16'h7d1a;
1887: douta=16'h5c37;
1888: douta=16'h855b;
1889: douta=16'h7d3a;
1890: douta=16'h855b;
1891: douta=16'h7d3a;
1892: douta=16'h7d3a;
1893: douta=16'h7d1a;
1894: douta=16'h74d9;
1895: douta=16'h7d1a;
1896: douta=16'h853b;
1897: douta=16'h74da;
1898: douta=16'h6cb9;
1899: douta=16'h7d5c;
1900: douta=16'h6c98;
1901: douta=16'h7d5c;
1902: douta=16'h6499;
1903: douta=16'h74fa;
1904: douta=16'h6436;
1905: douta=16'h29ca;
1906: douta=16'h08e5;
1907: douta=16'h1927;
1908: douta=16'h2a4e;
1909: douta=16'h4b51;
1910: douta=16'h84d6;
1911: douta=16'ha578;
1912: douta=16'h5bf5;
1913: douta=16'h2ab0;
1914: douta=16'hb63b;
1915: douta=16'h9579;
1916: douta=16'h6478;
1917: douta=16'h5395;
1918: douta=16'h6c77;
1919: douta=16'h6458;
1920: douta=16'h5416;
1921: douta=16'h7457;
1922: douta=16'h6416;
1923: douta=16'h5373;
1924: douta=16'h5372;
1925: douta=16'h7455;
1926: douta=16'ha599;
1927: douta=16'h73f3;
1928: douta=16'h8494;
1929: douta=16'h9d56;
1930: douta=16'hb597;
1931: douta=16'ha557;
1932: douta=16'hce58;
1933: douta=16'hc5f7;
1934: douta=16'hce17;
1935: douta=16'hb575;
1936: douta=16'ha4d4;
1937: douta=16'hbdb5;
1938: douta=16'hce57;
1939: douta=16'hde98;
1940: douta=16'hb532;
1941: douta=16'h73f0;
1942: douta=16'hde98;
1943: douta=16'hef19;
1944: douta=16'h426a;
1945: douta=16'hd655;
1946: douta=16'he6d7;
1947: douta=16'hff38;
1948: douta=16'h6aca;
1949: douta=16'hb510;
1950: douta=16'h946f;
1951: douta=16'h62cb;
1952: douta=16'h2127;
1953: douta=16'h18e5;
1954: douta=16'h0043;
1955: douta=16'h73ae;
1956: douta=16'h7410;
1957: douta=16'had32;
1958: douta=16'h8c50;
1959: douta=16'h9cb0;
1960: douta=16'hde97;
1961: douta=16'h5b4e;
1962: douta=16'h63d3;
1963: douta=16'h4a4b;
1964: douta=16'h18a2;
1965: douta=16'h1082;
1966: douta=16'h1882;
1967: douta=16'h3aaf;
1968: douta=16'h0907;
1969: douta=16'h5393;
1970: douta=16'h6477;
1971: douta=16'h6c56;
1972: douta=16'h5b93;
1973: douta=16'h4b53;
1974: douta=16'h63f5;
1975: douta=16'h6bf2;
1976: douta=16'h4acf;
1977: douta=16'h5352;
1978: douta=16'h42f1;
1979: douta=16'h32b1;
1980: douta=16'h6c56;
1981: douta=16'h63d3;
1982: douta=16'h9d57;
1983: douta=16'ha599;
1984: douta=16'h7413;
1985: douta=16'h4aad;
1986: douta=16'h31c7;
1987: douta=16'h41a6;
1988: douta=16'h8c52;
1989: douta=16'h84f8;
1990: douta=16'h84f8;
1991: douta=16'h7c97;
1992: douta=16'h8d39;
1993: douta=16'h84f9;
1994: douta=16'h7cb8;
1995: douta=16'h84f9;
1996: douta=16'h5373;
1997: douta=16'h8d7b;
1998: douta=16'h959b;
1999: douta=16'h8d5a;
2000: douta=16'h7477;
2001: douta=16'h84d9;
2002: douta=16'h959b;
2003: douta=16'h8d5b;
2004: douta=16'h853a;
2005: douta=16'h74b8;
2006: douta=16'h8d7b;
2007: douta=16'h957b;
2008: douta=16'h8d7b;
2009: douta=16'h95bc;
2010: douta=16'h959c;
2011: douta=16'h74da;
2012: douta=16'h5c58;
2013: douta=16'h859c;
2014: douta=16'h4b76;
2015: douta=16'h8dbc;
2016: douta=16'h74da;
2017: douta=16'h855b;
2018: douta=16'h7d3a;
2019: douta=16'h859c;
2020: douta=16'h855b;
2021: douta=16'h7d3b;
2022: douta=16'h5c17;
2023: douta=16'h8d9b;
2024: douta=16'h7d3a;
2025: douta=16'h7d3a;
2026: douta=16'h7d3b;
2027: douta=16'h753a;
2028: douta=16'h8d9b;
2029: douta=16'h7d7c;
2030: douta=16'h6458;
2031: douta=16'h74fa;
2032: douta=16'h6d1a;
2033: douta=16'h753b;
2034: douta=16'h42cf;
2035: douta=16'h21a8;
2036: douta=16'h1927;
2037: douta=16'h32af;
2038: douta=16'h8c94;
2039: douta=16'h63f5;
2040: douta=16'h3ab0;
2041: douta=16'haddb;
2042: douta=16'h63d4;
2043: douta=16'h2a90;
2044: douta=16'h4395;
2045: douta=16'h8518;
2046: douta=16'h9dbb;
2047: douta=16'h8d5a;
2048: douta=16'h53f6;
2049: douta=16'h5374;
2050: douta=16'h5bb4;
2051: douta=16'h6436;
2052: douta=16'h5b93;
2053: douta=16'h7c76;
2054: douta=16'hc5f9;
2055: douta=16'h7c74;
2056: douta=16'h6bd2;
2057: douta=16'h73f3;
2058: douta=16'ha4d4;
2059: douta=16'ha4f5;
2060: douta=16'hb596;
2061: douta=16'hbdb6;
2062: douta=16'heef9;
2063: douta=16'ha4d3;
2064: douta=16'ha4d3;
2065: douta=16'hde98;
2066: douta=16'hcdf6;
2067: douta=16'hd637;
2068: douta=16'ha4d2;
2069: douta=16'hc5d4;
2070: douta=16'h9cd1;
2071: douta=16'hd696;
2072: douta=16'h634d;
2073: douta=16'hb593;
2074: douta=16'hbdd3;
2075: douta=16'heeb7;
2076: douta=16'h7b4b;
2077: douta=16'h6b0b;
2078: douta=16'h5289;
2079: douta=16'h4a29;
2080: douta=16'h18e5;
2081: douta=16'h2146;
2082: douta=16'h10e4;
2083: douta=16'h1043;
2084: douta=16'h5b0e;
2085: douta=16'ha513;
2086: douta=16'h9450;
2087: douta=16'hbdf5;
2088: douta=16'h8c50;
2089: douta=16'h4b10;
2090: douta=16'h428d;
2091: douta=16'h52ee;
2092: douta=16'h3b11;
2093: douta=16'h0000;
2094: douta=16'h18e3;
2095: douta=16'h10c2;
2096: douta=16'h29a8;
2097: douta=16'h1127;
2098: douta=16'h32f0;
2099: douta=16'h53b4;
2100: douta=16'h19cc;
2101: douta=16'h53b4;
2102: douta=16'h42f1;
2103: douta=16'h7d19;
2104: douta=16'h5c14;
2105: douta=16'h426d;
2106: douta=16'h4b53;
2107: douta=16'h4b53;
2108: douta=16'h7c97;
2109: douta=16'h4b31;
2110: douta=16'h6c34;
2111: douta=16'h3a8f;
2112: douta=16'h4aac;
2113: douta=16'h29a8;
2114: douta=16'hac0e;
2115: douta=16'h94f7;
2116: douta=16'h8d19;
2117: douta=16'h6c15;
2118: douta=16'h84b7;
2119: douta=16'h6c15;
2120: douta=16'h8d39;
2121: douta=16'h957a;
2122: douta=16'h8d5a;
2123: douta=16'h7cd8;
2124: douta=16'h8d3a;
2125: douta=16'h84d8;
2126: douta=16'h7477;
2127: douta=16'h957b;
2128: douta=16'h853a;
2129: douta=16'h7cb8;
2130: douta=16'h8d5b;
2131: douta=16'h851a;
2132: douta=16'h855a;
2133: douta=16'h853a;
2134: douta=16'h8d5a;
2135: douta=16'h8d7b;
2136: douta=16'h8d5a;
2137: douta=16'h8d7b;
2138: douta=16'h8d3a;
2139: douta=16'h8d9b;
2140: douta=16'h8d9b;
2141: douta=16'h6cb9;
2142: douta=16'h5c37;
2143: douta=16'h6c99;
2144: douta=16'h7d7c;
2145: douta=16'h753b;
2146: douta=16'h6cb9;
2147: douta=16'h855a;
2148: douta=16'h8d9c;
2149: douta=16'h751a;
2150: douta=16'h859c;
2151: douta=16'h7d1b;
2152: douta=16'h74d9;
2153: douta=16'h859c;
2154: douta=16'h859c;
2155: douta=16'h6cda;
2156: douta=16'h751a;
2157: douta=16'h6cb9;
2158: douta=16'h8d9b;
2159: douta=16'h5bd6;
2160: douta=16'h7d7c;
2161: douta=16'h6cb9;
2162: douta=16'h6d1a;
2163: douta=16'h857b;
2164: douta=16'h21a9;
2165: douta=16'h1948;
2166: douta=16'h2a2d;
2167: douta=16'h220e;
2168: douta=16'h5393;
2169: douta=16'h6c36;
2170: douta=16'h3b34;
2171: douta=16'h53d5;
2172: douta=16'h7c96;
2173: douta=16'hcefe;
2174: douta=16'h5c16;
2175: douta=16'h4b95;
2176: douta=16'h4375;
2177: douta=16'h4312;
2178: douta=16'h6c78;
2179: douta=16'h2a70;
2180: douta=16'h5b73;
2181: douta=16'h6bd4;
2182: douta=16'h7c33;
2183: douta=16'h6bd2;
2184: douta=16'h6350;
2185: douta=16'h8c94;
2186: douta=16'h9cd4;
2187: douta=16'h8453;
2188: douta=16'had55;
2189: douta=16'hd657;
2190: douta=16'hdeb9;
2191: douta=16'ha4d2;
2192: douta=16'h9cd3;
2193: douta=16'hf738;
2194: douta=16'hc5d5;
2195: douta=16'hc5b5;
2196: douta=16'hcdf5;
2197: douta=16'hde76;
2198: douta=16'ha48f;
2199: douta=16'hce16;
2200: douta=16'h6b4d;
2201: douta=16'hb551;
2202: douta=16'hc5d3;
2203: douta=16'hde96;
2204: douta=16'h7b4b;
2205: douta=16'h62ca;
2206: douta=16'h31a7;
2207: douta=16'h2167;
2208: douta=16'h31e9;
2209: douta=16'h2988;
2210: douta=16'h10e4;
2211: douta=16'h0084;
2212: douta=16'h4aac;
2213: douta=16'h530c;
2214: douta=16'h840f;
2215: douta=16'h7bce;
2216: douta=16'h6c34;
2217: douta=16'h4b31;
2218: douta=16'h29c9;
2219: douta=16'h9472;
2220: douta=16'h4331;
2221: douta=16'h4b0f;
2222: douta=16'h3a0c;
2223: douta=16'h1061;
2224: douta=16'h18e4;
2225: douta=16'h1061;
2226: douta=16'h5bb4;
2227: douta=16'h00e7;
2228: douta=16'h32d1;
2229: douta=16'h3b31;
2230: douta=16'h4b73;
2231: douta=16'h29ec;
2232: douta=16'h216a;
2233: douta=16'h4b31;
2234: douta=16'h6477;
2235: douta=16'h74b8;
2236: douta=16'h74f9;
2237: douta=16'h6bd2;
2238: douta=16'h21cc;
2239: douta=16'h52f0;
2240: douta=16'h4229;
2241: douta=16'h836c;
2242: douta=16'h84d8;
2243: douta=16'h9d9a;
2244: douta=16'h7435;
2245: douta=16'h9519;
2246: douta=16'h84f8;
2247: douta=16'h7456;
2248: douta=16'h8d18;
2249: douta=16'h84d8;
2250: douta=16'h7cb8;
2251: douta=16'h84f9;
2252: douta=16'h6c56;
2253: douta=16'h8d3a;
2254: douta=16'h7cd8;
2255: douta=16'h8519;
2256: douta=16'h8519;
2257: douta=16'h7cb9;
2258: douta=16'h853a;
2259: douta=16'h8d7b;
2260: douta=16'h853a;
2261: douta=16'h853a;
2262: douta=16'h8d9b;
2263: douta=16'h959c;
2264: douta=16'h853a;
2265: douta=16'h8d7a;
2266: douta=16'h959b;
2267: douta=16'h8519;
2268: douta=16'h8d5a;
2269: douta=16'h851a;
2270: douta=16'h959c;
2271: douta=16'h853a;
2272: douta=16'h6458;
2273: douta=16'h74fa;
2274: douta=16'h64b9;
2275: douta=16'h7d7b;
2276: douta=16'h8dfd;
2277: douta=16'h8dbd;
2278: douta=16'h7d5b;
2279: douta=16'h95bc;
2280: douta=16'h7d3b;
2281: douta=16'h7d3a;
2282: douta=16'h857c;
2283: douta=16'h74fa;
2284: douta=16'h8d9b;
2285: douta=16'h6499;
2286: douta=16'h7d5a;
2287: douta=16'h74d9;
2288: douta=16'h7d3a;
2289: douta=16'h5c16;
2290: douta=16'h7d7b;
2291: douta=16'h6cb9;
2292: douta=16'h7cfa;
2293: douta=16'h29a8;
2294: douta=16'h1968;
2295: douta=16'h53d4;
2296: douta=16'hb61b;
2297: douta=16'h5c16;
2298: douta=16'h220d;
2299: douta=16'h5392;
2300: douta=16'hbe3b;
2301: douta=16'h7456;
2302: douta=16'h6c77;
2303: douta=16'h84d7;
2304: douta=16'h4bf6;
2305: douta=16'h5416;
2306: douta=16'h5c16;
2307: douta=16'h32b1;
2308: douta=16'h6c14;
2309: douta=16'h8d18;
2310: douta=16'h5b30;
2311: douta=16'h7c53;
2312: douta=16'h8c53;
2313: douta=16'hb5f9;
2314: douta=16'hce17;
2315: douta=16'h9494;
2316: douta=16'h94b3;
2317: douta=16'hc5f6;
2318: douta=16'ha4f4;
2319: douta=16'hbdb6;
2320: douta=16'hb533;
2321: douta=16'hde77;
2322: douta=16'hc5f5;
2323: douta=16'hbdb5;
2324: douta=16'had11;
2325: douta=16'had11;
2326: douta=16'hb531;
2327: douta=16'heef9;
2328: douta=16'h630c;
2329: douta=16'hc5f4;
2330: douta=16'hb532;
2331: douta=16'h83ed;
2332: douta=16'h7b4b;
2333: douta=16'h62ca;
2334: douta=16'h4a27;
2335: douta=16'h10a4;
2336: douta=16'h18e5;
2337: douta=16'h1105;
2338: douta=16'h2167;
2339: douta=16'h10e5;
2340: douta=16'h62aa;
2341: douta=16'h4a4a;
2342: douta=16'h9cf2;
2343: douta=16'h63b2;
2344: douta=16'h532f;
2345: douta=16'h8c72;
2346: douta=16'h7c30;
2347: douta=16'h840f;
2348: douta=16'h52ac;
2349: douta=16'h63b1;
2350: douta=16'h42ce;
2351: douta=16'h63d1;
2352: douta=16'h3a6b;
2353: douta=16'h1082;
2354: douta=16'h0040;
2355: douta=16'h1925;
2356: douta=16'h19ab;
2357: douta=16'h328f;
2358: douta=16'h53f5;
2359: douta=16'h324e;
2360: douta=16'h21ec;
2361: douta=16'h32af;
2362: douta=16'h4374;
2363: douta=16'h853a;
2364: douta=16'h224f;
2365: douta=16'h6415;
2366: douta=16'h5b93;
2367: douta=16'h3a4a;
2368: douta=16'ha44f;
2369: douta=16'h7cb7;
2370: douta=16'h959a;
2371: douta=16'h5b93;
2372: douta=16'h8d5a;
2373: douta=16'h957b;
2374: douta=16'h7c96;
2375: douta=16'h84b8;
2376: douta=16'h9559;
2377: douta=16'h6c56;
2378: douta=16'h7c97;
2379: douta=16'h8519;
2380: douta=16'h7cb8;
2381: douta=16'h8d7a;
2382: douta=16'h7c98;
2383: douta=16'h6c56;
2384: douta=16'h6c36;
2385: douta=16'h7cd9;
2386: douta=16'h8d7b;
2387: douta=16'h959b;
2388: douta=16'h8d5a;
2389: douta=16'h7498;
2390: douta=16'h959b;
2391: douta=16'h8d5b;
2392: douta=16'h959b;
2393: douta=16'h84f9;
2394: douta=16'h95bc;
2395: douta=16'h959b;
2396: douta=16'h959b;
2397: douta=16'h8d5a;
2398: douta=16'h851a;
2399: douta=16'h95bc;
2400: douta=16'h95bc;
2401: douta=16'h853b;
2402: douta=16'h74da;
2403: douta=16'h7d5b;
2404: douta=16'h6cda;
2405: douta=16'h85bd;
2406: douta=16'h753a;
2407: douta=16'h8ddc;
2408: douta=16'h7d5b;
2409: douta=16'h7d3b;
2410: douta=16'h7d5b;
2411: douta=16'h751a;
2412: douta=16'h857b;
2413: douta=16'h6498;
2414: douta=16'h7d5b;
2415: douta=16'h74b9;
2416: douta=16'h74b9;
2417: douta=16'h8d9c;
2418: douta=16'h6498;
2419: douta=16'h6cda;
2420: douta=16'h7d7b;
2421: douta=16'h6cba;
2422: douta=16'h2167;
2423: douta=16'h21a9;
2424: douta=16'h7477;
2425: douta=16'h32d2;
2426: douta=16'h5bb4;
2427: douta=16'hadba;
2428: douta=16'h5bb4;
2429: douta=16'h3290;
2430: douta=16'h32b0;
2431: douta=16'h7c75;
2432: douta=16'h32d2;
2433: douta=16'h5c57;
2434: douta=16'h4b32;
2435: douta=16'h5bd5;
2436: douta=16'h7c56;
2437: douta=16'h9d59;
2438: douta=16'h7c12;
2439: douta=16'h5b70;
2440: douta=16'ha516;
2441: douta=16'hce39;
2442: douta=16'ha515;
2443: douta=16'had35;
2444: douta=16'h8c52;
2445: douta=16'hde77;
2446: douta=16'h8c72;
2447: douta=16'h6b4d;
2448: douta=16'h8410;
2449: douta=16'hde76;
2450: douta=16'had33;
2451: douta=16'h52ed;
2452: douta=16'h9c90;
2453: douta=16'hbdd3;
2454: douta=16'hcdd3;
2455: douta=16'hd636;
2456: douta=16'h842e;
2457: douta=16'hc614;
2458: douta=16'h7b6c;
2459: douta=16'h83ac;
2460: douta=16'h7b4b;
2461: douta=16'h62a9;
2462: douta=16'h4a49;
2463: douta=16'h2167;
2464: douta=16'h39a7;
2465: douta=16'h10e5;
2466: douta=16'h10e4;
2467: douta=16'h18e5;
2468: douta=16'h4229;
2469: douta=16'h39a8;
2470: douta=16'h738d;
2471: douta=16'h63d2;
2472: douta=16'h5b0e;
2473: douta=16'h1927;
2474: douta=16'h530d;
2475: douta=16'h8430;
2476: douta=16'h7bef;
2477: douta=16'h8474;
2478: douta=16'h7c33;
2479: douta=16'h5370;
2480: douta=16'h4b10;
2481: douta=16'h5393;
2482: douta=16'h0841;
2483: douta=16'h10e3;
2484: douta=16'h1060;
2485: douta=16'h428d;
2486: douta=16'h220c;
2487: douta=16'h4374;
2488: douta=16'h29ec;
2489: douta=16'h3b11;
2490: douta=16'h4373;
2491: douta=16'h53b4;
2492: douta=16'h198b;
2493: douta=16'h6498;
2494: douta=16'h4a4a;
2495: douta=16'hacaf;
2496: douta=16'h95bc;
2497: douta=16'h6478;
2498: douta=16'h7cd8;
2499: douta=16'h957a;
2500: douta=16'h6416;
2501: douta=16'h5bb5;
2502: douta=16'h7457;
2503: douta=16'h7c76;
2504: douta=16'h7cb8;
2505: douta=16'h6c36;
2506: douta=16'h6415;
2507: douta=16'h8d1a;
2508: douta=16'h84f9;
2509: douta=16'h959b;
2510: douta=16'h7477;
2511: douta=16'h7cb8;
2512: douta=16'h7497;
2513: douta=16'h6c56;
2514: douta=16'h7478;
2515: douta=16'h851a;
2516: douta=16'h7cd8;
2517: douta=16'h8d7a;
2518: douta=16'h8d3b;
2519: douta=16'h7cd9;
2520: douta=16'h959c;
2521: douta=16'h8d5a;
2522: douta=16'h7d19;
2523: douta=16'h8d3a;
2524: douta=16'h851a;
2525: douta=16'h8d3a;
2526: douta=16'h853a;
2527: douta=16'h8d5b;
2528: douta=16'h7cf9;
2529: douta=16'h851a;
2530: douta=16'h8d7b;
2531: douta=16'h855a;
2532: douta=16'h6499;
2533: douta=16'h8e1e;
2534: douta=16'h6478;
2535: douta=16'h6cfa;
2536: douta=16'h74da;
2537: douta=16'h857c;
2538: douta=16'h751a;
2539: douta=16'h857b;
2540: douta=16'h74d9;
2541: douta=16'h74fa;
2542: douta=16'h751a;
2543: douta=16'h6458;
2544: douta=16'h859b;
2545: douta=16'h8d5b;
2546: douta=16'h6c98;
2547: douta=16'h6cfa;
2548: douta=16'h6478;
2549: douta=16'h74fa;
2550: douta=16'h751b;
2551: douta=16'h1906;
2552: douta=16'h1107;
2553: douta=16'h5353;
2554: douta=16'h7497;
2555: douta=16'h19cc;
2556: douta=16'h32d0;
2557: douta=16'h4b51;
2558: douta=16'h7c75;
2559: douta=16'h42d0;
2560: douta=16'h4353;
2561: douta=16'h6c99;
2562: douta=16'h324f;
2563: douta=16'h4311;
2564: douta=16'h6bd4;
2565: douta=16'h84d7;
2566: douta=16'h530f;
2567: douta=16'h530f;
2568: douta=16'hbd96;
2569: douta=16'hd69a;
2570: douta=16'h9c94;
2571: douta=16'h6b8f;
2572: douta=16'hbd95;
2573: douta=16'hde78;
2574: douta=16'h9cb3;
2575: douta=16'h7bae;
2576: douta=16'h632d;
2577: douta=16'hb573;
2578: douta=16'hacf2;
2579: douta=16'h9491;
2580: douta=16'h83ed;
2581: douta=16'hb572;
2582: douta=16'hbd93;
2583: douta=16'hdeb7;
2584: douta=16'h944e;
2585: douta=16'h838b;
2586: douta=16'h8bac;
2587: douta=16'h8bcb;
2588: douta=16'h93ec;
2589: douta=16'h62a9;
2590: douta=16'h2147;
2591: douta=16'h2946;
2592: douta=16'h2126;
2593: douta=16'h10a4;
2594: douta=16'h10e5;
2595: douta=16'h10e4;
2596: douta=16'h10a4;
2597: douta=16'h528a;
2598: douta=16'h8c2e;
2599: douta=16'h5b71;
2600: douta=16'h322b;
2601: douta=16'h1988;
2602: douta=16'h426b;
2603: douta=16'h4acd;
2604: douta=16'h9cf3;
2605: douta=16'h08c6;
2606: douta=16'h6bb1;
2607: douta=16'h4b0f;
2608: douta=16'h5b71;
2609: douta=16'h5bb2;
2610: douta=16'h2a0c;
2611: douta=16'h5b70;
2612: douta=16'h10c2;
2613: douta=16'h10c4;
2614: douta=16'h0000;
2615: douta=16'h320c;
2616: douta=16'h32af;
2617: douta=16'h3333;
2618: douta=16'h6415;
2619: douta=16'h5394;
2620: douta=16'h4310;
2621: douta=16'h5a6a;
2622: douta=16'hc54f;
2623: douta=16'hae5e;
2624: douta=16'h959b;
2625: douta=16'h959b;
2626: douta=16'h8519;
2627: douta=16'h957a;
2628: douta=16'h959c;
2629: douta=16'h959b;
2630: douta=16'h7cf8;
2631: douta=16'h7cd8;
2632: douta=16'h7498;
2633: douta=16'h7cb8;
2634: douta=16'h7478;
2635: douta=16'h84d9;
2636: douta=16'h851a;
2637: douta=16'h957a;
2638: douta=16'h6c35;
2639: douta=16'h8d5a;
2640: douta=16'h7cd8;
2641: douta=16'h8d3a;
2642: douta=16'h84f9;
2643: douta=16'h6435;
2644: douta=16'h6c16;
2645: douta=16'h7477;
2646: douta=16'h9ddc;
2647: douta=16'h7cf9;
2648: douta=16'h959c;
2649: douta=16'h853a;
2650: douta=16'h855a;
2651: douta=16'h95bc;
2652: douta=16'h8519;
2653: douta=16'h8519;
2654: douta=16'h8d5a;
2655: douta=16'h959b;
2656: douta=16'h8d5b;
2657: douta=16'h8d5a;
2658: douta=16'h853b;
2659: douta=16'h959c;
2660: douta=16'h855b;
2661: douta=16'h959c;
2662: douta=16'h1a2f;
2663: douta=16'h85bd;
2664: douta=16'h6cda;
2665: douta=16'h6c99;
2666: douta=16'h74fa;
2667: douta=16'h751a;
2668: douta=16'h855b;
2669: douta=16'h855b;
2670: douta=16'h6cd9;
2671: douta=16'h7d3a;
2672: douta=16'h7d3a;
2673: douta=16'h7d3a;
2674: douta=16'h857b;
2675: douta=16'h95bc;
2676: douta=16'h6c99;
2677: douta=16'h74da;
2678: douta=16'h6c57;
2679: douta=16'h7498;
2680: douta=16'h2168;
2681: douta=16'ha5fc;
2682: douta=16'h63f4;
2683: douta=16'h7496;
2684: douta=16'hb5f8;
2685: douta=16'h7c33;
2686: douta=16'h6416;
2687: douta=16'h324e;
2688: douta=16'h3b33;
2689: douta=16'h4333;
2690: douta=16'h42d1;
2691: douta=16'h322e;
2692: douta=16'h63d3;
2693: douta=16'h84b7;
2694: douta=16'h6392;
2695: douta=16'h7c35;
2696: douta=16'h9cd6;
2697: douta=16'hd69b;
2698: douta=16'h94b4;
2699: douta=16'hbd95;
2700: douta=16'hd657;
2701: douta=16'hde97;
2702: douta=16'hb574;
2703: douta=16'h5aed;
2704: douta=16'h7bcf;
2705: douta=16'hbd94;
2706: douta=16'h940f;
2707: douta=16'h8c4f;
2708: douta=16'h62c9;
2709: douta=16'hb530;
2710: douta=16'hb592;
2711: douta=16'hbd93;
2712: douta=16'h7b2b;
2713: douta=16'h8bcc;
2714: douta=16'h93cc;
2715: douta=16'h9c0d;
2716: douta=16'h9c0d;
2717: douta=16'h6aea;
2718: douta=16'h2125;
2719: douta=16'h2987;
2720: douta=16'h1905;
2721: douta=16'h1926;
2722: douta=16'h18e5;
2723: douta=16'h18e5;
2724: douta=16'h1105;
2725: douta=16'hacd0;
2726: douta=16'h0000;
2727: douta=16'h5b90;
2728: douta=16'h2147;
2729: douta=16'h634d;
2730: douta=16'h3209;
2731: douta=16'h29a9;
2732: douta=16'h3a4c;
2733: douta=16'h1106;
2734: douta=16'h5b2e;
2735: douta=16'h29cb;
2736: douta=16'h2a0c;
2737: douta=16'h3b10;
2738: douta=16'h3acf;
2739: douta=16'h42f1;
2740: douta=16'h5bf5;
2741: douta=16'h4acd;
2742: douta=16'h0861;
2743: douta=16'h0820;
2744: douta=16'h31ea;
2745: douta=16'h3a8f;
2746: douta=16'h5bf5;
2747: douta=16'h5c36;
2748: douta=16'h524a;
2749: douta=16'hd550;
2750: douta=16'h8d18;
2751: douta=16'h5375;
2752: douta=16'h8d9b;
2753: douta=16'h853a;
2754: douta=16'h8d7b;
2755: douta=16'hae1c;
2756: douta=16'h959b;
2757: douta=16'h853a;
2758: douta=16'h959b;
2759: douta=16'ha5db;
2760: douta=16'h7478;
2761: douta=16'h7cb8;
2762: douta=16'h855a;
2763: douta=16'h9dbb;
2764: douta=16'h851a;
2765: douta=16'h7cd9;
2766: douta=16'h7cd8;
2767: douta=16'h9ddb;
2768: douta=16'h6c15;
2769: douta=16'h957a;
2770: douta=16'h6c16;
2771: douta=16'h7cd8;
2772: douta=16'h8d5a;
2773: douta=16'h74b8;
2774: douta=16'h7cd9;
2775: douta=16'h7cb8;
2776: douta=16'h8d5b;
2777: douta=16'h6c36;
2778: douta=16'h7cf9;
2779: douta=16'h8d5b;
2780: douta=16'h853a;
2781: douta=16'h95bc;
2782: douta=16'h853a;
2783: douta=16'h959c;
2784: douta=16'h8d5b;
2785: douta=16'h959b;
2786: douta=16'h95bc;
2787: douta=16'h8d7b;
2788: douta=16'h853a;
2789: douta=16'h857b;
2790: douta=16'h851a;
2791: douta=16'h95bd;
2792: douta=16'h74d9;
2793: douta=16'h857b;
2794: douta=16'h53f6;
2795: douta=16'h751b;
2796: douta=16'h6498;
2797: douta=16'h751b;
2798: douta=16'h859c;
2799: douta=16'h6cb9;
2800: douta=16'h6c79;
2801: douta=16'h7d5a;
2802: douta=16'h859b;
2803: douta=16'h8d7b;
2804: douta=16'h74f9;
2805: douta=16'h857b;
2806: douta=16'h74da;
2807: douta=16'h74fa;
2808: douta=16'h6415;
2809: douta=16'h2189;
2810: douta=16'h8cd5;
2811: douta=16'h8cf5;
2812: douta=16'h6391;
2813: douta=16'h63b2;
2814: douta=16'h5b91;
2815: douta=16'h8453;
2816: douta=16'h32f2;
2817: douta=16'h4354;
2818: douta=16'h4b52;
2819: douta=16'h5bb4;
2820: douta=16'h5b72;
2821: douta=16'h84b7;
2822: douta=16'h5b31;
2823: douta=16'h6bb2;
2824: douta=16'ha537;
2825: douta=16'hc5d7;
2826: douta=16'h8432;
2827: douta=16'h7c12;
2828: douta=16'h8410;
2829: douta=16'ha534;
2830: douta=16'hb553;
2831: douta=16'h632d;
2832: douta=16'h632d;
2833: douta=16'h942f;
2834: douta=16'ha4d0;
2835: douta=16'h9490;
2836: douta=16'h942d;
2837: douta=16'hacf0;
2838: douta=16'hce34;
2839: douta=16'h736b;
2840: douta=16'h7b6b;
2841: douta=16'h9c0c;
2842: douta=16'h9c0c;
2843: douta=16'h9c2d;
2844: douta=16'hb4ad;
2845: douta=16'h836c;
2846: douta=16'h838c;
2847: douta=16'h5249;
2848: douta=16'h1905;
2849: douta=16'h1926;
2850: douta=16'h1905;
2851: douta=16'h10e5;
2852: douta=16'h1905;
2853: douta=16'h10c3;
2854: douta=16'h0000;
2855: douta=16'h6c14;
2856: douta=16'h4249;
2857: douta=16'h5aeb;
2858: douta=16'h7bce;
2859: douta=16'h31ca;
2860: douta=16'h29ea;
2861: douta=16'h320a;
2862: douta=16'h3a4a;
2863: douta=16'h52cc;
2864: douta=16'h29aa;
2865: douta=16'h322c;
2866: douta=16'h73d1;
2867: douta=16'h5351;
2868: douta=16'h326e;
2869: douta=16'h3ad1;
2870: douta=16'h328e;
2871: douta=16'h18c3;
2872: douta=16'h20e4;
2873: douta=16'h1061;
2874: douta=16'h5350;
2875: douta=16'h220c;
2876: douta=16'h7289;
2877: douta=16'h5b0f;
2878: douta=16'h959a;
2879: douta=16'h8d39;
2880: douta=16'h8d7b;
2881: douta=16'h851a;
2882: douta=16'h53d6;
2883: douta=16'h74d9;
2884: douta=16'hae1c;
2885: douta=16'h95bb;
2886: douta=16'h959b;
2887: douta=16'h8539;
2888: douta=16'h7476;
2889: douta=16'h9d9a;
2890: douta=16'h5311;
2891: douta=16'h851a;
2892: douta=16'h8d7a;
2893: douta=16'h8d5a;
2894: douta=16'h84f9;
2895: douta=16'h8d7a;
2896: douta=16'h7497;
2897: douta=16'h8d3a;
2898: douta=16'h84f9;
2899: douta=16'h63d4;
2900: douta=16'h959a;
2901: douta=16'h7cd8;
2902: douta=16'h851a;
2903: douta=16'h855a;
2904: douta=16'h7cd8;
2905: douta=16'h6c57;
2906: douta=16'h851a;
2907: douta=16'h5bd5;
2908: douta=16'h851a;
2909: douta=16'h959b;
2910: douta=16'h7cf9;
2911: douta=16'h8d7b;
2912: douta=16'h7cd9;
2913: douta=16'h95bc;
2914: douta=16'h851a;
2915: douta=16'h8d5a;
2916: douta=16'h95dc;
2917: douta=16'h8d7b;
2918: douta=16'h853a;
2919: douta=16'h7cf9;
2920: douta=16'h8d5b;
2921: douta=16'h8d9b;
2922: douta=16'h7d1a;
2923: douta=16'h6498;
2924: douta=16'h6cb9;
2925: douta=16'h7d5b;
2926: douta=16'h6c99;
2927: douta=16'h6cd9;
2928: douta=16'h859c;
2929: douta=16'h7d5b;
2930: douta=16'h6cda;
2931: douta=16'h74ba;
2932: douta=16'h855b;
2933: douta=16'h95dc;
2934: douta=16'h5c17;
2935: douta=16'h7d1a;
2936: douta=16'h74f9;
2937: douta=16'h2988;
2938: douta=16'h7c74;
2939: douta=16'h6c35;
2940: douta=16'h4b11;
2941: douta=16'h32b0;
2942: douta=16'ha598;
2943: douta=16'h5310;
2944: douta=16'h3b54;
2945: douta=16'h4b95;
2946: douta=16'h3ab0;
2947: douta=16'h2a2e;
2948: douta=16'h7cb7;
2949: douta=16'h7c76;
2950: douta=16'h7414;
2951: douta=16'h8cb5;
2952: douta=16'h6bd3;
2953: douta=16'h9c93;
2954: douta=16'ha4d4;
2955: douta=16'h39eb;
2956: douta=16'h8451;
2957: douta=16'h9470;
2958: douta=16'hbd73;
2959: douta=16'h9450;
2960: douta=16'h5acb;
2961: douta=16'ha4d0;
2962: douta=16'h9c6f;
2963: douta=16'hb572;
2964: douta=16'h83ad;
2965: douta=16'hce34;
2966: douta=16'ha4f1;
2967: douta=16'h8bac;
2968: douta=16'h93cb;
2969: douta=16'h9c0c;
2970: douta=16'ha44c;
2971: douta=16'hb4ad;
2972: douta=16'hac8d;
2973: douta=16'hac6d;
2974: douta=16'h6aea;
2975: douta=16'h6b0a;
2976: douta=16'h39c8;
2977: douta=16'h18e5;
2978: douta=16'h18e5;
2979: douta=16'h1905;
2980: douta=16'h1905;
2981: douta=16'h0883;
2982: douta=16'h0002;
2983: douta=16'h84b6;
2984: douta=16'h3186;
2985: douta=16'h4229;
2986: douta=16'h630b;
2987: douta=16'h632d;
2988: douta=16'h422a;
2989: douta=16'h428c;
2990: douta=16'h5b0d;
2991: douta=16'h6b6f;
2992: douta=16'h2189;
2993: douta=16'h1927;
2994: douta=16'h636f;
2995: douta=16'h6bd2;
2996: douta=16'h5372;
2997: douta=16'h328f;
2998: douta=16'h1969;
2999: douta=16'h3a4b;
3000: douta=16'h532f;
3001: douta=16'h18c3;
3002: douta=16'h10c2;
3003: douta=16'h0860;
3004: douta=16'h5269;
3005: douta=16'h9579;
3006: douta=16'h959a;
3007: douta=16'h7cd7;
3008: douta=16'h7c98;
3009: douta=16'h8d5a;
3010: douta=16'h63d5;
3011: douta=16'h84f9;
3012: douta=16'h7cf8;
3013: douta=16'h7cd9;
3014: douta=16'ha5db;
3015: douta=16'h8519;
3016: douta=16'h7c97;
3017: douta=16'h84b8;
3018: douta=16'ha5ba;
3019: douta=16'ha5fc;
3020: douta=16'hae1c;
3021: douta=16'h957a;
3022: douta=16'h957a;
3023: douta=16'h84f9;
3024: douta=16'h7cf9;
3025: douta=16'h8d5a;
3026: douta=16'h7cd8;
3027: douta=16'h8d3a;
3028: douta=16'h95bb;
3029: douta=16'h7477;
3030: douta=16'h8d39;
3031: douta=16'h8d5a;
3032: douta=16'h8519;
3033: douta=16'h6c15;
3034: douta=16'h6c57;
3035: douta=16'h8d3a;
3036: douta=16'h8d5a;
3037: douta=16'h853a;
3038: douta=16'h6c16;
3039: douta=16'h7cf9;
3040: douta=16'h851a;
3041: douta=16'h957b;
3042: douta=16'h8d7b;
3043: douta=16'h851a;
3044: douta=16'h95bc;
3045: douta=16'h7d3a;
3046: douta=16'h8d7b;
3047: douta=16'h7d1b;
3048: douta=16'h7cfa;
3049: douta=16'h7d1a;
3050: douta=16'h853a;
3051: douta=16'h7cfa;
3052: douta=16'h95dd;
3053: douta=16'h53b5;
3054: douta=16'h74da;
3055: douta=16'h8dfd;
3056: douta=16'h74fb;
3057: douta=16'h6cba;
3058: douta=16'h7d5b;
3059: douta=16'h859c;
3060: douta=16'h74fa;
3061: douta=16'h8dbc;
3062: douta=16'h7d5b;
3063: douta=16'h7d1a;
3064: douta=16'h8d9c;
3065: douta=16'h5b72;
3066: douta=16'h326d;
3067: douta=16'h8496;
3068: douta=16'h3aaf;
3069: douta=16'h6c13;
3070: douta=16'h6c14;
3071: douta=16'h5331;
3072: douta=16'h4354;
3073: douta=16'h2a6f;
3074: douta=16'h4333;
3075: douta=16'h6c15;
3076: douta=16'h42f1;
3077: douta=16'h73f4;
3078: douta=16'h5330;
3079: douta=16'h8cb5;
3080: douta=16'h6371;
3081: douta=16'had56;
3082: douta=16'had15;
3083: douta=16'ha4f4;
3084: douta=16'h73af;
3085: douta=16'had13;
3086: douta=16'hbd93;
3087: douta=16'ha4b0;
3088: douta=16'h5269;
3089: douta=16'h8c6f;
3090: douta=16'h942e;
3091: douta=16'h940e;
3092: douta=16'h940d;
3093: douta=16'hc614;
3094: douta=16'h838b;
3095: douta=16'h93cc;
3096: douta=16'h9c0c;
3097: douta=16'hac6c;
3098: douta=16'hb48d;
3099: douta=16'hbcce;
3100: douta=16'hb46d;
3101: douta=16'h9c0c;
3102: douta=16'h9c0d;
3103: douta=16'h732b;
3104: douta=16'h4a29;
3105: douta=16'h2987;
3106: douta=16'h0884;
3107: douta=16'h2126;
3108: douta=16'h18e5;
3109: douta=16'h1105;
3110: douta=16'h0000;
3111: douta=16'h528c;
3112: douta=16'h530e;
3113: douta=16'h2987;
3114: douta=16'h7bef;
3115: douta=16'h6b4c;
3116: douta=16'h426b;
3117: douta=16'h3a8c;
3118: douta=16'h5b2e;
3119: douta=16'h5b0d;
3120: douta=16'h4a8c;
3121: douta=16'h29c9;
3122: douta=16'h2a0b;
3123: douta=16'h5b4f;
3124: douta=16'h5bd3;
3125: douta=16'h5372;
3126: douta=16'h428e;
3127: douta=16'h5b2f;
3128: douta=16'h5b70;
3129: douta=16'h4b0f;
3130: douta=16'h29a8;
3131: douta=16'h3166;
3132: douta=16'h9d39;
3133: douta=16'h8d59;
3134: douta=16'h8539;
3135: douta=16'h7cb8;
3136: douta=16'h7cb8;
3137: douta=16'h957a;
3138: douta=16'h7477;
3139: douta=16'h8d5a;
3140: douta=16'h6415;
3141: douta=16'h7cd8;
3142: douta=16'h7c77;
3143: douta=16'h7cd8;
3144: douta=16'h8518;
3145: douta=16'h8cf8;
3146: douta=16'h8cf8;
3147: douta=16'h9ddc;
3148: douta=16'hb63d;
3149: douta=16'h959b;
3150: douta=16'hb65d;
3151: douta=16'h9dbc;
3152: douta=16'h8d7b;
3153: douta=16'h8d3a;
3154: douta=16'h7cd8;
3155: douta=16'h853a;
3156: douta=16'h84f9;
3157: douta=16'h95bb;
3158: douta=16'h84f9;
3159: douta=16'h853a;
3160: douta=16'h7497;
3161: douta=16'h7477;
3162: douta=16'h8d5a;
3163: douta=16'h6c16;
3164: douta=16'h84f9;
3165: douta=16'h63f5;
3166: douta=16'h7cf9;
3167: douta=16'h8d5b;
3168: douta=16'h7498;
3169: douta=16'h6c57;
3170: douta=16'h7d1a;
3171: douta=16'h74d9;
3172: douta=16'h8d9b;
3173: douta=16'h74b8;
3174: douta=16'h8d7c;
3175: douta=16'h74b9;
3176: douta=16'h959c;
3177: douta=16'h853a;
3178: douta=16'h8d5b;
3179: douta=16'h7d1a;
3180: douta=16'h855a;
3181: douta=16'h855b;
3182: douta=16'h8ddd;
3183: douta=16'h5bd5;
3184: douta=16'h74fa;
3185: douta=16'h6cda;
3186: douta=16'h6cda;
3187: douta=16'h7d5b;
3188: douta=16'h857b;
3189: douta=16'h7d5b;
3190: douta=16'h7d3b;
3191: douta=16'h7d3b;
3192: douta=16'h855b;
3193: douta=16'h7cd9;
3194: douta=16'h10c5;
3195: douta=16'h6bf4;
3196: douta=16'h7434;
3197: douta=16'h9d78;
3198: douta=16'ha5b9;
3199: douta=16'h42d0;
3200: douta=16'h4b95;
3201: douta=16'h4312;
3202: douta=16'h4b74;
3203: douta=16'h7477;
3204: douta=16'h5352;
3205: douta=16'h6bf3;
3206: douta=16'h5b92;
3207: douta=16'h8cb5;
3208: douta=16'h6bd2;
3209: douta=16'hb535;
3210: douta=16'h7c12;
3211: douta=16'h7b90;
3212: douta=16'h4a6c;
3213: douta=16'ha4f2;
3214: douta=16'hb552;
3215: douta=16'h944f;
3216: douta=16'h7bac;
3217: douta=16'hbd92;
3218: douta=16'h7b4c;
3219: douta=16'hb531;
3220: douta=16'haccf;
3221: douta=16'h7309;
3222: douta=16'h9c0d;
3223: douta=16'h9c0d;
3224: douta=16'hac4c;
3225: douta=16'hb4cd;
3226: douta=16'hcd4e;
3227: douta=16'hd570;
3228: douta=16'hcd6f;
3229: douta=16'hac4d;
3230: douta=16'h8b8c;
3231: douta=16'h5a68;
3232: douta=16'h5a6a;
3233: douta=16'h2967;
3234: douta=16'h528a;
3235: douta=16'h08a4;
3236: douta=16'h10e5;
3237: douta=16'h10e4;
3238: douta=16'h1926;
3239: douta=16'h0000;
3240: douta=16'h6391;
3241: douta=16'h428b;
3242: douta=16'h52cb;
3243: douta=16'h6b4d;
3244: douta=16'h3a2a;
3245: douta=16'h29ea;
3246: douta=16'h29a8;
3247: douta=16'h73ae;
3248: douta=16'h4aee;
3249: douta=16'h42ce;
3250: douta=16'h08a5;
3251: douta=16'h29c9;
3252: douta=16'h2189;
3253: douta=16'h32ae;
3254: douta=16'h3a6d;
3255: douta=16'h3a4c;
3256: douta=16'h3aaf;
3257: douta=16'h5371;
3258: douta=16'h4aaf;
3259: douta=16'hb48d;
3260: douta=16'h84f9;
3261: douta=16'h84d8;
3262: douta=16'h955a;
3263: douta=16'h7477;
3264: douta=16'h84d8;
3265: douta=16'h7477;
3266: douta=16'h955a;
3267: douta=16'h8cf8;
3268: douta=16'h84d8;
3269: douta=16'h8d3a;
3270: douta=16'h6415;
3271: douta=16'h7cb7;
3272: douta=16'h8d39;
3273: douta=16'h84f8;
3274: douta=16'hae1b;
3275: douta=16'h957b;
3276: douta=16'h9dfb;
3277: douta=16'h7d19;
3278: douta=16'h84f9;
3279: douta=16'h95db;
3280: douta=16'h9ddb;
3281: douta=16'h7cd9;
3282: douta=16'h8d7a;
3283: douta=16'h8d7a;
3284: douta=16'h8519;
3285: douta=16'h8d39;
3286: douta=16'h957b;
3287: douta=16'h8d5a;
3288: douta=16'h74b8;
3289: douta=16'h853a;
3290: douta=16'h7cd9;
3291: douta=16'h7477;
3292: douta=16'h7498;
3293: douta=16'h8d3a;
3294: douta=16'h851a;
3295: douta=16'h851a;
3296: douta=16'h7498;
3297: douta=16'h74b8;
3298: douta=16'h7cfa;
3299: douta=16'h6c77;
3300: douta=16'h6c77;
3301: douta=16'h6436;
3302: douta=16'h95dc;
3303: douta=16'h855b;
3304: douta=16'h7cf9;
3305: douta=16'h7d1a;
3306: douta=16'h8d5b;
3307: douta=16'h95dc;
3308: douta=16'h855c;
3309: douta=16'h7cfa;
3310: douta=16'h853b;
3311: douta=16'h857c;
3312: douta=16'h74f9;
3313: douta=16'h8d9c;
3314: douta=16'h6479;
3315: douta=16'h7d3b;
3316: douta=16'h6cb9;
3317: douta=16'h7d5a;
3318: douta=16'h95dc;
3319: douta=16'h7cf9;
3320: douta=16'h7d5b;
3321: douta=16'h7d3a;
3322: douta=16'h2167;
3323: douta=16'hb5d9;
3324: douta=16'h5b72;
3325: douta=16'h8474;
3326: douta=16'h9cf5;
3327: douta=16'h73b0;
3328: douta=16'h4394;
3329: douta=16'h2a8f;
3330: douta=16'h5c36;
3331: douta=16'h7497;
3332: douta=16'h5b93;
3333: douta=16'h7414;
3334: douta=16'h8cd7;
3335: douta=16'h9537;
3336: douta=16'h9d36;
3337: douta=16'h9492;
3338: douta=16'h9cf3;
3339: douta=16'ha4d2;
3340: douta=16'h4aad;
3341: douta=16'h9c90;
3342: douta=16'hbd72;
3343: douta=16'hc5b3;
3344: douta=16'hbd72;
3345: douta=16'hb552;
3346: douta=16'h83cd;
3347: douta=16'hcdf3;
3348: douta=16'h7b0a;
3349: douta=16'h838b;
3350: douta=16'h93cc;
3351: douta=16'hac6c;
3352: douta=16'hbd0e;
3353: douta=16'hcd6f;
3354: douta=16'hddd2;
3355: douta=16'hddd1;
3356: douta=16'hd5b1;
3357: douta=16'hddf3;
3358: douta=16'hc50e;
3359: douta=16'h940d;
3360: douta=16'h4a2a;
3361: douta=16'h52ab;
3362: douta=16'h62cb;
3363: douta=16'h2967;
3364: douta=16'h10e5;
3365: douta=16'h1905;
3366: douta=16'h1904;
3367: douta=16'h0000;
3368: douta=16'h0000;
3369: douta=16'h6370;
3370: douta=16'h2987;
3371: douta=16'h6b0b;
3372: douta=16'h18e4;
3373: douta=16'h10e5;
3374: douta=16'h1106;
3375: douta=16'h4a8d;
3376: douta=16'h2a0c;
3377: douta=16'h118a;
3378: douta=16'h2188;
3379: douta=16'h4a8a;
3380: douta=16'h6baf;
3381: douta=16'h1947;
3382: douta=16'h29a9;
3383: douta=16'h320b;
3384: douta=16'h0927;
3385: douta=16'h2a0c;
3386: douta=16'h326d;
3387: douta=16'h5acb;
3388: douta=16'h84d8;
3389: douta=16'h7cd8;
3390: douta=16'h8d39;
3391: douta=16'h74b8;
3392: douta=16'h957a;
3393: douta=16'h7477;
3394: douta=16'h6c36;
3395: douta=16'h8518;
3396: douta=16'h84d9;
3397: douta=16'h7cb8;
3398: douta=16'ha5db;
3399: douta=16'h6416;
3400: douta=16'h8d39;
3401: douta=16'ha5fc;
3402: douta=16'ha5fb;
3403: douta=16'h8d3a;
3404: douta=16'h9dbc;
3405: douta=16'h851a;
3406: douta=16'ha61d;
3407: douta=16'h7cf9;
3408: douta=16'h6c97;
3409: douta=16'ha5fb;
3410: douta=16'h851a;
3411: douta=16'h8519;
3412: douta=16'h7cd9;
3413: douta=16'h9ddc;
3414: douta=16'h7cd9;
3415: douta=16'h8519;
3416: douta=16'h7cf9;
3417: douta=16'h855a;
3418: douta=16'h7498;
3419: douta=16'h851a;
3420: douta=16'h6c57;
3421: douta=16'h6c77;
3422: douta=16'h7478;
3423: douta=16'h6456;
3424: douta=16'h6416;
3425: douta=16'h6c77;
3426: douta=16'h6c36;
3427: douta=16'h6416;
3428: douta=16'h7477;
3429: douta=16'h7498;
3430: douta=16'h6c36;
3431: douta=16'h6c77;
3432: douta=16'h6c98;
3433: douta=16'h8d9c;
3434: douta=16'h7d3b;
3435: douta=16'h853b;
3436: douta=16'h7d1b;
3437: douta=16'h8dbc;
3438: douta=16'h853b;
3439: douta=16'h8d7c;
3440: douta=16'h7d3a;
3441: douta=16'h7d3a;
3442: douta=16'h74b9;
3443: douta=16'h857b;
3444: douta=16'h74da;
3445: douta=16'h6458;
3446: douta=16'h857b;
3447: douta=16'h857b;
3448: douta=16'h8d9c;
3449: douta=16'h74fa;
3450: douta=16'h6c77;
3451: douta=16'h7c75;
3452: douta=16'h7433;
3453: douta=16'h7413;
3454: douta=16'h94b4;
3455: douta=16'h3a4c;
3456: douta=16'h3b32;
3457: douta=16'h2a2e;
3458: douta=16'h6417;
3459: douta=16'h84b8;
3460: douta=16'h6c76;
3461: douta=16'h7c75;
3462: douta=16'h8cd7;
3463: douta=16'h9d16;
3464: douta=16'h8475;
3465: douta=16'h7bf1;
3466: douta=16'hc5b5;
3467: douta=16'hc5f5;
3468: douta=16'h632c;
3469: douta=16'h8bee;
3470: douta=16'ha4d1;
3471: douta=16'heef8;
3472: douta=16'h732b;
3473: douta=16'hb531;
3474: douta=16'h946d;
3475: douta=16'h6ae9;
3476: douta=16'h72ea;
3477: douta=16'h93eb;
3478: douta=16'h93cb;
3479: douta=16'hb48d;
3480: douta=16'hcd6f;
3481: douta=16'hddf3;
3482: douta=16'hde13;
3483: douta=16'he634;
3484: douta=16'hddf3;
3485: douta=16'hcd6f;
3486: douta=16'he653;
3487: douta=16'h3165;
3488: douta=16'hacd0;
3489: douta=16'h39e9;
3490: douta=16'h6aeb;
3491: douta=16'h29a8;
3492: douta=16'h2126;
3493: douta=16'h10a3;
3494: douta=16'h18e4;
3495: douta=16'h2145;
3496: douta=16'h0001;
3497: douta=16'h1106;
3498: douta=16'h1905;
3499: douta=16'h10e5;
3500: douta=16'h0842;
3501: douta=16'h4208;
3502: douta=16'h4208;
3503: douta=16'h630d;
3504: douta=16'h4aac;
3505: douta=16'h1948;
3506: douta=16'h31c9;
3507: douta=16'h4aab;
3508: douta=16'h8410;
3509: douta=16'h3a09;
3510: douta=16'h1947;
3511: douta=16'h29ca;
3512: douta=16'h3187;
3513: douta=16'h530f;
3514: douta=16'h6ace;
3515: douta=16'ha598;
3516: douta=16'h6436;
3517: douta=16'h9dbb;
3518: douta=16'h8519;
3519: douta=16'h8519;
3520: douta=16'h9d9a;
3521: douta=16'h7cd8;
3522: douta=16'h6c56;
3523: douta=16'ha5dc;
3524: douta=16'h5bf5;
3525: douta=16'h9dbb;
3526: douta=16'h8519;
3527: douta=16'h9559;
3528: douta=16'h8d39;
3529: douta=16'h8d3a;
3530: douta=16'h7cd8;
3531: douta=16'h853a;
3532: douta=16'h957a;
3533: douta=16'h959a;
3534: douta=16'h84f9;
3535: douta=16'h7cd9;
3536: douta=16'hae1c;
3537: douta=16'h6417;
3538: douta=16'h851a;
3539: douta=16'h959b;
3540: douta=16'h84f9;
3541: douta=16'h955a;
3542: douta=16'h53b4;
3543: douta=16'h853a;
3544: douta=16'h6cb8;
3545: douta=16'h7d3b;
3546: douta=16'h7cd9;
3547: douta=16'h7d1a;
3548: douta=16'h6c36;
3549: douta=16'h6c57;
3550: douta=16'h7477;
3551: douta=16'h6c77;
3552: douta=16'h7cf9;
3553: douta=16'h6436;
3554: douta=16'h7498;
3555: douta=16'h6c15;
3556: douta=16'h853a;
3557: douta=16'h6415;
3558: douta=16'h5bd4;
3559: douta=16'h6c78;
3560: douta=16'h855a;
3561: douta=16'h6c78;
3562: douta=16'h8d9c;
3563: douta=16'h855c;
3564: douta=16'h74fa;
3565: douta=16'h859c;
3566: douta=16'h7d3a;
3567: douta=16'h7cfa;
3568: douta=16'h855c;
3569: douta=16'h857b;
3570: douta=16'h74d9;
3571: douta=16'h7d1a;
3572: douta=16'h6c99;
3573: douta=16'h857c;
3574: douta=16'h53f6;
3575: douta=16'h7d3a;
3576: douta=16'h857b;
3577: douta=16'h8dbc;
3578: douta=16'h7d1b;
3579: douta=16'h52cd;
3580: douta=16'h8453;
3581: douta=16'h63b2;
3582: douta=16'h42cf;
3583: douta=16'h73d2;
3584: douta=16'h3312;
3585: douta=16'h2a50;
3586: douta=16'h5bf6;
3587: douta=16'h7c97;
3588: douta=16'h7c97;
3589: douta=16'h4acf;
3590: douta=16'h5b92;
3591: douta=16'h8454;
3592: douta=16'h8c94;
3593: douta=16'h8c71;
3594: douta=16'h7bd0;
3595: douta=16'hbd74;
3596: douta=16'h7b8e;
3597: douta=16'hd635;
3598: douta=16'h7bce;
3599: douta=16'hbd52;
3600: douta=16'h738c;
3601: douta=16'h8c2d;
3602: douta=16'h9c90;
3603: douta=16'h730a;
3604: douta=16'h8bab;
3605: douta=16'ha40c;
3606: douta=16'hac6c;
3607: douta=16'hc50e;
3608: douta=16'hddd2;
3609: douta=16'hde33;
3610: douta=16'he654;
3611: douta=16'hddd2;
3612: douta=16'hddf3;
3613: douta=16'hbcce;
3614: douta=16'hac4d;
3615: douta=16'ha46e;
3616: douta=16'ha46e;
3617: douta=16'h39ea;
3618: douta=16'h734c;
3619: douta=16'h39c9;
3620: douta=16'h2188;
3621: douta=16'h2967;
3622: douta=16'h0883;
3623: douta=16'h10e4;
3624: douta=16'h1905;
3625: douta=16'h0042;
3626: douta=16'h2168;
3627: douta=16'h18e5;
3628: douta=16'h18e6;
3629: douta=16'h18e4;
3630: douta=16'h944e;
3631: douta=16'h9c8f;
3632: douta=16'h5b0c;
3633: douta=16'h320b;
3634: douta=16'h530d;
3635: douta=16'h29ea;
3636: douta=16'h3a4c;
3637: douta=16'h322a;
3638: douta=16'h1127;
3639: douta=16'h1969;
3640: douta=16'h5b0c;
3641: douta=16'h39c8;
3642: douta=16'hac6f;
3643: douta=16'h8d7a;
3644: douta=16'h6c56;
3645: douta=16'h5b93;
3646: douta=16'h5353;
3647: douta=16'h8d19;
3648: douta=16'h74b7;
3649: douta=16'h9d7b;
3650: douta=16'h7497;
3651: douta=16'h9ddc;
3652: douta=16'h7cd9;
3653: douta=16'h955a;
3654: douta=16'h7478;
3655: douta=16'h84f9;
3656: douta=16'h8d5a;
3657: douta=16'ha5db;
3658: douta=16'h9559;
3659: douta=16'ha5fb;
3660: douta=16'h6c77;
3661: douta=16'h8d7a;
3662: douta=16'h959a;
3663: douta=16'hae5d;
3664: douta=16'h7cb7;
3665: douta=16'h5bf5;
3666: douta=16'h851a;
3667: douta=16'h7477;
3668: douta=16'h4b74;
3669: douta=16'h7cd9;
3670: douta=16'h857c;
3671: douta=16'h6498;
3672: douta=16'h6437;
3673: douta=16'h53d5;
3674: douta=16'h7d1a;
3675: douta=16'h7d1a;
3676: douta=16'h7497;
3677: douta=16'h6c36;
3678: douta=16'h7c97;
3679: douta=16'h63d4;
3680: douta=16'h63f4;
3681: douta=16'h7c96;
3682: douta=16'h7496;
3683: douta=16'h7456;
3684: douta=16'h7c97;
3685: douta=16'h63f4;
3686: douta=16'h7457;
3687: douta=16'h74d9;
3688: douta=16'h5c16;
3689: douta=16'h6478;
3690: douta=16'h6498;
3691: douta=16'h74fa;
3692: douta=16'h859c;
3693: douta=16'h6cba;
3694: douta=16'h855b;
3695: douta=16'h74da;
3696: douta=16'h855b;
3697: douta=16'h7d1a;
3698: douta=16'h8d7c;
3699: douta=16'h853a;
3700: douta=16'h7d1a;
3701: douta=16'h8d7b;
3702: douta=16'h7d3a;
3703: douta=16'h855b;
3704: douta=16'h74b8;
3705: douta=16'h8d9c;
3706: douta=16'h751a;
3707: douta=16'h2126;
3708: douta=16'h6370;
3709: douta=16'h8c94;
3710: douta=16'h532f;
3711: douta=16'h6390;
3712: douta=16'h4374;
3713: douta=16'h2a90;
3714: douta=16'h4353;
3715: douta=16'h5352;
3716: douta=16'h84f8;
3717: douta=16'h3a4e;
3718: douta=16'h6bf4;
3719: douta=16'h7c33;
3720: douta=16'h8c93;
3721: douta=16'h94d3;
3722: douta=16'h7c31;
3723: douta=16'hbd74;
3724: douta=16'had12;
3725: douta=16'ha4b1;
3726: douta=16'h736d;
3727: douta=16'ha4d1;
3728: douta=16'h7bad;
3729: douta=16'h8c0e;
3730: douta=16'h8b8c;
3731: douta=16'h836a;
3732: douta=16'h93aa;
3733: douta=16'hb4ad;
3734: douta=16'hbcac;
3735: douta=16'hcd90;
3736: douta=16'he654;
3737: douta=16'he654;
3738: douta=16'he654;
3739: douta=16'hd5b1;
3740: douta=16'hc52f;
3741: douta=16'hb48e;
3742: douta=16'hc52f;
3743: douta=16'hbd30;
3744: douta=16'hacaf;
3745: douta=16'h6aec;
3746: douta=16'h83ae;
3747: douta=16'h422a;
3748: douta=16'h29a8;
3749: douta=16'h1926;
3750: douta=16'h2147;
3751: douta=16'h1905;
3752: douta=16'h10a3;
3753: douta=16'h10c4;
3754: douta=16'h0000;
3755: douta=16'h1106;
3756: douta=16'h10a5;
3757: douta=16'h29a7;
3758: douta=16'h8bed;
3759: douta=16'h734c;
3760: douta=16'h2966;
3761: douta=16'h5aec;
3762: douta=16'h3a4b;
3763: douta=16'h1147;
3764: douta=16'h31ca;
3765: douta=16'h426c;
3766: douta=16'h1129;
3767: douta=16'h0044;
3768: douta=16'h52ed;
3769: douta=16'h2167;
3770: douta=16'h836a;
3771: douta=16'h8d39;
3772: douta=16'h9dba;
3773: douta=16'h9d9a;
3774: douta=16'h8d59;
3775: douta=16'hadfc;
3776: douta=16'h5b93;
3777: douta=16'h6435;
3778: douta=16'h8d7a;
3779: douta=16'h957a;
3780: douta=16'h8d3a;
3781: douta=16'h957b;
3782: douta=16'h853a;
3783: douta=16'h8d5a;
3784: douta=16'h8d1a;
3785: douta=16'h959b;
3786: douta=16'h8d3a;
3787: douta=16'h7cd9;
3788: douta=16'h9dbb;
3789: douta=16'h6c77;
3790: douta=16'h957a;
3791: douta=16'hbe9e;
3792: douta=16'h5331;
3793: douta=16'h6c56;
3794: douta=16'h6c56;
3795: douta=16'h6436;
3796: douta=16'h5373;
3797: douta=16'h6416;
3798: douta=16'h328f;
3799: douta=16'h6cb9;
3800: douta=16'h5bd6;
3801: douta=16'h6457;
3802: douta=16'h6416;
3803: douta=16'h4b53;
3804: douta=16'h7cd8;
3805: douta=16'h7497;
3806: douta=16'h7436;
3807: douta=16'h7c77;
3808: douta=16'h7c97;
3809: douta=16'h7c96;
3810: douta=16'h7457;
3811: douta=16'h6c35;
3812: douta=16'h7455;
3813: douta=16'h5373;
3814: douta=16'h4311;
3815: douta=16'h3b13;
3816: douta=16'h6cb9;
3817: douta=16'h5c58;
3818: douta=16'h6c99;
3819: douta=16'h6458;
3820: douta=16'h74da;
3821: douta=16'h74da;
3822: douta=16'h857c;
3823: douta=16'h74d9;
3824: douta=16'h7d3a;
3825: douta=16'h7d3a;
3826: douta=16'h74fa;
3827: douta=16'h7d3b;
3828: douta=16'h8d9c;
3829: douta=16'h7499;
3830: douta=16'h8d9c;
3831: douta=16'h7cd9;
3832: douta=16'h8d7b;
3833: douta=16'h7d1a;
3834: douta=16'h6417;
3835: douta=16'h1906;
3836: douta=16'h7c13;
3837: douta=16'h63d3;
3838: douta=16'h42cf;
3839: douta=16'h6bb1;
3840: douta=16'h4353;
3841: douta=16'h4bd6;
3842: douta=16'h32d2;
3843: douta=16'h326e;
3844: douta=16'h7456;
3845: douta=16'h5330;
3846: douta=16'h7414;
3847: douta=16'h7c32;
3848: douta=16'ha516;
3849: douta=16'h8c93;
3850: douta=16'h6bb0;
3851: douta=16'h8c51;
3852: douta=16'hce36;
3853: douta=16'hd678;
3854: douta=16'ha4b2;
3855: douta=16'had12;
3856: douta=16'hc5d4;
3857: douta=16'h6aa9;
3858: douta=16'h9beb;
3859: douta=16'h93ec;
3860: douta=16'hb48c;
3861: douta=16'hb4ad;
3862: douta=16'hcd2f;
3863: douta=16'he634;
3864: douta=16'he633;
3865: douta=16'hddd2;
3866: douta=16'hc50f;
3867: douta=16'hd590;
3868: douta=16'hb48e;
3869: douta=16'h9beb;
3870: douta=16'hb48e;
3871: douta=16'hcd71;
3872: douta=16'hb4cf;
3873: douta=16'h940e;
3874: douta=16'h8bef;
3875: douta=16'h4a8b;
3876: douta=16'h4a4a;
3877: douta=16'h29ca;
3878: douta=16'h2168;
3879: douta=16'h422a;
3880: douta=16'h18e5;
3881: douta=16'h10e4;
3882: douta=16'h10a4;
3883: douta=16'h10e5;
3884: douta=16'h0000;
3885: douta=16'h4ace;
3886: douta=16'h4a28;
3887: douta=16'h39e8;
3888: douta=16'h732c;
3889: douta=16'h1063;
3890: douta=16'h1105;
3891: douta=16'h52aa;
3892: douta=16'h9470;
3893: douta=16'h6b4d;
3894: douta=16'h1128;
3895: douta=16'h320b;
3896: douta=16'h52cc;
3897: douta=16'h2169;
3898: douta=16'h62ca;
3899: douta=16'h9d9a;
3900: douta=16'h8d18;
3901: douta=16'h9d9a;
3902: douta=16'h957a;
3903: douta=16'h9559;
3904: douta=16'h9d9a;
3905: douta=16'h9d9a;
3906: douta=16'ha5fb;
3907: douta=16'h5bf6;
3908: douta=16'h8519;
3909: douta=16'h7cd9;
3910: douta=16'h957b;
3911: douta=16'ha5dc;
3912: douta=16'h957b;
3913: douta=16'h9dbc;
3914: douta=16'h6457;
3915: douta=16'h8d3a;
3916: douta=16'h7497;
3917: douta=16'hb65d;
3918: douta=16'h7477;
3919: douta=16'h8d59;
3920: douta=16'h940f;
3921: douta=16'h10e5;
3922: douta=16'h1948;
3923: douta=16'h4bf6;
3924: douta=16'h4374;
3925: douta=16'h5bf5;
3926: douta=16'h5bd4;
3927: douta=16'h5bb3;
3928: douta=16'h328e;
3929: douta=16'h7436;
3930: douta=16'h6c97;
3931: douta=16'h6c98;
3932: douta=16'h5c16;
3933: douta=16'h6436;
3934: douta=16'h5bb4;
3935: douta=16'h955a;
3936: douta=16'h7435;
3937: douta=16'h6c14;
3938: douta=16'h7c75;
3939: douta=16'h4a6a;
3940: douta=16'h2125;
3941: douta=16'h1a4f;
3942: douta=16'h3b75;
3943: douta=16'h4395;
3944: douta=16'h5c58;
3945: douta=16'h4395;
3946: douta=16'h6cba;
3947: douta=16'h7d3b;
3948: douta=16'h6c99;
3949: douta=16'h74fa;
3950: douta=16'h5bf7;
3951: douta=16'h7d1a;
3952: douta=16'h7d3a;
3953: douta=16'h7cfa;
3954: douta=16'h857c;
3955: douta=16'h7d1a;
3956: douta=16'h855c;
3957: douta=16'h7499;
3958: douta=16'h8d7b;
3959: douta=16'h855b;
3960: douta=16'h8d7b;
3961: douta=16'h6478;
3962: douta=16'h857b;
3963: douta=16'h1906;
3964: douta=16'h84b6;
3965: douta=16'h6bb1;
3966: douta=16'h1149;
3967: douta=16'h7c74;
3968: douta=16'h19cc;
3969: douta=16'h3333;
3970: douta=16'h2a90;
3971: douta=16'h53d4;
3972: douta=16'h6c15;
3973: douta=16'h5331;
3974: douta=16'h8cf8;
3975: douta=16'h8c54;
3976: douta=16'h9cd6;
3977: douta=16'had56;
3978: douta=16'ha514;
3979: douta=16'h8c50;
3980: douta=16'hc5f6;
3981: douta=16'hd657;
3982: douta=16'h8c50;
3983: douta=16'h8c71;
3984: douta=16'h8bac;
3985: douta=16'h8bab;
3986: douta=16'hb48d;
3987: douta=16'hac6b;
3988: douta=16'hac8d;
3989: douta=16'hd56f;
3990: douta=16'hde33;
3991: douta=16'he675;
3992: douta=16'hde33;
3993: douta=16'hddf3;
3994: douta=16'h9c0d;
3995: douta=16'hbcae;
3996: douta=16'h8b8a;
3997: douta=16'hb4ae;
3998: douta=16'hc54f;
3999: douta=16'hd5d2;
4000: douta=16'hc550;
4001: douta=16'hb4d0;
4002: douta=16'ha470;
4003: douta=16'h736e;
4004: douta=16'h630e;
4005: douta=16'h428c;
4006: douta=16'h31eb;
4007: douta=16'h1906;
4008: douta=16'h526b;
4009: douta=16'h18a4;
4010: douta=16'h10a4;
4011: douta=16'h08a4;
4012: douta=16'h18e5;
4013: douta=16'h2988;
4014: douta=16'h4acd;
4015: douta=16'h0001;
4016: douta=16'h0842;
4017: douta=16'h62aa;
4018: douta=16'h5289;
4019: douta=16'h6b4c;
4020: douta=16'h52ec;
4021: douta=16'hb532;
4022: douta=16'h6b2d;
4023: douta=16'h636f;
4024: douta=16'h8430;
4025: douta=16'h7bef;
4026: douta=16'h732b;
4027: douta=16'h84b7;
4028: douta=16'h8d39;
4029: douta=16'h9579;
4030: douta=16'h9579;
4031: douta=16'h8d39;
4032: douta=16'h8d38;
4033: douta=16'ha5ba;
4034: douta=16'h957a;
4035: douta=16'h9d9a;
4036: douta=16'h9dba;
4037: douta=16'h8d39;
4038: douta=16'h5bf6;
4039: douta=16'h9dbb;
4040: douta=16'h955b;
4041: douta=16'h95bb;
4042: douta=16'h959b;
4043: douta=16'h6c58;
4044: douta=16'h7cf9;
4045: douta=16'ha5fc;
4046: douta=16'h6c56;
4047: douta=16'h8518;
4048: douta=16'h94d6;
4049: douta=16'h1925;
4050: douta=16'h0883;
4051: douta=16'h4b32;
4052: douta=16'h7cd8;
4053: douta=16'h7497;
4054: douta=16'h7498;
4055: douta=16'h7cb7;
4056: douta=16'h7456;
4057: douta=16'h6415;
4058: douta=16'h5393;
4059: douta=16'h5b73;
4060: douta=16'h6c77;
4061: douta=16'h6c77;
4062: douta=16'h5373;
4063: douta=16'h5bb3;
4064: douta=16'h5372;
4065: douta=16'h9d9a;
4066: douta=16'h7c34;
4067: douta=16'h2967;
4068: douta=16'h10e5;
4069: douta=16'h7cd9;
4070: douta=16'h6c57;
4071: douta=16'h6cb9;
4072: douta=16'h53b6;
4073: douta=16'h6479;
4074: douta=16'h74fa;
4075: douta=16'h5c37;
4076: douta=16'h53f6;
4077: douta=16'h74f9;
4078: douta=16'h7d1a;
4079: douta=16'h7d3a;
4080: douta=16'h7478;
4081: douta=16'h6416;
4082: douta=16'h855b;
4083: douta=16'h8d9c;
4084: douta=16'h7d3a;
4085: douta=16'h7d1a;
4086: douta=16'h8dbc;
4087: douta=16'h7cd9;
4088: douta=16'h855b;
4089: douta=16'h853a;
4090: douta=16'h7d3a;
4091: douta=16'h39ea;
4092: douta=16'h9d57;
4093: douta=16'h7413;
4094: douta=16'h73f3;
4095: douta=16'h9517;
4096: douta=16'h2a90;
4097: douta=16'h3313;
4098: douta=16'h2a90;
4099: douta=16'h6457;
4100: douta=16'h8519;
4101: douta=16'h5b93;
4102: douta=16'h6392;
4103: douta=16'h7c54;
4104: douta=16'h94b5;
4105: douta=16'hb5b6;
4106: douta=16'ha4f3;
4107: douta=16'hb533;
4108: douta=16'had54;
4109: douta=16'hd677;
4110: douta=16'h9491;
4111: douta=16'h72c8;
4112: douta=16'h8b8b;
4113: douta=16'ha42b;
4114: douta=16'h8b69;
4115: douta=16'hbccd;
4116: douta=16'hcd2e;
4117: douta=16'he634;
4118: douta=16'hee96;
4119: douta=16'heeb6;
4120: douta=16'hddf4;
4121: douta=16'hbd0f;
4122: douta=16'hac4d;
4123: douta=16'h7b07;
4124: douta=16'hc52f;
4125: douta=16'ha42c;
4126: douta=16'hd5b2;
4127: douta=16'hd5b2;
4128: douta=16'hcd71;
4129: douta=16'hc530;
4130: douta=16'h9c70;
4131: douta=16'h83ef;
4132: douta=16'h6b6f;
4133: douta=16'h5b2e;
4134: douta=16'h428d;
4135: douta=16'h29aa;
4136: douta=16'h08e6;
4137: douta=16'h08a4;
4138: douta=16'h10a4;
4139: douta=16'h10c4;
4140: douta=16'h10e4;
4141: douta=16'h2125;
4142: douta=16'h2a2c;
4143: douta=16'h5b0e;
4144: douta=16'h8c50;
4145: douta=16'had11;
4146: douta=16'h5aaa;
4147: douta=16'h0000;
4148: douta=16'h0042;
4149: douta=16'h83ee;
4150: douta=16'h73ef;
4151: douta=16'h39ea;
4152: douta=16'h29a8;
4153: douta=16'h5b0d;
4154: douta=16'h7b6c;
4155: douta=16'h8517;
4156: douta=16'h8d18;
4157: douta=16'h84f8;
4158: douta=16'h8d18;
4159: douta=16'h8d38;
4160: douta=16'h9559;
4161: douta=16'h8d59;
4162: douta=16'h9dba;
4163: douta=16'h9559;
4164: douta=16'h9559;
4165: douta=16'h957a;
4166: douta=16'ha5ba;
4167: douta=16'h9dda;
4168: douta=16'h9d9a;
4169: douta=16'h7498;
4170: douta=16'h8d5a;
4171: douta=16'h95bb;
4172: douta=16'ha5fc;
4173: douta=16'h8d3a;
4174: douta=16'h7c77;
4175: douta=16'h7cb7;
4176: douta=16'h84f9;
4177: douta=16'h4a09;
4178: douta=16'h10c4;
4179: douta=16'h9539;
4180: douta=16'h7c97;
4181: douta=16'h84d8;
4182: douta=16'h9d9b;
4183: douta=16'h84d8;
4184: douta=16'h63f4;
4185: douta=16'h959b;
4186: douta=16'h853a;
4187: douta=16'h8d19;
4188: douta=16'h63b4;
4189: douta=16'h63d4;
4190: douta=16'h84f8;
4191: douta=16'h7456;
4192: douta=16'h7cd8;
4193: douta=16'h6bf5;
4194: douta=16'h6c35;
4195: douta=16'h2125;
4196: douta=16'h10e4;
4197: douta=16'h6456;
4198: douta=16'h6436;
4199: douta=16'h74d9;
4200: douta=16'h74d9;
4201: douta=16'h6cda;
4202: douta=16'h6c78;
4203: douta=16'h6457;
4204: douta=16'h6c98;
4205: douta=16'h7498;
4206: douta=16'h6c36;
4207: douta=16'h7cd9;
4208: douta=16'h74b8;
4209: douta=16'h7cd9;
4210: douta=16'h855b;
4211: douta=16'h7cb8;
4212: douta=16'h74d9;
4213: douta=16'h7cf9;
4214: douta=16'h855b;
4215: douta=16'h74d9;
4216: douta=16'h8d7b;
4217: douta=16'h7cb9;
4218: douta=16'h7d3a;
4219: douta=16'h7c53;
4220: douta=16'h84b6;
4221: douta=16'h6391;
4222: douta=16'h6391;
4223: douta=16'h20e3;
4224: douta=16'h4375;
4225: douta=16'h4b54;
4226: douta=16'h32d1;
4227: douta=16'h6458;
4228: douta=16'h84f9;
4229: douta=16'h63d4;
4230: douta=16'h73f3;
4231: douta=16'h5b92;
4232: douta=16'h9cf5;
4233: douta=16'hb576;
4234: douta=16'had35;
4235: douta=16'hb534;
4236: douta=16'hbdb5;
4237: douta=16'hce36;
4238: douta=16'h7b09;
4239: douta=16'h93cb;
4240: douta=16'hac4c;
4241: douta=16'hbc8b;
4242: douta=16'hb48c;
4243: douta=16'hd5b0;
4244: douta=16'hde12;
4245: douta=16'hee75;
4246: douta=16'he634;
4247: douta=16'he674;
4248: douta=16'hc550;
4249: douta=16'hc551;
4250: douta=16'h72e8;
4251: douta=16'h93ec;
4252: douta=16'h9c0d;
4253: douta=16'hde13;
4254: douta=16'hd5f3;
4255: douta=16'hddf3;
4256: douta=16'hd591;
4257: douta=16'hcd50;
4258: douta=16'hacb0;
4259: douta=16'h8c10;
4260: douta=16'h6b6f;
4261: douta=16'h6b70;
4262: douta=16'h5b50;
4263: douta=16'h42af;
4264: douta=16'h324d;
4265: douta=16'h2988;
4266: douta=16'h0063;
4267: douta=16'h10e4;
4268: douta=16'h10e4;
4269: douta=16'h10a4;
4270: douta=16'h2967;
4271: douta=16'h3acf;
4272: douta=16'h1926;
4273: douta=16'h2167;
4274: douta=16'h6b0a;
4275: douta=16'h39a6;
4276: douta=16'h3145;
4277: douta=16'h4228;
4278: douta=16'h528a;
4279: douta=16'h942f;
4280: douta=16'h0064;
4281: douta=16'h1105;
4282: douta=16'h72eb;
4283: douta=16'h5bb4;
4284: douta=16'h8d37;
4285: douta=16'h9579;
4286: douta=16'h9539;
4287: douta=16'h8d18;
4288: douta=16'h84f8;
4289: douta=16'h8d18;
4290: douta=16'h8d18;
4291: douta=16'h957a;
4292: douta=16'h9559;
4293: douta=16'h9d9a;
4294: douta=16'h8d39;
4295: douta=16'h9559;
4296: douta=16'ha5db;
4297: douta=16'ha5db;
4298: douta=16'h959a;
4299: douta=16'h9d9a;
4300: douta=16'h7497;
4301: douta=16'h9ddc;
4302: douta=16'h8d39;
4303: douta=16'h84f8;
4304: douta=16'h6c14;
4305: douta=16'h838b;
4306: douta=16'h1905;
4307: douta=16'h8cf8;
4308: douta=16'h8d18;
4309: douta=16'h9d7a;
4310: douta=16'h9dba;
4311: douta=16'h8d39;
4312: douta=16'h7cb7;
4313: douta=16'h8d39;
4314: douta=16'h84f8;
4315: douta=16'h8539;
4316: douta=16'h8d7a;
4317: douta=16'h957a;
4318: douta=16'h9559;
4319: douta=16'h63d3;
4320: douta=16'h9539;
4321: douta=16'h8518;
4322: douta=16'h6c15;
4323: douta=16'h2146;
4324: douta=16'h1905;
4325: douta=16'h5c16;
4326: douta=16'h751a;
4327: douta=16'h6cb9;
4328: douta=16'h6cb8;
4329: douta=16'h74da;
4330: douta=16'h6cb9;
4331: douta=16'h74d9;
4332: douta=16'h7cf9;
4333: douta=16'h74b9;
4334: douta=16'h7457;
4335: douta=16'h7d1a;
4336: douta=16'h5bd5;
4337: douta=16'h8d5b;
4338: douta=16'h7498;
4339: douta=16'h851a;
4340: douta=16'h853a;
4341: douta=16'h853b;
4342: douta=16'h855a;
4343: douta=16'h8519;
4344: douta=16'h853a;
4345: douta=16'h851a;
4346: douta=16'h6c77;
4347: douta=16'hdefd;
4348: douta=16'h8496;
4349: douta=16'ha558;
4350: douta=16'h8cd4;
4351: douta=16'h3a2a;
4352: douta=16'h2a6f;
4353: douta=16'h3b33;
4354: douta=16'h2ab0;
4355: douta=16'h4b75;
4356: douta=16'h63d4;
4357: douta=16'h7477;
4358: douta=16'h6bf3;
4359: douta=16'h5b72;
4360: douta=16'h8c74;
4361: douta=16'hb5b7;
4362: douta=16'ha515;
4363: douta=16'h9cb3;
4364: douta=16'hbdb6;
4365: douta=16'hbdb6;
4366: douta=16'h8b8a;
4367: douta=16'h93ca;
4368: douta=16'hb46c;
4369: douta=16'hcd0d;
4370: douta=16'hcd2e;
4371: douta=16'hddd1;
4372: douta=16'hee75;
4373: douta=16'hee95;
4374: douta=16'he634;
4375: douta=16'hddd1;
4376: douta=16'hb4ad;
4377: douta=16'h9c0b;
4378: douta=16'h9c2c;
4379: douta=16'hbcef;
4380: douta=16'hb4ae;
4381: douta=16'hcd70;
4382: douta=16'hde13;
4383: douta=16'hde13;
4384: douta=16'hd591;
4385: douta=16'hcd71;
4386: douta=16'hbd11;
4387: douta=16'h9430;
4388: douta=16'h73b0;
4389: douta=16'h7390;
4390: douta=16'h6b71;
4391: douta=16'h4aef;
4392: douta=16'h3a4d;
4393: douta=16'h3a0b;
4394: douta=16'h528d;
4395: douta=16'h0883;
4396: douta=16'h10c4;
4397: douta=16'h10e4;
4398: douta=16'h10a4;
4399: douta=16'h1906;
4400: douta=16'h0884;
4401: douta=16'h1947;
4402: douta=16'h62ea;
4403: douta=16'h62e9;
4404: douta=16'h732b;
4405: douta=16'h5248;
4406: douta=16'h2966;
4407: douta=16'h6b6e;
4408: douta=16'h3a29;
4409: douta=16'h632e;
4410: douta=16'hb532;
4411: douta=16'h9559;
4412: douta=16'h7455;
4413: douta=16'h957a;
4414: douta=16'h8d18;
4415: douta=16'h63f4;
4416: douta=16'h84f7;
4417: douta=16'h9d7a;
4418: douta=16'h9599;
4419: douta=16'h8518;
4420: douta=16'h8d39;
4421: douta=16'h9d9a;
4422: douta=16'h8d39;
4423: douta=16'h9d9a;
4424: douta=16'h9d9a;
4425: douta=16'h959a;
4426: douta=16'h9dbb;
4427: douta=16'h957a;
4428: douta=16'h9dbb;
4429: douta=16'h9ddb;
4430: douta=16'h9d9a;
4431: douta=16'h6c36;
4432: douta=16'h957a;
4433: douta=16'ha46f;
4434: douta=16'h10e5;
4435: douta=16'h322c;
4436: douta=16'h84f8;
4437: douta=16'h9539;
4438: douta=16'h9d7a;
4439: douta=16'h9518;
4440: douta=16'h9559;
4441: douta=16'h957a;
4442: douta=16'h9dfc;
4443: douta=16'h9d9a;
4444: douta=16'h84b6;
4445: douta=16'h7c13;
4446: douta=16'h8d17;
4447: douta=16'h84d7;
4448: douta=16'h84d7;
4449: douta=16'h7456;
4450: douta=16'h6392;
4451: douta=16'h1925;
4452: douta=16'h2106;
4453: douta=16'h4313;
4454: douta=16'h5c78;
4455: douta=16'h6458;
4456: douta=16'h5bf6;
4457: douta=16'h74d9;
4458: douta=16'h74f9;
4459: douta=16'h7cf9;
4460: douta=16'h6c77;
4461: douta=16'h7cf9;
4462: douta=16'h7d19;
4463: douta=16'h7cf9;
4464: douta=16'h74b8;
4465: douta=16'h851a;
4466: douta=16'h6436;
4467: douta=16'h8d9b;
4468: douta=16'h6c77;
4469: douta=16'h8d5b;
4470: douta=16'h8d7b;
4471: douta=16'h7d1a;
4472: douta=16'h8d7b;
4473: douta=16'h7cf9;
4474: douta=16'h428d;
4475: douta=16'h63b1;
4476: douta=16'hb5d9;
4477: douta=16'h5b71;
4478: douta=16'h5aee;
4479: douta=16'ha557;
4480: douta=16'h32f2;
4481: douta=16'h3af2;
4482: douta=16'h5416;
4483: douta=16'h3b12;
4484: douta=16'h63f5;
4485: douta=16'h5bb4;
4486: douta=16'h6392;
4487: douta=16'h6392;
4488: douta=16'h7bf2;
4489: douta=16'ha536;
4490: douta=16'hc618;
4491: douta=16'h8411;
4492: douta=16'hc5f6;
4493: douta=16'h834a;
4494: douta=16'hb44b;
4495: douta=16'hb4ac;
4496: douta=16'hc4ed;
4497: douta=16'hd5b0;
4498: douta=16'hd5b0;
4499: douta=16'hee75;
4500: douta=16'hde13;
4501: douta=16'he634;
4502: douta=16'hd5b1;
4503: douta=16'hbcf0;
4504: douta=16'hac8d;
4505: douta=16'hb4ce;
4506: douta=16'hacae;
4507: douta=16'hc54f;
4508: douta=16'hcd71;
4509: douta=16'he634;
4510: douta=16'hee75;
4511: douta=16'hde13;
4512: douta=16'hd5d2;
4513: douta=16'hcd50;
4514: douta=16'hbd11;
4515: douta=16'ha471;
4516: douta=16'h8c31;
4517: douta=16'h8411;
4518: douta=16'h73d1;
4519: douta=16'h5b50;
4520: douta=16'h5b30;
4521: douta=16'h6372;
4522: douta=16'h18e5;
4523: douta=16'h2146;
4524: douta=16'h0862;
4525: douta=16'h10e4;
4526: douta=16'h10c4;
4527: douta=16'h10a3;
4528: douta=16'h1905;
4529: douta=16'h0042;
4530: douta=16'h08a5;
4531: douta=16'h840d;
4532: douta=16'hbd72;
4533: douta=16'h39a7;
4534: douta=16'h5269;
4535: douta=16'h630c;
4536: douta=16'h632d;
4537: douta=16'h2187;
4538: douta=16'h2146;
4539: douta=16'h7c95;
4540: douta=16'h8d38;
4541: douta=16'h84f8;
4542: douta=16'h9559;
4543: douta=16'h7c97;
4544: douta=16'h9559;
4545: douta=16'h7456;
4546: douta=16'h5bb2;
4547: douta=16'ha5ba;
4548: douta=16'h9579;
4549: douta=16'h9579;
4550: douta=16'h959a;
4551: douta=16'ha5da;
4552: douta=16'h9579;
4553: douta=16'h9d9a;
4554: douta=16'h9559;
4555: douta=16'ha5db;
4556: douta=16'ha5db;
4557: douta=16'ha5fb;
4558: douta=16'h7cd8;
4559: douta=16'h959a;
4560: douta=16'h8d39;
4561: douta=16'h94f6;
4562: douta=16'h2126;
4563: douta=16'h0042;
4564: douta=16'h957a;
4565: douta=16'h8d39;
4566: douta=16'h84d8;
4567: douta=16'h957a;
4568: douta=16'h84b7;
4569: douta=16'h9d9a;
4570: douta=16'h8518;
4571: douta=16'h9d99;
4572: douta=16'h8cd6;
4573: douta=16'h8c75;
4574: douta=16'h9539;
4575: douta=16'h7455;
4576: douta=16'h84b8;
4577: douta=16'h7cd8;
4578: douta=16'h31a7;
4579: douta=16'h10e5;
4580: douta=16'h426d;
4581: douta=16'h6478;
4582: douta=16'h7d3b;
4583: douta=16'h3b34;
4584: douta=16'h7d5c;
4585: douta=16'h53f6;
4586: douta=16'h5bf6;
4587: douta=16'h857b;
4588: douta=16'h855b;
4589: douta=16'h7498;
4590: douta=16'h74b8;
4591: douta=16'h7cf9;
4592: douta=16'h7cd9;
4593: douta=16'h7cd9;
4594: douta=16'h7cf9;
4595: douta=16'h8d5a;
4596: douta=16'h6c77;
4597: douta=16'h853a;
4598: douta=16'h7478;
4599: douta=16'h853a;
4600: douta=16'h855b;
4601: douta=16'h8d7b;
4602: douta=16'h39ca;
4603: douta=16'hbe3a;
4604: douta=16'h5330;
4605: douta=16'h9d16;
4606: douta=16'h0000;
4607: douta=16'h5310;
4608: douta=16'h2a4f;
4609: douta=16'h21ec;
4610: douta=16'h53d6;
4611: douta=16'h32f2;
4612: douta=16'h4b31;
4613: douta=16'h6416;
4614: douta=16'h4acf;
4615: douta=16'h8cd7;
4616: douta=16'h8453;
4617: douta=16'h8433;
4618: douta=16'hbdd7;
4619: douta=16'h9c93;
4620: douta=16'h7b0a;
4621: douta=16'h9c0b;
4622: douta=16'hc50e;
4623: douta=16'hc52e;
4624: douta=16'hd590;
4625: douta=16'he634;
4626: douta=16'he655;
4627: douta=16'he654;
4628: douta=16'hee96;
4629: douta=16'hd5d3;
4630: douta=16'hb4ad;
4631: douta=16'hb4ae;
4632: douta=16'h9c0c;
4633: douta=16'ha42d;
4634: douta=16'hbd0f;
4635: douta=16'hcd91;
4636: douta=16'hde13;
4637: douta=16'he654;
4638: douta=16'he654;
4639: douta=16'hde13;
4640: douta=16'hd5b3;
4641: douta=16'hc551;
4642: douta=16'hbd11;
4643: douta=16'h9451;
4644: douta=16'h9c72;
4645: douta=16'h8c73;
4646: douta=16'h8433;
4647: douta=16'h8c74;
4648: douta=16'h5352;
4649: douta=16'h9bca;
4650: douta=16'h39ea;
4651: douta=16'h2167;
4652: douta=16'h0042;
4653: douta=16'h1083;
4654: douta=16'h10c5;
4655: douta=16'h18e4;
4656: douta=16'h10e4;
4657: douta=16'h18e5;
4658: douta=16'h21a8;
4659: douta=16'h52cd;
4660: douta=16'h4a28;
4661: douta=16'h2946;
4662: douta=16'h3145;
4663: douta=16'h2945;
4664: douta=16'h7b6d;
4665: douta=16'h944f;
4666: douta=16'h630c;
4667: douta=16'h62ec;
4668: douta=16'h9559;
4669: douta=16'h7c96;
4670: douta=16'h84d7;
4671: douta=16'h8d39;
4672: douta=16'h7cb7;
4673: douta=16'h84d7;
4674: douta=16'h84d7;
4675: douta=16'h9579;
4676: douta=16'h7c96;
4677: douta=16'h84b6;
4678: douta=16'h9d9a;
4679: douta=16'h9d99;
4680: douta=16'ha5da;
4681: douta=16'ha5ba;
4682: douta=16'h9579;
4683: douta=16'ha5da;
4684: douta=16'hae1b;
4685: douta=16'h9d9a;
4686: douta=16'h9d9a;
4687: douta=16'ha5da;
4688: douta=16'h8d39;
4689: douta=16'h8d39;
4690: douta=16'hac6d;
4691: douta=16'h10c4;
4692: douta=16'ha5fc;
4693: douta=16'h84d8;
4694: douta=16'h8d5a;
4695: douta=16'h8d39;
4696: douta=16'h9d59;
4697: douta=16'h7c76;
4698: douta=16'h7c55;
4699: douta=16'h9d58;
4700: douta=16'ha578;
4701: douta=16'h9d37;
4702: douta=16'h8d18;
4703: douta=16'h8d7a;
4704: douta=16'h959b;
4705: douta=16'h851a;
4706: douta=16'h3167;
4707: douta=16'h10a4;
4708: douta=16'h6457;
4709: douta=16'h74b9;
4710: douta=16'h6cb9;
4711: douta=16'h855b;
4712: douta=16'h7d1b;
4713: douta=16'h53d5;
4714: douta=16'h855b;
4715: douta=16'h6437;
4716: douta=16'h53d4;
4717: douta=16'h6c98;
4718: douta=16'h853a;
4719: douta=16'h7478;
4720: douta=16'h8d7b;
4721: douta=16'h8d5b;
4722: douta=16'h84f9;
4723: douta=16'h851a;
4724: douta=16'h855a;
4725: douta=16'h851a;
4726: douta=16'h851a;
4727: douta=16'h7457;
4728: douta=16'h95bc;
4729: douta=16'h6bf3;
4730: douta=16'h84d6;
4731: douta=16'h8cf7;
4732: douta=16'h4b11;
4733: douta=16'h7413;
4734: douta=16'h7454;
4735: douta=16'h8c95;
4736: douta=16'h324d;
4737: douta=16'h21ed;
4738: douta=16'h19cc;
4739: douta=16'h32f2;
4740: douta=16'h5352;
4741: douta=16'h74b8;
4742: douta=16'h6392;
4743: douta=16'h8497;
4744: douta=16'h8c95;
4745: douta=16'h5b30;
4746: douta=16'h8c52;
4747: douta=16'h8bcb;
4748: douta=16'h938b;
4749: douta=16'hbcad;
4750: douta=16'hcd4f;
4751: douta=16'hcd6f;
4752: douta=16'he633;
4753: douta=16'hee96;
4754: douta=16'he634;
4755: douta=16'heeb6;
4756: douta=16'hddf2;
4757: douta=16'hc50e;
4758: douta=16'hb4ce;
4759: douta=16'h8b8a;
4760: douta=16'ha42d;
4761: douta=16'hc54f;
4762: douta=16'hd5b0;
4763: douta=16'hde13;
4764: douta=16'hee75;
4765: douta=16'hde14;
4766: douta=16'hde33;
4767: douta=16'he613;
4768: douta=16'hcd72;
4769: douta=16'hbcf1;
4770: douta=16'hb4d1;
4771: douta=16'h8c12;
4772: douta=16'h8412;
4773: douta=16'h8c33;
4774: douta=16'h73f2;
4775: douta=16'h5b2f;
4776: douta=16'h8b28;
4777: douta=16'h9c2e;
4778: douta=16'h5aac;
4779: douta=16'h31ea;
4780: douta=16'h10e5;
4781: douta=16'h1906;
4782: douta=16'h10a4;
4783: douta=16'h10e4;
4784: douta=16'h10a4;
4785: douta=16'h10e4;
4786: douta=16'h1906;
4787: douta=16'h0000;
4788: douta=16'h6bb0;
4789: douta=16'h940d;
4790: douta=16'haccf;
4791: douta=16'h0861;
4792: douta=16'h9cd1;
4793: douta=16'h8c0d;
4794: douta=16'h83ee;
4795: douta=16'h8bef;
4796: douta=16'h8cf8;
4797: douta=16'h8d39;
4798: douta=16'h9d9a;
4799: douta=16'h8d38;
4800: douta=16'h8517;
4801: douta=16'h7c96;
4802: douta=16'h9579;
4803: douta=16'h9538;
4804: douta=16'h8d38;
4805: douta=16'h8d58;
4806: douta=16'h84f8;
4807: douta=16'h9579;
4808: douta=16'h8d59;
4809: douta=16'ha5ba;
4810: douta=16'h8d39;
4811: douta=16'h7cb7;
4812: douta=16'ha5da;
4813: douta=16'h959a;
4814: douta=16'h9d9a;
4815: douta=16'ha5ba;
4816: douta=16'h9d7a;
4817: douta=16'h9579;
4818: douta=16'hc4ee;
4819: douta=16'h2926;
4820: douta=16'h29ca;
4821: douta=16'h9559;
4822: douta=16'h9dba;
4823: douta=16'h6c35;
4824: douta=16'h7c96;
4825: douta=16'h84d7;
4826: douta=16'h84b6;
4827: douta=16'h7c13;
4828: douta=16'h7c33;
4829: douta=16'h8cb6;
4830: douta=16'h7cb7;
4831: douta=16'h7497;
4832: douta=16'h959a;
4833: douta=16'h7476;
4834: douta=16'h0884;
4835: douta=16'h31c8;
4836: douta=16'h74d9;
4837: douta=16'h7d3a;
4838: douta=16'h6436;
4839: douta=16'h6457;
4840: douta=16'h74d9;
4841: douta=16'h7cd9;
4842: douta=16'h9e1d;
4843: douta=16'h7cd9;
4844: douta=16'h7498;
4845: douta=16'h74fa;
4846: douta=16'h53f6;
4847: douta=16'h853a;
4848: douta=16'h8d5a;
4849: douta=16'h6c36;
4850: douta=16'h6c57;
4851: douta=16'h8d7a;
4852: douta=16'h851a;
4853: douta=16'h6c77;
4854: douta=16'h959c;
4855: douta=16'h7cb8;
4856: douta=16'h8d9b;
4857: douta=16'h6391;
4858: douta=16'h7454;
4859: douta=16'h9d58;
4860: douta=16'h8475;
4861: douta=16'h73f3;
4862: douta=16'hadb8;
4863: douta=16'h5351;
4864: douta=16'h2126;
4865: douta=16'h2a4f;
4866: douta=16'h4bb6;
4867: douta=16'h2a6f;
4868: douta=16'h5bb4;
4869: douta=16'h7cd9;
4870: douta=16'h5b93;
4871: douta=16'h5351;
4872: douta=16'h94f6;
4873: douta=16'h8454;
4874: douta=16'h6b70;
4875: douta=16'h8bab;
4876: douta=16'ha40b;
4877: douta=16'hcd2e;
4878: douta=16'hddf1;
4879: douta=16'hddf2;
4880: douta=16'heeb6;
4881: douta=16'heeb6;
4882: douta=16'he654;
4883: douta=16'hc50e;
4884: douta=16'hcd70;
4885: douta=16'hc4ee;
4886: douta=16'h8baa;
4887: douta=16'h9c0c;
4888: douta=16'hc52f;
4889: douta=16'hd5b1;
4890: douta=16'hde13;
4891: douta=16'he654;
4892: douta=16'he675;
4893: douta=16'hde13;
4894: douta=16'hddf3;
4895: douta=16'hd5b2;
4896: douta=16'hc552;
4897: douta=16'ha491;
4898: douta=16'h9c72;
4899: douta=16'h6371;
4900: douta=16'h9472;
4901: douta=16'h6b2e;
4902: douta=16'h73d1;
4903: douta=16'h7309;
4904: douta=16'he613;
4905: douta=16'h9c2e;
4906: douta=16'h734d;
4907: douta=16'h5acd;
4908: douta=16'h29c9;
4909: douta=16'h2126;
4910: douta=16'h0883;
4911: douta=16'h4a6b;
4912: douta=16'h10e4;
4913: douta=16'h10e4;
4914: douta=16'h18a4;
4915: douta=16'h10a4;
4916: douta=16'h0863;
4917: douta=16'h6bd2;
4918: douta=16'h0884;
4919: douta=16'h7bad;
4920: douta=16'h1125;
4921: douta=16'h39e7;
4922: douta=16'h5269;
4923: douta=16'h732a;
4924: douta=16'ha5fc;
4925: douta=16'h8d39;
4926: douta=16'h957a;
4927: douta=16'h8d39;
4928: douta=16'h8d18;
4929: douta=16'h9d79;
4930: douta=16'h8d38;
4931: douta=16'h8d38;
4932: douta=16'h8d18;
4933: douta=16'h84b7;
4934: douta=16'h8d59;
4935: douta=16'h8539;
4936: douta=16'h6415;
4937: douta=16'h84d8;
4938: douta=16'h84f9;
4939: douta=16'h959a;
4940: douta=16'h9d79;
4941: douta=16'hadfa;
4942: douta=16'ha5ba;
4943: douta=16'hb61b;
4944: douta=16'h9d59;
4945: douta=16'h9d9a;
4946: douta=16'h8d39;
4947: douta=16'hff37;
4948: douta=16'h0043;
4949: douta=16'h8d38;
4950: douta=16'h9d9a;
4951: douta=16'h84f8;
4952: douta=16'h84b6;
4953: douta=16'hb61a;
4954: douta=16'h7413;
4955: douta=16'h73f2;
4956: douta=16'h7c55;
4957: douta=16'h9559;
4958: douta=16'h957b;
4959: douta=16'h7cd9;
4960: douta=16'h8d7c;
4961: douta=16'h1905;
4962: douta=16'h29c9;
4963: douta=16'h3a2b;
4964: douta=16'h5351;
4965: douta=16'h7cb8;
4966: douta=16'h7cf9;
4967: douta=16'h84f9;
4968: douta=16'h853a;
4969: douta=16'h7cb9;
4970: douta=16'h855a;
4971: douta=16'h857b;
4972: douta=16'h9ddc;
4973: douta=16'h8d7b;
4974: douta=16'h8d5a;
4975: douta=16'h8d9c;
4976: douta=16'h5bf6;
4977: douta=16'h8d5b;
4978: douta=16'h7d5a;
4979: douta=16'h8d5b;
4980: douta=16'h6436;
4981: douta=16'h8d3a;
4982: douta=16'h7cd9;
4983: douta=16'h7cd9;
4984: douta=16'h5bf5;
4985: douta=16'h7c56;
4986: douta=16'h2a2d;
4987: douta=16'h6c35;
4988: douta=16'hb65c;
4989: douta=16'h0800;
4990: douta=16'h84b6;
4991: douta=16'h9537;
4992: douta=16'h18a4;
4993: douta=16'h2250;
4994: douta=16'h4374;
4995: douta=16'h32d1;
4996: douta=16'h5394;
4997: douta=16'h5bb4;
4998: douta=16'h6c36;
4999: douta=16'h7435;
5000: douta=16'h8454;
5001: douta=16'h94b5;
5002: douta=16'h93ca;
5003: douta=16'ha42c;
5004: douta=16'hc4cd;
5005: douta=16'hd570;
5006: douta=16'he654;
5007: douta=16'heed7;
5008: douta=16'he654;
5009: douta=16'hddd2;
5010: douta=16'hde13;
5011: douta=16'hc52f;
5012: douta=16'hc52f;
5013: douta=16'h8b69;
5014: douta=16'hac6d;
5015: douta=16'hb4ed;
5016: douta=16'hd5f2;
5017: douta=16'he655;
5018: douta=16'he654;
5019: douta=16'heeb6;
5020: douta=16'he675;
5021: douta=16'he654;
5022: douta=16'hddd2;
5023: douta=16'hbd10;
5024: douta=16'h9c51;
5025: douta=16'h9c72;
5026: douta=16'h8412;
5027: douta=16'h73d1;
5028: douta=16'h31ea;
5029: douta=16'h4a6b;
5030: douta=16'hac2c;
5031: douta=16'hcd2e;
5032: douta=16'he634;
5033: douta=16'hb48d;
5034: douta=16'h7b6e;
5035: douta=16'h630e;
5036: douta=16'h52ee;
5037: douta=16'h322c;
5038: douta=16'h29a9;
5039: douta=16'h1906;
5040: douta=16'h42ad;
5041: douta=16'h10a3;
5042: douta=16'h18e5;
5043: douta=16'h10a4;
5044: douta=16'h1083;
5045: douta=16'h29a8;
5046: douta=16'h1926;
5047: douta=16'h1926;
5048: douta=16'hd633;
5049: douta=16'h8c2e;
5050: douta=16'h10a4;
5051: douta=16'h31a6;
5052: douta=16'h5aaa;
5053: douta=16'h7cb7;
5054: douta=16'h9579;
5055: douta=16'h9559;
5056: douta=16'h9579;
5057: douta=16'h8d38;
5058: douta=16'h8d38;
5059: douta=16'h8d18;
5060: douta=16'h8d39;
5061: douta=16'h8d58;
5062: douta=16'h9559;
5063: douta=16'h9559;
5064: douta=16'h8518;
5065: douta=16'h9559;
5066: douta=16'h957a;
5067: douta=16'h8518;
5068: douta=16'h8d39;
5069: douta=16'h9d9a;
5070: douta=16'h8d18;
5071: douta=16'h8d39;
5072: douta=16'h9d9a;
5073: douta=16'h9d9a;
5074: douta=16'h9d99;
5075: douta=16'had34;
5076: douta=16'he590;
5077: douta=16'h1106;
5078: douta=16'h7cb7;
5079: douta=16'h9d79;
5080: douta=16'h9558;
5081: douta=16'h9d58;
5082: douta=16'h94f6;
5083: douta=16'h9d16;
5084: douta=16'h7c35;
5085: douta=16'h6cb8;
5086: douta=16'h6457;
5087: douta=16'h7d5c;
5088: douta=16'h2125;
5089: douta=16'h322c;
5090: douta=16'h1107;
5091: douta=16'h7d3a;
5092: douta=16'h8d7b;
5093: douta=16'h8d5a;
5094: douta=16'h6415;
5095: douta=16'h7498;
5096: douta=16'h855a;
5097: douta=16'h853a;
5098: douta=16'h7498;
5099: douta=16'h8d5a;
5100: douta=16'h8519;
5101: douta=16'h855a;
5102: douta=16'h853a;
5103: douta=16'h853b;
5104: douta=16'h74d9;
5105: douta=16'h855a;
5106: douta=16'h5c16;
5107: douta=16'h7cd9;
5108: douta=16'h7cf9;
5109: douta=16'h7498;
5110: douta=16'h6457;
5111: douta=16'h6cda;
5112: douta=16'h630e;
5113: douta=16'h7414;
5114: douta=16'h5310;
5115: douta=16'h7cb7;
5116: douta=16'hb69f;
5117: douta=16'h5330;
5118: douta=16'h7434;
5119: douta=16'h7c95;
5120: douta=16'h1062;
5121: douta=16'h4394;
5122: douta=16'h32b0;
5123: douta=16'h2a4f;
5124: douta=16'h6436;
5125: douta=16'h5393;
5126: douta=16'h63d4;
5127: douta=16'h6bd3;
5128: douta=16'h7c55;
5129: douta=16'h732c;
5130: douta=16'hac4c;
5131: douta=16'hac6c;
5132: douta=16'hcd4f;
5133: douta=16'hd5d0;
5134: douta=16'heeb6;
5135: douta=16'heeb6;
5136: douta=16'hee75;
5137: douta=16'he654;
5138: douta=16'hd591;
5139: douta=16'hb46c;
5140: douta=16'h8b69;
5141: douta=16'h9c2b;
5142: douta=16'hbcee;
5143: douta=16'hcd6f;
5144: douta=16'he655;
5145: douta=16'he675;
5146: douta=16'hee96;
5147: douta=16'he675;
5148: douta=16'he654;
5149: douta=16'hddd2;
5150: douta=16'hcd90;
5151: douta=16'ha450;
5152: douta=16'h8c11;
5153: douta=16'h7bd1;
5154: douta=16'h7b6f;
5155: douta=16'h630e;
5156: douta=16'h524a;
5157: douta=16'h9389;
5158: douta=16'h938b;
5159: douta=16'hddf2;
5160: douta=16'he613;
5161: douta=16'hd52f;
5162: douta=16'ha40e;
5163: douta=16'h6b2e;
5164: douta=16'h632f;
5165: douta=16'h5330;
5166: douta=16'h42cf;
5167: douta=16'h322c;
5168: douta=16'h2168;
5169: douta=16'h424c;
5170: douta=16'h10a4;
5171: douta=16'h18e5;
5172: douta=16'h10e4;
5173: douta=16'h1905;
5174: douta=16'h1925;
5175: douta=16'h2126;
5176: douta=16'h0043;
5177: douta=16'h2167;
5178: douta=16'h2967;
5179: douta=16'h2166;
5180: douta=16'h62cb;
5181: douta=16'h4aae;
5182: douta=16'h8d18;
5183: douta=16'h84d7;
5184: douta=16'h7cb6;
5185: douta=16'ha5fb;
5186: douta=16'h9599;
5187: douta=16'h8d18;
5188: douta=16'h84f7;
5189: douta=16'h84f8;
5190: douta=16'h84d7;
5191: douta=16'h8d39;
5192: douta=16'h8d18;
5193: douta=16'h8d38;
5194: douta=16'h84b7;
5195: douta=16'h84d7;
5196: douta=16'h9559;
5197: douta=16'h9d9a;
5198: douta=16'h9559;
5199: douta=16'h8d19;
5200: douta=16'h8d39;
5201: douta=16'h8d59;
5202: douta=16'h8d59;
5203: douta=16'h9d99;
5204: douta=16'h838e;
5205: douta=16'h6b0f;
5206: douta=16'h1948;
5207: douta=16'h0001;
5208: douta=16'h42cf;
5209: douta=16'hadfb;
5210: douta=16'h5aea;
5211: douta=16'h19ab;
5212: douta=16'h54fb;
5213: douta=16'h4311;
5214: douta=16'h2082;
5215: douta=16'h4a09;
5216: douta=16'h42d0;
5217: douta=16'h1105;
5218: douta=16'h857b;
5219: douta=16'h7cd9;
5220: douta=16'h7cf9;
5221: douta=16'h8519;
5222: douta=16'h957a;
5223: douta=16'h9dbc;
5224: douta=16'h8d5b;
5225: douta=16'h84d9;
5226: douta=16'h853a;
5227: douta=16'h8d7b;
5228: douta=16'h8d5a;
5229: douta=16'h8d19;
5230: douta=16'h8d5a;
5231: douta=16'h8d5a;
5232: douta=16'h7cf9;
5233: douta=16'h853a;
5234: douta=16'h851a;
5235: douta=16'h7d1a;
5236: douta=16'h6478;
5237: douta=16'h6c57;
5238: douta=16'h6cb9;
5239: douta=16'h6a46;
5240: douta=16'h4372;
5241: douta=16'h84b6;
5242: douta=16'h84b8;
5243: douta=16'h5bf3;
5244: douta=16'h4a28;
5245: douta=16'h9539;
5246: douta=16'h7c54;
5247: douta=16'h638f;
5248: douta=16'h18e4;
5249: douta=16'h328f;
5250: douta=16'h2a6f;
5251: douta=16'h4374;
5252: douta=16'h6415;
5253: douta=16'h84d8;
5254: douta=16'h7c77;
5255: douta=16'h5b51;
5256: douta=16'h5b71;
5257: douta=16'h9bca;
5258: douta=16'hbccd;
5259: douta=16'hc4ed;
5260: douta=16'hddd1;
5261: douta=16'he633;
5262: douta=16'hee96;
5263: douta=16'heeb6;
5264: douta=16'he654;
5265: douta=16'hd5b1;
5266: douta=16'hbd0f;
5267: douta=16'h8308;
5268: douta=16'h93ca;
5269: douta=16'hbccd;
5270: douta=16'hc52e;
5271: douta=16'hde12;
5272: douta=16'hee96;
5273: douta=16'hee95;
5274: douta=16'heeb6;
5275: douta=16'he613;
5276: douta=16'hddd2;
5277: douta=16'hc530;
5278: douta=16'hb4af;
5279: douta=16'h9431;
5280: douta=16'h8412;
5281: douta=16'h630e;
5282: douta=16'h734e;
5283: douta=16'h49e8;
5284: douta=16'ha40b;
5285: douta=16'h9bcb;
5286: douta=16'hcd6f;
5287: douta=16'he654;
5288: douta=16'he5f2;
5289: douta=16'hc4ee;
5290: douta=16'ha40d;
5291: douta=16'h7b4d;
5292: douta=16'h6b4f;
5293: douta=16'h6b71;
5294: douta=16'h5331;
5295: douta=16'h3a8e;
5296: douta=16'h29eb;
5297: douta=16'h2168;
5298: douta=16'h4ace;
5299: douta=16'h10e4;
5300: douta=16'h10c4;
5301: douta=16'h10a4;
5302: douta=16'h10c4;
5303: douta=16'h1905;
5304: douta=16'h29a8;
5305: douta=16'h6b90;
5306: douta=16'h83ee;
5307: douta=16'h5269;
5308: douta=16'h18e5;
5309: douta=16'h6b2b;
5310: douta=16'h6c13;
5311: douta=16'h8d38;
5312: douta=16'h84d7;
5313: douta=16'h84b7;
5314: douta=16'h9579;
5315: douta=16'h8d39;
5316: douta=16'ha5da;
5317: douta=16'h9558;
5318: douta=16'h7cb7;
5319: douta=16'h7496;
5320: douta=16'h84f7;
5321: douta=16'h84d7;
5322: douta=16'h8d18;
5323: douta=16'h8d39;
5324: douta=16'h84d7;
5325: douta=16'h8d18;
5326: douta=16'h8d39;
5327: douta=16'h8d18;
5328: douta=16'h957a;
5329: douta=16'h84f8;
5330: douta=16'h7cd7;
5331: douta=16'h9559;
5332: douta=16'h7cd7;
5333: douta=16'h9db9;
5334: douta=16'h6bd3;
5335: douta=16'h1989;
5336: douta=16'h21aa;
5337: douta=16'h10e5;
5338: douta=16'h10c5;
5339: douta=16'h1905;
5340: douta=16'h3186;
5341: douta=16'h834c;
5342: douta=16'h832b;
5343: douta=16'h63f4;
5344: douta=16'h4a8d;
5345: douta=16'h853b;
5346: douta=16'h7cb8;
5347: douta=16'h6c37;
5348: douta=16'h959b;
5349: douta=16'h7cb8;
5350: douta=16'h7cb8;
5351: douta=16'h8d5a;
5352: douta=16'ha5fc;
5353: douta=16'h8d5b;
5354: douta=16'h8d5b;
5355: douta=16'h95bc;
5356: douta=16'h84d9;
5357: douta=16'h74b8;
5358: douta=16'h74b8;
5359: douta=16'h8d7b;
5360: douta=16'h851a;
5361: douta=16'h5bf5;
5362: douta=16'h853a;
5363: douta=16'h851a;
5364: douta=16'h74d9;
5365: douta=16'h857b;
5366: douta=16'h73b1;
5367: douta=16'h63d4;
5368: douta=16'h63d3;
5369: douta=16'h3965;
5370: douta=16'h7d3b;
5371: douta=16'h6c56;
5372: douta=16'h2924;
5373: douta=16'h84b6;
5374: douta=16'h3a4c;
5375: douta=16'h1083;
5376: douta=16'h2104;
5377: douta=16'h29ca;
5378: douta=16'h32b0;
5379: douta=16'h4374;
5380: douta=16'h53b4;
5381: douta=16'h5351;
5382: douta=16'h5bb4;
5383: douta=16'h6bb2;
5384: douta=16'h7c55;
5385: douta=16'hbcad;
5386: douta=16'hc50e;
5387: douta=16'hcd4f;
5388: douta=16'he634;
5389: douta=16'hee95;
5390: douta=16'hee75;
5391: douta=16'hddf1;
5392: douta=16'he633;
5393: douta=16'hc4ee;
5394: douta=16'ha40b;
5395: douta=16'hac6d;
5396: douta=16'hac4c;
5397: douta=16'hbcee;
5398: douta=16'hddd1;
5399: douta=16'he654;
5400: douta=16'hee96;
5401: douta=16'hee95;
5402: douta=16'he654;
5403: douta=16'he654;
5404: douta=16'hcd50;
5405: douta=16'hac8f;
5406: douta=16'h8c10;
5407: douta=16'h8bf1;
5408: douta=16'h6b2e;
5409: douta=16'h6b0d;
5410: douta=16'h2904;
5411: douta=16'h93ca;
5412: douta=16'ha46c;
5413: douta=16'hd5b1;
5414: douta=16'hee75;
5415: douta=16'he655;
5416: douta=16'hdd90;
5417: douta=16'hc4cd;
5418: douta=16'ha40d;
5419: douta=16'h9bef;
5420: douta=16'h8bd0;
5421: douta=16'h6370;
5422: douta=16'h6371;
5423: douta=16'h42cf;
5424: douta=16'h428e;
5425: douta=16'h322c;
5426: douta=16'h29ea;
5427: douta=16'h530e;
5428: douta=16'h18c4;
5429: douta=16'h10a4;
5430: douta=16'h08a3;
5431: douta=16'h10c4;
5432: douta=16'h10e4;
5433: douta=16'h0021;
5434: douta=16'h6bf1;
5435: douta=16'had33;
5436: douta=16'ha4b0;
5437: douta=16'had31;
5438: douta=16'h62aa;
5439: douta=16'h7cb7;
5440: douta=16'h7455;
5441: douta=16'h84d7;
5442: douta=16'h8d18;
5443: douta=16'h84b7;
5444: douta=16'h84f7;
5445: douta=16'h7cb7;
5446: douta=16'h84f7;
5447: douta=16'h84b6;
5448: douta=16'h9dba;
5449: douta=16'h84b6;
5450: douta=16'h957a;
5451: douta=16'h9d79;
5452: douta=16'h959a;
5453: douta=16'h9d79;
5454: douta=16'h84b6;
5455: douta=16'h84d7;
5456: douta=16'ha5bb;
5457: douta=16'h8d18;
5458: douta=16'h8518;
5459: douta=16'h8d19;
5460: douta=16'h8518;
5461: douta=16'h955a;
5462: douta=16'h8519;
5463: douta=16'h634f;
5464: douta=16'h52ee;
5465: douta=16'h4b51;
5466: douta=16'h1927;
5467: douta=16'h5acd;
5468: douta=16'h6b71;
5469: douta=16'h4a6e;
5470: douta=16'h5ace;
5471: douta=16'ha63d;
5472: douta=16'h9559;
5473: douta=16'h9ddb;
5474: douta=16'h9ddb;
5475: douta=16'h8d5a;
5476: douta=16'hae1c;
5477: douta=16'h7cb8;
5478: douta=16'h7cd8;
5479: douta=16'h8519;
5480: douta=16'h8d7a;
5481: douta=16'h7cd8;
5482: douta=16'h7cb9;
5483: douta=16'h8d9b;
5484: douta=16'h9d9b;
5485: douta=16'h959a;
5486: douta=16'h959b;
5487: douta=16'h7498;
5488: douta=16'h7498;
5489: douta=16'h853a;
5490: douta=16'h7cf9;
5491: douta=16'h7d19;
5492: douta=16'h6477;
5493: douta=16'h6aec;
5494: douta=16'h5bb3;
5495: douta=16'h63f5;
5496: douta=16'h84f9;
5497: douta=16'h9559;
5498: douta=16'h9517;
5499: douta=16'h5164;
5500: douta=16'h3b30;
5501: douta=16'h84d7;
5502: douta=16'h7cb7;
5503: douta=16'h10a3;
5504: douta=16'h2926;
5505: douta=16'h31ca;
5506: douta=16'h3312;
5507: douta=16'h4bb5;
5508: douta=16'h4b53;
5509: douta=16'h63d4;
5510: douta=16'h6c36;
5511: douta=16'h6392;
5512: douta=16'h8d18;
5513: douta=16'hc4ed;
5514: douta=16'hd56f;
5515: douta=16'hde13;
5516: douta=16'hee95;
5517: douta=16'hee95;
5518: douta=16'he654;
5519: douta=16'hd5b0;
5520: douta=16'hac4d;
5521: douta=16'hbcee;
5522: douta=16'hb4ae;
5523: douta=16'hb4cd;
5524: douta=16'hbcee;
5525: douta=16'hde33;
5526: douta=16'he634;
5527: douta=16'he675;
5528: douta=16'heeb6;
5529: douta=16'hee75;
5530: douta=16'he654;
5531: douta=16'hd590;
5532: douta=16'hbcb0;
5533: douta=16'h83d0;
5534: douta=16'h7370;
5535: douta=16'h734f;
5536: douta=16'h5aaa;
5537: douta=16'h2925;
5538: douta=16'ha3eb;
5539: douta=16'hcd2f;
5540: douta=16'he613;
5541: douta=16'hee95;
5542: douta=16'hee75;
5543: douta=16'hee54;
5544: douta=16'hcd0f;
5545: douta=16'hc4cf;
5546: douta=16'hac4e;
5547: douta=16'h93ce;
5548: douta=16'h8c10;
5549: douta=16'h7bf2;
5550: douta=16'h6bb2;
5551: douta=16'h5b91;
5552: douta=16'h42ce;
5553: douta=16'h29cb;
5554: douta=16'h322c;
5555: douta=16'h31eb;
5556: douta=16'h3a4c;
5557: douta=16'h1905;
5558: douta=16'h1927;
5559: douta=16'h2147;
5560: douta=16'h1906;
5561: douta=16'h18e5;
5562: douta=16'h18e5;
5563: douta=16'h10e4;
5564: douta=16'h0022;
5565: douta=16'h6b6d;
5566: douta=16'h83ee;
5567: douta=16'h8bed;
5568: douta=16'h8518;
5569: douta=16'h7cb7;
5570: douta=16'h8d38;
5571: douta=16'h84f8;
5572: douta=16'h7476;
5573: douta=16'h63f4;
5574: douta=16'h8d18;
5575: douta=16'h8d38;
5576: douta=16'h7c96;
5577: douta=16'h8d18;
5578: douta=16'h9599;
5579: douta=16'hbe7c;
5580: douta=16'h84d8;
5581: douta=16'h8d39;
5582: douta=16'h8d39;
5583: douta=16'h9559;
5584: douta=16'h9559;
5585: douta=16'h8d39;
5586: douta=16'h8d18;
5587: douta=16'h8d18;
5588: douta=16'h7476;
5589: douta=16'h957a;
5590: douta=16'h8518;
5591: douta=16'h9d9a;
5592: douta=16'h8d39;
5593: douta=16'h853a;
5594: douta=16'h49e6;
5595: douta=16'h2188;
5596: douta=16'hae3e;
5597: douta=16'h8d59;
5598: douta=16'h7cf8;
5599: douta=16'h959a;
5600: douta=16'h8d79;
5601: douta=16'h8539;
5602: douta=16'h9dbb;
5603: douta=16'h7cf8;
5604: douta=16'ha5db;
5605: douta=16'h9dbb;
5606: douta=16'h959b;
5607: douta=16'h959a;
5608: douta=16'h7498;
5609: douta=16'h8d3a;
5610: douta=16'h959b;
5611: douta=16'h855a;
5612: douta=16'h7478;
5613: douta=16'h7498;
5614: douta=16'h8d3a;
5615: douta=16'h853a;
5616: douta=16'h853a;
5617: douta=16'h95bc;
5618: douta=16'h7d19;
5619: douta=16'h74b8;
5620: douta=16'h52ac;
5621: douta=16'h32ae;
5622: douta=16'h6415;
5623: douta=16'hae1c;
5624: douta=16'h6c76;
5625: douta=16'h4b33;
5626: douta=16'h8d18;
5627: douta=16'h0000;
5628: douta=16'h7c96;
5629: douta=16'h61e4;
5630: douta=16'h64d9;
5631: douta=16'h0882;
5632: douta=16'h3146;
5633: douta=16'h2126;
5634: douta=16'h3b33;
5635: douta=16'h4333;
5636: douta=16'h4b53;
5637: douta=16'h4b11;
5638: douta=16'h5bb4;
5639: douta=16'h63b3;
5640: douta=16'h63f4;
5641: douta=16'hc50d;
5642: douta=16'hcd70;
5643: douta=16'he654;
5644: douta=16'heeb6;
5645: douta=16'he675;
5646: douta=16'hd5b1;
5647: douta=16'hc4cf;
5648: douta=16'h938a;
5649: douta=16'ha42c;
5650: douta=16'hb4ad;
5651: douta=16'hd591;
5652: douta=16'hddf2;
5653: douta=16'hee95;
5654: douta=16'hddf2;
5655: douta=16'heeb6;
5656: douta=16'hee95;
5657: douta=16'hee54;
5658: douta=16'hddd1;
5659: douta=16'hd550;
5660: douta=16'h9c10;
5661: douta=16'h7bb0;
5662: douta=16'h62ed;
5663: douta=16'h5a6a;
5664: douta=16'h2904;
5665: douta=16'hb46c;
5666: douta=16'hcd2d;
5667: douta=16'he613;
5668: douta=16'hee96;
5669: douta=16'hee75;
5670: douta=16'hee75;
5671: douta=16'hddd2;
5672: douta=16'hcd0f;
5673: douta=16'hbccf;
5674: douta=16'hb46e;
5675: douta=16'h9410;
5676: douta=16'h8c31;
5677: douta=16'h8c73;
5678: douta=16'h7c13;
5679: douta=16'h7434;
5680: douta=16'h6bd2;
5681: douta=16'h6392;
5682: douta=16'h0909;
5683: douta=16'h4b0e;
5684: douta=16'h4a8e;
5685: douta=16'h0042;
5686: douta=16'h1905;
5687: douta=16'h10a4;
5688: douta=16'h10a4;
5689: douta=16'h1905;
5690: douta=16'h18e5;
5691: douta=16'h1084;
5692: douta=16'h18c4;
5693: douta=16'h10e4;
5694: douta=16'h736d;
5695: douta=16'hde97;
5696: douta=16'h4a8c;
5697: douta=16'h9d7a;
5698: douta=16'h7cb7;
5699: douta=16'h7cb7;
5700: douta=16'h959a;
5701: douta=16'h9599;
5702: douta=16'h84f8;
5703: douta=16'h84d6;
5704: douta=16'h6c14;
5705: douta=16'h8d18;
5706: douta=16'h8d18;
5707: douta=16'h84d7;
5708: douta=16'h7455;
5709: douta=16'ha5db;
5710: douta=16'h9dba;
5711: douta=16'h8d19;
5712: douta=16'h9559;
5713: douta=16'h84d7;
5714: douta=16'h84b7;
5715: douta=16'h8518;
5716: douta=16'h84f8;
5717: douta=16'h957a;
5718: douta=16'h7497;
5719: douta=16'h84f8;
5720: douta=16'h8d7a;
5721: douta=16'h8d19;
5722: douta=16'h8b6b;
5723: douta=16'h1882;
5724: douta=16'h7cb8;
5725: douta=16'h9dbb;
5726: douta=16'h95bb;
5727: douta=16'h959a;
5728: douta=16'h8d18;
5729: douta=16'h8d59;
5730: douta=16'h74b8;
5731: douta=16'h9dbb;
5732: douta=16'h8d7a;
5733: douta=16'h95bb;
5734: douta=16'h957a;
5735: douta=16'h959b;
5736: douta=16'h959a;
5737: douta=16'h957a;
5738: douta=16'h7477;
5739: douta=16'h7cd8;
5740: douta=16'h959b;
5741: douta=16'h8d3a;
5742: douta=16'h9d9a;
5743: douta=16'h7477;
5744: douta=16'h7cf9;
5745: douta=16'h8d7b;
5746: douta=16'h8d5b;
5747: douta=16'h632e;
5748: douta=16'h5921;
5749: douta=16'h3af1;
5750: douta=16'h6c56;
5751: douta=16'h6c57;
5752: douta=16'h8d39;
5753: douta=16'h4311;
5754: douta=16'h84fa;
5755: douta=16'h63f4;
5756: douta=16'h5bf4;
5757: douta=16'h7456;
5758: douta=16'h7477;
5759: douta=16'h5a25;
5760: douta=16'h3145;
5761: douta=16'h1083;
5762: douta=16'h32d1;
5763: douta=16'h32b1;
5764: douta=16'h53b5;
5765: douta=16'h7456;
5766: douta=16'h7cb8;
5767: douta=16'h6372;
5768: douta=16'h8496;
5769: douta=16'hbcef;
5770: douta=16'hddf3;
5771: douta=16'hee76;
5772: douta=16'hee95;
5773: douta=16'he613;
5774: douta=16'hcd70;
5775: douta=16'h7b07;
5776: douta=16'hb48d;
5777: douta=16'hbcee;
5778: douta=16'hd613;
5779: douta=16'hd5d3;
5780: douta=16'he675;
5781: douta=16'hddf3;
5782: douta=16'heeb7;
5783: douta=16'hee95;
5784: douta=16'he613;
5785: douta=16'hde12;
5786: douta=16'hcd2f;
5787: douta=16'ha46f;
5788: douta=16'h838f;
5789: douta=16'h6b2c;
5790: douta=16'h5a6b;
5791: douta=16'h3145;
5792: douta=16'hac4a;
5793: douta=16'hc4cc;
5794: douta=16'he654;
5795: douta=16'hde33;
5796: douta=16'he654;
5797: douta=16'heeb6;
5798: douta=16'he654;
5799: douta=16'hd572;
5800: douta=16'hc510;
5801: douta=16'hac50;
5802: douta=16'h9430;
5803: douta=16'h8c31;
5804: douta=16'h8432;
5805: douta=16'h8412;
5806: douta=16'h7bf2;
5807: douta=16'h736f;
5808: douta=16'h52ac;
5809: douta=16'h6a8a;
5810: douta=16'hde13;
5811: douta=16'h4ace;
5812: douta=16'h632e;
5813: douta=16'h2147;
5814: douta=16'h10c5;
5815: douta=16'h5b0e;
5816: douta=16'h1083;
5817: douta=16'h10e5;
5818: douta=16'h18e5;
5819: douta=16'h18c4;
5820: douta=16'h18e5;
5821: douta=16'h0883;
5822: douta=16'h73f2;
5823: douta=16'h9492;
5824: douta=16'hacf2;
5825: douta=16'h634d;
5826: douta=16'h42ae;
5827: douta=16'h8d18;
5828: douta=16'h7cb7;
5829: douta=16'h9579;
5830: douta=16'h8d38;
5831: douta=16'h9579;
5832: douta=16'h84f7;
5833: douta=16'h8d18;
5834: douta=16'h7cb6;
5835: douta=16'h84d7;
5836: douta=16'h84f8;
5837: douta=16'h7c96;
5838: douta=16'h84d8;
5839: douta=16'h5352;
5840: douta=16'h8d39;
5841: douta=16'h9dbb;
5842: douta=16'h7496;
5843: douta=16'h8518;
5844: douta=16'h8d5a;
5845: douta=16'h8539;
5846: douta=16'h8539;
5847: douta=16'h7cf8;
5848: douta=16'h84d8;
5849: douta=16'h8518;
5850: douta=16'h7b2a;
5851: douta=16'h18a2;
5852: douta=16'h8d7a;
5853: douta=16'h8538;
5854: douta=16'h95ba;
5855: douta=16'h8518;
5856: douta=16'h8d5a;
5857: douta=16'h9ddb;
5858: douta=16'h8539;
5859: douta=16'h95ba;
5860: douta=16'hae1c;
5861: douta=16'h8d9a;
5862: douta=16'h8d59;
5863: douta=16'ha5db;
5864: douta=16'h9dda;
5865: douta=16'h957a;
5866: douta=16'h8d5a;
5867: douta=16'h7cd9;
5868: douta=16'h8d3a;
5869: douta=16'h7497;
5870: douta=16'h7cb8;
5871: douta=16'h957b;
5872: douta=16'h8d5a;
5873: douta=16'h84f9;
5874: douta=16'h4964;
5875: douta=16'h10a2;
5876: douta=16'h5bb4;
5877: douta=16'h4060;
5878: douta=16'h4b73;
5879: douta=16'h84f9;
5880: douta=16'ha61c;
5881: douta=16'h42f1;
5882: douta=16'h6288;
5883: douta=16'h8d7a;
5884: douta=16'h955a;
5885: douta=16'h8497;
5886: douta=16'h74b8;
5887: douta=16'h0020;
5888: douta=16'h3966;
5889: douta=16'h20c3;
5890: douta=16'h32d2;
5891: douta=16'h3290;
5892: douta=16'h5bf6;
5893: douta=16'h4b32;
5894: douta=16'h3a8f;
5895: douta=16'h7414;
5896: douta=16'h8cf7;
5897: douta=16'ha578;
5898: douta=16'hde34;
5899: douta=16'hee96;
5900: douta=16'hddf3;
5901: douta=16'hd591;
5902: douta=16'hac6c;
5903: douta=16'hb48d;
5904: douta=16'hb4ad;
5905: douta=16'hc530;
5906: douta=16'he654;
5907: douta=16'he675;
5908: douta=16'he634;
5909: douta=16'heeb7;
5910: douta=16'hd571;
5911: douta=16'hee95;
5912: douta=16'hd5b1;
5913: douta=16'hcd50;
5914: douta=16'ha46f;
5915: douta=16'h7b6f;
5916: douta=16'h730e;
5917: douta=16'h62ab;
5918: douta=16'h51c4;
5919: douta=16'hac0b;
5920: douta=16'hc50d;
5921: douta=16'he634;
5922: douta=16'he654;
5923: douta=16'hee95;
5924: douta=16'he655;
5925: douta=16'he654;
5926: douta=16'hddd2;
5927: douta=16'hbcd1;
5928: douta=16'hacb2;
5929: douta=16'h9c71;
5930: douta=16'h9472;
5931: douta=16'h8412;
5932: douta=16'h7bd1;
5933: douta=16'h734e;
5934: douta=16'h62ed;
5935: douta=16'h49e8;
5936: douta=16'hb42b;
5937: douta=16'he633;
5938: douta=16'hcd71;
5939: douta=16'h6b70;
5940: douta=16'h83d0;
5941: douta=16'h31eb;
5942: douta=16'h39ea;
5943: douta=16'h18e5;
5944: douta=16'h1927;
5945: douta=16'h10e6;
5946: douta=16'h18e5;
5947: douta=16'h1905;
5948: douta=16'h1905;
5949: douta=16'h10e4;
5950: douta=16'h08a4;
5951: douta=16'h6bb1;
5952: douta=16'h6c33;
5953: douta=16'h8c30;
5954: douta=16'ha512;
5955: douta=16'h2967;
5956: douta=16'h9dfc;
5957: douta=16'h8d18;
5958: douta=16'h9559;
5959: douta=16'h84f8;
5960: douta=16'h8d38;
5961: douta=16'h9538;
5962: douta=16'h84d7;
5963: douta=16'h7cb7;
5964: douta=16'h8d39;
5965: douta=16'h8d59;
5966: douta=16'h84f8;
5967: douta=16'h84f8;
5968: douta=16'h8cd8;
5969: douta=16'h6c15;
5970: douta=16'h7c96;
5971: douta=16'h8d19;
5972: douta=16'h7cd7;
5973: douta=16'h7cf8;
5974: douta=16'h8d7a;
5975: douta=16'h8539;
5976: douta=16'h8d3a;
5977: douta=16'h8d5a;
5978: douta=16'h6246;
5979: douta=16'h0820;
5980: douta=16'h8519;
5981: douta=16'h9559;
5982: douta=16'h955a;
5983: douta=16'h8d59;
5984: douta=16'h957a;
5985: douta=16'h84d8;
5986: douta=16'h8d39;
5987: douta=16'h84f9;
5988: douta=16'h9dbb;
5989: douta=16'h8d7a;
5990: douta=16'h8d7a;
5991: douta=16'h9dbb;
5992: douta=16'h8d7a;
5993: douta=16'h8d7a;
5994: douta=16'h9dba;
5995: douta=16'h9ddb;
5996: douta=16'h84f9;
5997: douta=16'h959a;
5998: douta=16'h959b;
5999: douta=16'ha61d;
6000: douta=16'h5aad;
6001: douta=16'h8ddf;
6002: douta=16'h7ac8;
6003: douta=16'h3123;
6004: douta=16'h0000;
6005: douta=16'h4374;
6006: douta=16'h2840;
6007: douta=16'h5392;
6008: douta=16'h959a;
6009: douta=16'h7498;
6010: douta=16'h18a2;
6011: douta=16'ha5db;
6012: douta=16'h9d9b;
6013: douta=16'h6c77;
6014: douta=16'h84f8;
6015: douta=16'h0000;
6016: douta=16'h3966;
6017: douta=16'h3146;
6018: douta=16'h3af1;
6019: douta=16'h32b0;
6020: douta=16'h5394;
6021: douta=16'h3aaf;
6022: douta=16'h6c56;
6023: douta=16'h42af;
6024: douta=16'h7414;
6025: douta=16'ha557;
6026: douta=16'hd593;
6027: douta=16'hee75;
6028: douta=16'hd5d2;
6029: douta=16'hc50e;
6030: douta=16'hac6c;
6031: douta=16'hbd0f;
6032: douta=16'hd5d2;
6033: douta=16'he634;
6034: douta=16'hee96;
6035: douta=16'heeb7;
6036: douta=16'hf6d8;
6037: douta=16'hee75;
6038: douta=16'he634;
6039: douta=16'hac2d;
6040: douta=16'hc550;
6041: douta=16'hac70;
6042: douta=16'h8bf0;
6043: douta=16'h6b4d;
6044: douta=16'h628b;
6045: douta=16'h6206;
6046: douta=16'hac2b;
6047: douta=16'hcd2e;
6048: douta=16'he634;
6049: douta=16'he654;
6050: douta=16'hee95;
6051: douta=16'hde13;
6052: douta=16'hd5b2;
6053: douta=16'hcd52;
6054: douta=16'hbd12;
6055: douta=16'hb4f2;
6056: douta=16'h9cb3;
6057: douta=16'h9473;
6058: douta=16'h8433;
6059: douta=16'h736f;
6060: douta=16'h630e;
6061: douta=16'h6b0e;
6062: douta=16'h6227;
6063: douta=16'hc46c;
6064: douta=16'hd590;
6065: douta=16'hde12;
6066: douta=16'hddf2;
6067: douta=16'h8c10;
6068: douta=16'h9432;
6069: douta=16'h5b91;
6070: douta=16'h4aae;
6071: douta=16'h324d;
6072: douta=16'h29c9;
6073: douta=16'h08a4;
6074: douta=16'h428d;
6075: douta=16'h18e5;
6076: douta=16'h10e4;
6077: douta=16'h10e4;
6078: douta=16'h1905;
6079: douta=16'h1906;
6080: douta=16'h0000;
6081: douta=16'h31ea;
6082: douta=16'h0885;
6083: douta=16'h4a6a;
6084: douta=16'h4209;
6085: douta=16'h2169;
6086: douta=16'h959a;
6087: douta=16'h8d18;
6088: douta=16'h8d18;
6089: douta=16'h7c96;
6090: douta=16'h84d7;
6091: douta=16'h84d7;
6092: douta=16'h9579;
6093: douta=16'h7c76;
6094: douta=16'h84d7;
6095: douta=16'h8d18;
6096: douta=16'h8d59;
6097: douta=16'h8d39;
6098: douta=16'h8d39;
6099: douta=16'h7cb7;
6100: douta=16'h8d39;
6101: douta=16'h63b2;
6102: douta=16'h7cb7;
6103: douta=16'h8d7a;
6104: douta=16'h8539;
6105: douta=16'h8519;
6106: douta=16'h8d5b;
6107: douta=16'h95bc;
6108: douta=16'h959a;
6109: douta=16'h74b8;
6110: douta=16'h8519;
6111: douta=16'h957a;
6112: douta=16'h957a;
6113: douta=16'h8d19;
6114: douta=16'h9dbb;
6115: douta=16'h957a;
6116: douta=16'h8d7a;
6117: douta=16'ha5db;
6118: douta=16'ha5db;
6119: douta=16'ha5db;
6120: douta=16'ha5db;
6121: douta=16'h959a;
6122: douta=16'ha5fb;
6123: douta=16'h959a;
6124: douta=16'h959a;
6125: douta=16'ha5dc;
6126: douta=16'h8c95;
6127: douta=16'h5c38;
6128: douta=16'h857c;
6129: douta=16'h5373;
6130: douta=16'h630c;
6131: douta=16'h6245;
6132: douta=16'h0842;
6133: douta=16'h5331;
6134: douta=16'h6458;
6135: douta=16'h10a5;
6136: douta=16'h7cd7;
6137: douta=16'h7c32;
6138: douta=16'h7498;
6139: douta=16'h5352;
6140: douta=16'h6415;
6141: douta=16'h84d8;
6142: douta=16'h0000;
6143: douta=16'h4acd;
6144: douta=16'h3966;
6145: douta=16'h2925;
6146: douta=16'h3a6e;
6147: douta=16'h42f1;
6148: douta=16'h32b0;
6149: douta=16'h6436;
6150: douta=16'h7456;
6151: douta=16'h5b93;
6152: douta=16'h8cb6;
6153: douta=16'h9d16;
6154: douta=16'h6bb1;
6155: douta=16'he653;
6156: douta=16'hac8f;
6157: douta=16'h9389;
6158: douta=16'hcd50;
6159: douta=16'hcd90;
6160: douta=16'he634;
6161: douta=16'heeb7;
6162: douta=16'he675;
6163: douta=16'heeb7;
6164: douta=16'he675;
6165: douta=16'hddf3;
6166: douta=16'hd5d2;
6167: douta=16'hd591;
6168: douta=16'ha450;
6169: douta=16'h8c10;
6170: douta=16'h736e;
6171: douta=16'h6b0c;
6172: douta=16'h3966;
6173: douta=16'hb48c;
6174: douta=16'hd5b0;
6175: douta=16'he634;
6176: douta=16'hee76;
6177: douta=16'he634;
6178: douta=16'hde13;
6179: douta=16'hd5d1;
6180: douta=16'hcd71;
6181: douta=16'hacb1;
6182: douta=16'hc552;
6183: douta=16'h9473;
6184: douta=16'h9c93;
6185: douta=16'h8432;
6186: douta=16'h7390;
6187: douta=16'h6b0e;
6188: douta=16'h6b2e;
6189: douta=16'h8b48;
6190: douta=16'hc4eb;
6191: douta=16'hddf2;
6192: douta=16'he654;
6193: douta=16'he674;
6194: douta=16'hd571;
6195: douta=16'h9c51;
6196: douta=16'h83f1;
6197: douta=16'h8c54;
6198: douta=16'h5b51;
6199: douta=16'h3a8d;
6200: douta=16'h322b;
6201: douta=16'h2168;
6202: douta=16'h10c3;
6203: douta=16'h5330;
6204: douta=16'h18e5;
6205: douta=16'h1905;
6206: douta=16'h10e4;
6207: douta=16'h10c4;
6208: douta=16'h10c5;
6209: douta=16'h0021;
6210: douta=16'h2146;
6211: douta=16'h1105;
6212: douta=16'h3188;
6213: douta=16'h3a28;
6214: douta=16'h31c8;
6215: douta=16'h7435;
6216: douta=16'h84d7;
6217: douta=16'ha5da;
6218: douta=16'h9559;
6219: douta=16'h8d59;
6220: douta=16'h8d18;
6221: douta=16'h8cd8;
6222: douta=16'h6c14;
6223: douta=16'h84f8;
6224: douta=16'h84d7;
6225: douta=16'h63d4;
6226: douta=16'h9d9a;
6227: douta=16'h8d59;
6228: douta=16'h8d39;
6229: douta=16'h84f7;
6230: douta=16'h7c56;
6231: douta=16'h8d59;
6232: douta=16'h8d39;
6233: douta=16'h7c77;
6234: douta=16'h8519;
6235: douta=16'h8539;
6236: douta=16'h8d39;
6237: douta=16'h8539;
6238: douta=16'h7cd8;
6239: douta=16'h8d5a;
6240: douta=16'h8d59;
6241: douta=16'h84f8;
6242: douta=16'h8d3a;
6243: douta=16'h84f8;
6244: douta=16'h8518;
6245: douta=16'h957a;
6246: douta=16'h8d5a;
6247: douta=16'h959a;
6248: douta=16'h8539;
6249: douta=16'h9d9a;
6250: douta=16'ha5db;
6251: douta=16'h95dc;
6252: douta=16'h6b70;
6253: douta=16'h4b32;
6254: douta=16'h4bf7;
6255: douta=16'h4bb5;
6256: douta=16'h53b5;
6257: douta=16'h6cba;
6258: douta=16'h7d5c;
6259: douta=16'h8328;
6260: douta=16'h20c2;
6261: douta=16'h0820;
6262: douta=16'h74d9;
6263: douta=16'h7d5b;
6264: douta=16'h2a8e;
6265: douta=16'h2000;
6266: douta=16'h955a;
6267: douta=16'h7455;
6268: douta=16'h957a;
6269: douta=16'h6bf3;
6270: douta=16'hbdb5;
6271: douta=16'hdeba;
6272: douta=16'h3966;
6273: douta=16'h3145;
6274: douta=16'h31a8;
6275: douta=16'h4333;
6276: douta=16'h3ad1;
6277: douta=16'h5bb4;
6278: douta=16'h7c98;
6279: douta=16'h6c35;
6280: douta=16'h6bd3;
6281: douta=16'h8433;
6282: douta=16'h94d5;
6283: douta=16'hb5b8;
6284: douta=16'ha40b;
6285: douta=16'hc530;
6286: douta=16'hd5f3;
6287: douta=16'hde15;
6288: douta=16'heeb6;
6289: douta=16'heeb6;
6290: douta=16'heeb6;
6291: douta=16'hd591;
6292: douta=16'he675;
6293: douta=16'hd5b2;
6294: douta=16'hbcf1;
6295: douta=16'h9450;
6296: douta=16'h8c10;
6297: douta=16'h838e;
6298: douta=16'h736d;
6299: douta=16'h3945;
6300: douta=16'hbccc;
6301: douta=16'hd570;
6302: douta=16'hee54;
6303: douta=16'hee74;
6304: douta=16'hddf2;
6305: douta=16'hf6b6;
6306: douta=16'hd5b2;
6307: douta=16'hcd71;
6308: douta=16'hb4d1;
6309: douta=16'ha491;
6310: douta=16'h9453;
6311: douta=16'ha4b4;
6312: douta=16'h7bf1;
6313: douta=16'h7bd1;
6314: douta=16'h6b2e;
6315: douta=16'h4a4a;
6316: douta=16'h9329;
6317: douta=16'hc4cc;
6318: douta=16'he632;
6319: douta=16'he654;
6320: douta=16'he633;
6321: douta=16'hddd3;
6322: douta=16'hc4f0;
6323: douta=16'ha491;
6324: douta=16'h9432;
6325: douta=16'h7c13;
6326: douta=16'h8454;
6327: douta=16'h5bb2;
6328: douta=16'h4aef;
6329: douta=16'h3a6d;
6330: douta=16'h3a4e;
6331: douta=16'h3aae;
6332: douta=16'h322b;
6333: douta=16'h10e5;
6334: douta=16'h10c4;
6335: douta=16'h10c4;
6336: douta=16'h18c4;
6337: douta=16'h18e5;
6338: douta=16'h2126;
6339: douta=16'h0883;
6340: douta=16'h424a;
6341: douta=16'h7412;
6342: douta=16'h3166;
6343: douta=16'h52cb;
6344: douta=16'h6b4d;
6345: douta=16'h6391;
6346: douta=16'h8d39;
6347: douta=16'h8497;
6348: douta=16'h8d39;
6349: douta=16'h8d18;
6350: douta=16'h9dba;
6351: douta=16'h8cf7;
6352: douta=16'h84b6;
6353: douta=16'h84b7;
6354: douta=16'h959a;
6355: douta=16'h84d7;
6356: douta=16'h84d7;
6357: douta=16'h8d39;
6358: douta=16'h8d39;
6359: douta=16'ha5db;
6360: douta=16'h6c55;
6361: douta=16'h7c96;
6362: douta=16'h957a;
6363: douta=16'h7476;
6364: douta=16'h7cd8;
6365: douta=16'h8519;
6366: douta=16'h7cd8;
6367: douta=16'h8d5a;
6368: douta=16'h8539;
6369: douta=16'h8519;
6370: douta=16'h7cb8;
6371: douta=16'h959b;
6372: douta=16'h8d5a;
6373: douta=16'h74b8;
6374: douta=16'h8d3a;
6375: douta=16'h959b;
6376: douta=16'h9ddb;
6377: douta=16'h8d9c;
6378: douta=16'h428d;
6379: douta=16'h3b12;
6380: douta=16'h6456;
6381: douta=16'h74b9;
6382: douta=16'h6cda;
6383: douta=16'h3b13;
6384: douta=16'h4353;
6385: douta=16'h4395;
6386: douta=16'h4bf6;
6387: douta=16'h732c;
6388: douta=16'h4144;
6389: douta=16'h0882;
6390: douta=16'h29ca;
6391: douta=16'h6436;
6392: douta=16'h6cd9;
6393: douta=16'h5c57;
6394: douta=16'h5bf6;
6395: douta=16'h63b1;
6396: douta=16'ha535;
6397: douta=16'hadd7;
6398: douta=16'h4aaa;
6399: douta=16'h1840;
6400: douta=16'h3986;
6401: douta=16'h3145;
6402: douta=16'h20e4;
6403: douta=16'h3af1;
6404: douta=16'h4353;
6405: douta=16'h5394;
6406: douta=16'h6c14;
6407: douta=16'h8d18;
6408: douta=16'h8454;
6409: douta=16'h94b5;
6410: douta=16'h94b4;
6411: douta=16'hc619;
6412: douta=16'hcd92;
6413: douta=16'hd613;
6414: douta=16'hde55;
6415: douta=16'heeb7;
6416: douta=16'heeb7;
6417: douta=16'heeb6;
6418: douta=16'hee96;
6419: douta=16'hde35;
6420: douta=16'hbcf0;
6421: douta=16'hcd91;
6422: douta=16'h8c31;
6423: douta=16'h7b90;
6424: douta=16'h83b0;
6425: douta=16'h7b6e;
6426: douta=16'h5207;
6427: douta=16'hb4cd;
6428: douta=16'hd570;
6429: douta=16'he654;
6430: douta=16'he654;
6431: douta=16'he654;
6432: douta=16'he634;
6433: douta=16'hddd2;
6434: douta=16'hcd72;
6435: douta=16'hacb2;
6436: douta=16'hb512;
6437: douta=16'h9473;
6438: douta=16'h9452;
6439: douta=16'h6b6f;
6440: douta=16'h7bd1;
6441: douta=16'h73b0;
6442: douta=16'h5a27;
6443: douta=16'ha3e9;
6444: douta=16'hddb1;
6445: douta=16'he654;
6446: douta=16'hde12;
6447: douta=16'hee54;
6448: douta=16'he633;
6449: douta=16'hd5b1;
6450: douta=16'hc510;
6451: douta=16'ha470;
6452: douta=16'h9432;
6453: douta=16'h8c74;
6454: douta=16'h7c13;
6455: douta=16'h73f3;
6456: douta=16'h6392;
6457: douta=16'h530f;
6458: douta=16'h4acf;
6459: douta=16'h3a6d;
6460: douta=16'h5330;
6461: douta=16'h3a2c;
6462: douta=16'h1926;
6463: douta=16'h1906;
6464: douta=16'h10e5;
6465: douta=16'h2146;
6466: douta=16'h1906;
6467: douta=16'h10e4;
6468: douta=16'h1083;
6469: douta=16'h0041;
6470: douta=16'h5b52;
6471: douta=16'h0001;
6472: douta=16'h29a8;
6473: douta=16'h7b8d;
6474: douta=16'h8c4f;
6475: douta=16'h7b6d;
6476: douta=16'h324d;
6477: douta=16'h8d18;
6478: douta=16'h9d9a;
6479: douta=16'h8d38;
6480: douta=16'h8d38;
6481: douta=16'h8d18;
6482: douta=16'h8d39;
6483: douta=16'h8d18;
6484: douta=16'h8d58;
6485: douta=16'h84d7;
6486: douta=16'h84d7;
6487: douta=16'h8d19;
6488: douta=16'h8d18;
6489: douta=16'h8d39;
6490: douta=16'h8d39;
6491: douta=16'h8d18;
6492: douta=16'h5392;
6493: douta=16'h7476;
6494: douta=16'h7456;
6495: douta=16'h8d39;
6496: douta=16'h8519;
6497: douta=16'h8519;
6498: douta=16'h8519;
6499: douta=16'h8539;
6500: douta=16'h7cf9;
6501: douta=16'h857b;
6502: douta=16'h8d39;
6503: douta=16'h528c;
6504: douta=16'h732d;
6505: douta=16'h1230;
6506: douta=16'h5459;
6507: douta=16'h3b53;
6508: douta=16'h4bd6;
6509: douta=16'h53d6;
6510: douta=16'h5416;
6511: douta=16'h5c37;
6512: douta=16'h53d6;
6513: douta=16'h4bb5;
6514: douta=16'h5416;
6515: douta=16'h5c9a;
6516: douta=16'h72c6;
6517: douta=16'h20e3;
6518: douta=16'h0861;
6519: douta=16'h7d7d;
6520: douta=16'h6436;
6521: douta=16'h8c0e;
6522: douta=16'hce15;
6523: douta=16'hb5d5;
6524: douta=16'h39c6;
6525: douta=16'h28c2;
6526: douta=16'h3944;
6527: douta=16'h3964;
6528: douta=16'h3124;
6529: douta=16'h3965;
6530: douta=16'h1882;
6531: douta=16'h2a4e;
6532: douta=16'h4b95;
6533: douta=16'h3ad1;
6534: douta=16'h6c56;
6535: douta=16'h6c15;
6536: douta=16'h73f3;
6537: douta=16'h73f3;
6538: douta=16'h7c12;
6539: douta=16'had77;
6540: douta=16'h9d16;
6541: douta=16'hee95;
6542: douta=16'he696;
6543: douta=16'heed8;
6544: douta=16'heed7;
6545: douta=16'hee96;
6546: douta=16'hee96;
6547: douta=16'hde13;
6548: douta=16'hc551;
6549: douta=16'h8c10;
6550: douta=16'h83f1;
6551: douta=16'h7390;
6552: douta=16'h734f;
6553: douta=16'h4985;
6554: douta=16'hac4c;
6555: douta=16'hd570;
6556: douta=16'he675;
6557: douta=16'he633;
6558: douta=16'hee75;
6559: douta=16'hde13;
6560: douta=16'hd591;
6561: douta=16'hc530;
6562: douta=16'hc531;
6563: douta=16'ha4b2;
6564: douta=16'h9453;
6565: douta=16'h9472;
6566: douta=16'h83f1;
6567: douta=16'h7bb0;
6568: douta=16'h734f;
6569: douta=16'h7a87;
6570: douta=16'ha3ca;
6571: douta=16'hddd1;
6572: douta=16'he654;
6573: douta=16'hee74;
6574: douta=16'hee54;
6575: douta=16'he632;
6576: douta=16'hddb0;
6577: douta=16'hbd0f;
6578: douta=16'ha450;
6579: douta=16'h9451;
6580: douta=16'h9432;
6581: douta=16'h8c94;
6582: douta=16'h8474;
6583: douta=16'h8475;
6584: douta=16'h7413;
6585: douta=16'h63b2;
6586: douta=16'h5b30;
6587: douta=16'h7b2d;
6588: douta=16'h428d;
6589: douta=16'h3a8d;
6590: douta=16'h10c4;
6591: douta=16'h4acf;
6592: douta=16'h0863;
6593: douta=16'h18e5;
6594: douta=16'h10e4;
6595: douta=16'h10c4;
6596: douta=16'h10e5;
6597: douta=16'h1926;
6598: douta=16'h0000;
6599: douta=16'h1905;
6600: douta=16'h2147;
6601: douta=16'h1926;
6602: douta=16'h5aec;
6603: douta=16'had11;
6604: douta=16'ha4b0;
6605: douta=16'h62eb;
6606: douta=16'h7b8c;
6607: douta=16'h4208;
6608: douta=16'h530e;
6609: douta=16'h7476;
6610: douta=16'h8d59;
6611: douta=16'h8d18;
6612: douta=16'h8518;
6613: douta=16'h9559;
6614: douta=16'h84d7;
6615: douta=16'h8d39;
6616: douta=16'h84f8;
6617: douta=16'h6c76;
6618: douta=16'h8518;
6619: douta=16'h8d39;
6620: douta=16'h84f8;
6621: douta=16'h84f8;
6622: douta=16'h957a;
6623: douta=16'h5371;
6624: douta=16'h74b6;
6625: douta=16'h8539;
6626: douta=16'h8d59;
6627: douta=16'h7496;
6628: douta=16'h42cf;
6629: douta=16'h4310;
6630: douta=16'h42d0;
6631: douta=16'h62ed;
6632: douta=16'h72a9;
6633: douta=16'h6248;
6634: douta=16'h3ad0;
6635: douta=16'h4395;
6636: douta=16'h3b95;
6637: douta=16'h3b33;
6638: douta=16'h3b74;
6639: douta=16'h4374;
6640: douta=16'h6cba;
6641: douta=16'h53d6;
6642: douta=16'h4334;
6643: douta=16'h5c37;
6644: douta=16'h8b26;
6645: douta=16'h51c4;
6646: douta=16'h0882;
6647: douta=16'h08e5;
6648: douta=16'hb593;
6649: douta=16'had10;
6650: douta=16'h3964;
6651: douta=16'h3944;
6652: douta=16'h4164;
6653: douta=16'h41a5;
6654: douta=16'h3985;
6655: douta=16'h49c7;
6656: douta=16'h4a8b;
6657: douta=16'h3965;
6658: douta=16'h20e3;
6659: douta=16'h29aa;
6660: douta=16'h4b94;
6661: douta=16'h4354;
6662: douta=16'h7cd9;
6663: douta=16'h5bb3;
6664: douta=16'h6c35;
6665: douta=16'h8cf6;
6666: douta=16'h9d16;
6667: douta=16'hb576;
6668: douta=16'hb5b8;
6669: douta=16'ha4b2;
6670: douta=16'he696;
6671: douta=16'heeb7;
6672: douta=16'heed7;
6673: douta=16'he675;
6674: douta=16'hde55;
6675: douta=16'hcd72;
6676: douta=16'ha491;
6677: douta=16'h8c11;
6678: douta=16'h7bb0;
6679: douta=16'h6b2e;
6680: douta=16'h49a4;
6681: douta=16'hac4c;
6682: douta=16'hcd2f;
6683: douta=16'he675;
6684: douta=16'heeb7;
6685: douta=16'he633;
6686: douta=16'hd590;
6687: douta=16'hcd50;
6688: douta=16'hc511;
6689: douta=16'hb4b1;
6690: douta=16'ha492;
6691: douta=16'h9432;
6692: douta=16'h8c11;
6693: douta=16'h6b4e;
6694: douta=16'h7b6f;
6695: douta=16'h41a7;
6696: douta=16'h9bca;
6697: douta=16'hc4cd;
6698: douta=16'heeb5;
6699: douta=16'hf6d7;
6700: douta=16'hf6b6;
6701: douta=16'hee95;
6702: douta=16'he613;
6703: douta=16'hd570;
6704: douta=16'hc4f1;
6705: douta=16'ha471;
6706: douta=16'h9c52;
6707: douta=16'h9c72;
6708: douta=16'h8c12;
6709: douta=16'h8412;
6710: douta=16'h7bb1;
6711: douta=16'h7bf2;
6712: douta=16'h6b0d;
6713: douta=16'h5a49;
6714: douta=16'hddaf;
6715: douta=16'hd592;
6716: douta=16'h5b50;
6717: douta=16'h6391;
6718: douta=16'h29ea;
6719: douta=16'h2148;
6720: douta=16'h10e5;
6721: douta=16'h320a;
6722: douta=16'h10c5;
6723: douta=16'h18e5;
6724: douta=16'h1905;
6725: douta=16'h18e5;
6726: douta=16'h10c4;
6727: douta=16'h10e5;
6728: douta=16'h0021;
6729: douta=16'h0884;
6730: douta=16'h4229;
6731: douta=16'h4b52;
6732: douta=16'h2988;
6733: douta=16'h83ed;
6734: douta=16'h83cd;
6735: douta=16'h83ef;
6736: douta=16'h9c4f;
6737: douta=16'h39e8;
6738: douta=16'had32;
6739: douta=16'h4a28;
6740: douta=16'h528a;
6741: douta=16'h29a8;
6742: douta=16'h428c;
6743: douta=16'h4a8c;
6744: douta=16'h4aae;
6745: douta=16'h5b2f;
6746: douta=16'h4aad;
6747: douta=16'h52ef;
6748: douta=16'h31ea;
6749: douta=16'h18c5;
6750: douta=16'h7b2b;
6751: douta=16'h82e6;
6752: douta=16'hb42c;
6753: douta=16'h1968;
6754: douta=16'h4aee;
6755: douta=16'h3a8d;
6756: douta=16'h2a0b;
6757: douta=16'h4310;
6758: douta=16'h63f3;
6759: douta=16'h5bd3;
6760: douta=16'h5372;
6761: douta=16'h6269;
6762: douta=16'h5a49;
6763: douta=16'h62aa;
6764: douta=16'h098c;
6765: douta=16'h3b54;
6766: douta=16'h32d1;
6767: douta=16'h32d1;
6768: douta=16'h4373;
6769: douta=16'h3b53;
6770: douta=16'h6498;
6771: douta=16'h7d9c;
6772: douta=16'h5351;
6773: douta=16'h8307;
6774: douta=16'h94d1;
6775: douta=16'hbd71;
6776: douta=16'h30e2;
6777: douta=16'h3964;
6778: douta=16'h41a5;
6779: douta=16'h41a5;
6780: douta=16'h41a6;
6781: douta=16'h4186;
6782: douta=16'h41a7;
6783: douta=16'h41c7;
6784: douta=16'h6c34;
6785: douta=16'h3945;
6786: douta=16'h2104;
6787: douta=16'h4acf;
6788: douta=16'h3b33;
6789: douta=16'h3ad1;
6790: douta=16'h6c56;
6791: douta=16'h5373;
6792: douta=16'h4b32;
6793: douta=16'h4aef;
6794: douta=16'hadb9;
6795: douta=16'h8411;
6796: douta=16'h94f6;
6797: douta=16'hb5b7;
6798: douta=16'he654;
6799: douta=16'hee96;
6800: douta=16'he696;
6801: douta=16'he675;
6802: douta=16'hd5b3;
6803: douta=16'hc531;
6804: douta=16'h9451;
6805: douta=16'h7b70;
6806: douta=16'h732e;
6807: douta=16'h2904;
6808: douta=16'hac2c;
6809: douta=16'hd570;
6810: douta=16'he634;
6811: douta=16'he655;
6812: douta=16'heeb6;
6813: douta=16'hee75;
6814: douta=16'h83ae;
6815: douta=16'ha491;
6816: douta=16'ha471;
6817: douta=16'h9432;
6818: douta=16'h83d1;
6819: douta=16'h7bd1;
6820: douta=16'h83f1;
6821: douta=16'h736f;
6822: douta=16'h41a7;
6823: douta=16'ha40a;
6824: douta=16'hccee;
6825: douta=16'hee75;
6826: douta=16'hf6d7;
6827: douta=16'hf6b6;
6828: douta=16'he633;
6829: douta=16'hddd2;
6830: douta=16'hbcf0;
6831: douta=16'hb4d1;
6832: douta=16'h9c72;
6833: douta=16'h9c72;
6834: douta=16'h9453;
6835: douta=16'h83f1;
6836: douta=16'h7bb0;
6837: douta=16'h7bb0;
6838: douta=16'h734d;
6839: douta=16'h62cd;
6840: douta=16'h8b29;
6841: douta=16'hddb0;
6842: douta=16'hee75;
6843: douta=16'hddb2;
6844: douta=16'h73f3;
6845: douta=16'h6bd2;
6846: douta=16'h5330;
6847: douta=16'h3a8e;
6848: douta=16'h328d;
6849: douta=16'h2168;
6850: douta=16'h31ca;
6851: douta=16'h2168;
6852: douta=16'h10e5;
6853: douta=16'h18e6;
6854: douta=16'h1926;
6855: douta=16'h1084;
6856: douta=16'h1926;
6857: douta=16'h1926;
6858: douta=16'h1927;
6859: douta=16'h0000;
6860: douta=16'h2146;
6861: douta=16'h2126;
6862: douta=16'h1906;
6863: douta=16'h7bef;
6864: douta=16'h10a4;
6865: douta=16'hde77;
6866: douta=16'h4a48;
6867: douta=16'h2986;
6868: douta=16'h736d;
6869: douta=16'ha4d2;
6870: douta=16'h52aa;
6871: douta=16'h52cb;
6872: douta=16'h39e9;
6873: douta=16'h5acb;
6874: douta=16'h4229;
6875: douta=16'h39c7;
6876: douta=16'hacae;
6877: douta=16'h9348;
6878: douta=16'hb44a;
6879: douta=16'h31c9;
6880: douta=16'h428d;
6881: douta=16'h42ae;
6882: douta=16'h52ee;
6883: douta=16'h42ae;
6884: douta=16'h530f;
6885: douta=16'h6370;
6886: douta=16'h6392;
6887: douta=16'h5b91;
6888: douta=16'h42d0;
6889: douta=16'h5b71;
6890: douta=16'h6371;
6891: douta=16'h5a48;
6892: douta=16'h5a08;
6893: douta=16'h4a8d;
6894: douta=16'h19ee;
6895: douta=16'h3334;
6896: douta=16'h222e;
6897: douta=16'h4bd5;
6898: douta=16'h5c16;
6899: douta=16'h3af1;
6900: douta=16'h7cb7;
6901: douta=16'hb573;
6902: douta=16'h1820;
6903: douta=16'h4985;
6904: douta=16'h49a5;
6905: douta=16'h41a6;
6906: douta=16'h4186;
6907: douta=16'h49e7;
6908: douta=16'h49c7;
6909: douta=16'h41c7;
6910: douta=16'h49c7;
6911: douta=16'h41a7;
6912: douta=16'h5b0d;
6913: douta=16'h3144;
6914: douta=16'h2903;
6915: douta=16'h6bf3;
6916: douta=16'h4bd6;
6917: douta=16'h4332;
6918: douta=16'h6416;
6919: douta=16'h5bb4;
6920: douta=16'h5b73;
6921: douta=16'h63b2;
6922: douta=16'h9d37;
6923: douta=16'h8c94;
6924: douta=16'hb5d8;
6925: douta=16'hb5d8;
6926: douta=16'hc639;
6927: douta=16'he654;
6928: douta=16'he675;
6929: douta=16'hde34;
6930: douta=16'hcdb3;
6931: douta=16'h9471;
6932: douta=16'h8bf2;
6933: douta=16'h6b2d;
6934: douta=16'h28e3;
6935: douta=16'hac8d;
6936: douta=16'hcd90;
6937: douta=16'hee75;
6938: douta=16'hee95;
6939: douta=16'hee96;
6940: douta=16'hddd2;
6941: douta=16'he655;
6942: douta=16'hcd71;
6943: douta=16'h8c12;
6944: douta=16'h5b2f;
6945: douta=16'h7bb1;
6946: douta=16'h83d1;
6947: douta=16'h6b6f;
6948: douta=16'h6b4f;
6949: douta=16'h30e1;
6950: douta=16'habeb;
6951: douta=16'hde12;
6952: douta=16'hf6d7;
6953: douta=16'heeb7;
6954: douta=16'hee96;
6955: douta=16'hee75;
6956: douta=16'he634;
6957: douta=16'hd591;
6958: douta=16'h9c92;
6959: douta=16'h9473;
6960: douta=16'h8432;
6961: douta=16'h8412;
6962: douta=16'h8bf1;
6963: douta=16'h83d0;
6964: douta=16'h7b6e;
6965: douta=16'h62cb;
6966: douta=16'h832b;
6967: douta=16'hbc6b;
6968: douta=16'he674;
6969: douta=16'hee75;
6970: douta=16'hde13;
6971: douta=16'hacb1;
6972: douta=16'h8453;
6973: douta=16'h7c54;
6974: douta=16'h6bf3;
6975: douta=16'h5b92;
6976: douta=16'h5351;
6977: douta=16'h3ad0;
6978: douta=16'h2a4d;
6979: douta=16'h1105;
6980: douta=16'h5311;
6981: douta=16'h1927;
6982: douta=16'h21a9;
6983: douta=16'h2168;
6984: douta=16'h1968;
6985: douta=16'h1927;
6986: douta=16'h1948;
6987: douta=16'h1926;
6988: douta=16'h1926;
6989: douta=16'h0863;
6990: douta=16'h0021;
6991: douta=16'h39ca;
6992: douta=16'h63d2;
6993: douta=16'h0000;
6994: douta=16'h1927;
6995: douta=16'h0084;
6996: douta=16'h2124;
6997: douta=16'h738d;
6998: douta=16'h1925;
6999: douta=16'h634c;
7000: douta=16'h3a29;
7001: douta=16'h2146;
7002: douta=16'h39a8;
7003: douta=16'h9348;
7004: douta=16'hbc4c;
7005: douta=16'h31a8;
7006: douta=16'h3a2a;
7007: douta=16'h426c;
7008: douta=16'h6bd1;
7009: douta=16'h322b;
7010: douta=16'h29cb;
7011: douta=16'h4aae;
7012: douta=16'h3a8d;
7013: douta=16'h5330;
7014: douta=16'h42ae;
7015: douta=16'h4af0;
7016: douta=16'h4b10;
7017: douta=16'h326d;
7018: douta=16'h3aaf;
7019: douta=16'h42d0;
7020: douta=16'h526b;
7021: douta=16'h5229;
7022: douta=16'h5a28;
7023: douta=16'h19cd;
7024: douta=16'h32f2;
7025: douta=16'h2a6f;
7026: douta=16'h2a90;
7027: douta=16'h7c97;
7028: douta=16'h2881;
7029: douta=16'h4184;
7030: douta=16'h51e6;
7031: douta=16'h49a7;
7032: douta=16'h5208;
7033: douta=16'h41a6;
7034: douta=16'h49e8;
7035: douta=16'h41a6;
7036: douta=16'h41c7;
7037: douta=16'h3966;
7038: douta=16'h3966;
7039: douta=16'h3987;
7040: douta=16'h3944;
7041: douta=16'h3103;
7042: douta=16'h2924;
7043: douta=16'h31a9;
7044: douta=16'h29a9;
7045: douta=16'h3a2c;
7046: douta=16'h6391;
7047: douta=16'h9cb4;
7048: douta=16'h8c95;
7049: douta=16'hadb9;
7050: douta=16'h9d56;
7051: douta=16'h94d5;
7052: douta=16'hd679;
7053: douta=16'h8431;
7054: douta=16'h7c12;
7055: douta=16'hde79;
7056: douta=16'hde14;
7057: douta=16'hd5f3;
7058: douta=16'hb512;
7059: douta=16'h8c11;
7060: douta=16'h7390;
7061: douta=16'h28e3;
7062: douta=16'hb4ad;
7063: douta=16'hd5b0;
7064: douta=16'he654;
7065: douta=16'hee75;
7066: douta=16'he634;
7067: douta=16'he654;
7068: douta=16'hd5f3;
7069: douta=16'hc550;
7070: douta=16'hb512;
7071: douta=16'h9c92;
7072: douta=16'h8432;
7073: douta=16'h632f;
7074: douta=16'h630e;
7075: douta=16'h4aae;
7076: douta=16'h82a7;
7077: douta=16'he590;
7078: douta=16'hee34;
7079: douta=16'hee96;
7080: douta=16'heeb6;
7081: douta=16'heeb6;
7082: douta=16'he634;
7083: douta=16'hcdb3;
7084: douta=16'hbd12;
7085: douta=16'h9452;
7086: douta=16'h9c73;
7087: douta=16'h8432;
7088: douta=16'h7bb0;
7089: douta=16'h736e;
7090: douta=16'h730d;
7091: douta=16'h732d;
7092: douta=16'h6228;
7093: douta=16'hb44b;
7094: douta=16'ha3ca;
7095: douta=16'hcd0e;
7096: douta=16'hd5d2;
7097: douta=16'hcd92;
7098: douta=16'hc532;
7099: douta=16'ha492;
7100: douta=16'h94b5;
7101: douta=16'h7413;
7102: douta=16'h7433;
7103: douta=16'h7413;
7104: douta=16'h6c14;
7105: douta=16'h5bd4;
7106: douta=16'h3a8e;
7107: douta=16'h29cb;
7108: douta=16'h320c;
7109: douta=16'h08c5;
7110: douta=16'h29ea;
7111: douta=16'h1106;
7112: douta=16'h10e5;
7113: douta=16'h10e5;
7114: douta=16'h10e5;
7115: douta=16'h10e5;
7116: douta=16'h1926;
7117: douta=16'h1927;
7118: douta=16'h1106;
7119: douta=16'h1927;
7120: douta=16'h1084;
7121: douta=16'h0062;
7122: douta=16'h0884;
7123: douta=16'h10e5;
7124: douta=16'h7c75;
7125: douta=16'h6c14;
7126: douta=16'h18e5;
7127: douta=16'h1905;
7128: douta=16'h08a5;
7129: douta=16'hd50d;
7130: douta=16'hbc8c;
7131: douta=16'h4a4a;
7132: douta=16'h8410;
7133: douta=16'h2168;
7134: douta=16'h426b;
7135: douta=16'h4a8c;
7136: douta=16'h3a4b;
7137: douta=16'h320b;
7138: douta=16'h4ace;
7139: douta=16'h4b10;
7140: douta=16'h4ace;
7141: douta=16'h4b0f;
7142: douta=16'h42ae;
7143: douta=16'h530f;
7144: douta=16'h3a6d;
7145: douta=16'h5372;
7146: douta=16'h5b71;
7147: douta=16'h42f0;
7148: douta=16'h63d4;
7149: douta=16'h3a6c;
7150: douta=16'h5a49;
7151: douta=16'h49c7;
7152: douta=16'h3187;
7153: douta=16'h32f2;
7154: douta=16'h3923;
7155: douta=16'h4185;
7156: douta=16'h51c6;
7157: douta=16'h49a6;
7158: douta=16'h5228;
7159: douta=16'h4186;
7160: douta=16'h49c7;
7161: douta=16'h49c7;
7162: douta=16'h41a7;
7163: douta=16'h39a6;
7164: douta=16'h49e8;
7165: douta=16'h49e8;
7166: douta=16'h4a08;
7167: douta=16'h49e7;
7168: douta=16'h3944;
7169: douta=16'h3965;
7170: douta=16'h3125;
7171: douta=16'h20e5;
7172: douta=16'h29ca;
7173: douta=16'h2189;
7174: douta=16'h29a9;
7175: douta=16'hb490;
7176: douta=16'hac2e;
7177: douta=16'h9bed;
7178: douta=16'hc4af;
7179: douta=16'h630d;
7180: douta=16'h7bd0;
7181: douta=16'h6baf;
7182: douta=16'h6b8f;
7183: douta=16'h634e;
7184: douta=16'h8c52;
7185: douta=16'h9450;
7186: douta=16'hacb1;
7187: douta=16'h736f;
7188: douta=16'h7288;
7189: douta=16'hc52f;
7190: douta=16'hddd2;
7191: douta=16'hee75;
7192: douta=16'hee75;
7193: douta=16'he654;
7194: douta=16'hddd2;
7195: douta=16'hd591;
7196: douta=16'hcd92;
7197: douta=16'ha4b2;
7198: douta=16'h9472;
7199: douta=16'h7bf1;
7200: douta=16'h7bd1;
7201: douta=16'h6b2e;
7202: douta=16'h31a7;
7203: douta=16'h9b88;
7204: douta=16'hd56e;
7205: douta=16'hcdb2;
7206: douta=16'hf6b6;
7207: douta=16'hee75;
7208: douta=16'he654;
7209: douta=16'hcd72;
7210: douta=16'hcd73;
7211: douta=16'hb4f3;
7212: douta=16'ha493;
7213: douta=16'h9452;
7214: douta=16'h7bd0;
7215: douta=16'h8c11;
7216: douta=16'h736d;
7217: douta=16'h732d;
7218: douta=16'h72ea;
7219: douta=16'h932a;
7220: douta=16'hd54e;
7221: douta=16'heeb6;
7222: douta=16'hee75;
7223: douta=16'he674;
7224: douta=16'hddd3;
7225: douta=16'hbd12;
7226: douta=16'ha492;
7227: douta=16'h9432;
7228: douta=16'h8433;
7229: douta=16'h8474;
7230: douta=16'h73f2;
7231: douta=16'h6371;
7232: douta=16'h5331;
7233: douta=16'h5351;
7234: douta=16'h428f;
7235: douta=16'h324d;
7236: douta=16'h42f1;
7237: douta=16'h21ca;
7238: douta=16'h3a2c;
7239: douta=16'h2168;
7240: douta=16'h1084;
7241: douta=16'h320c;
7242: douta=16'h1906;
7243: douta=16'h1926;
7244: douta=16'h2168;
7245: douta=16'h1927;
7246: douta=16'h1927;
7247: douta=16'h1927;
7248: douta=16'h1926;
7249: douta=16'h1906;
7250: douta=16'h1926;
7251: douta=16'h2127;
7252: douta=16'h1905;
7253: douta=16'h0021;
7254: douta=16'h0021;
7255: douta=16'h0021;
7256: douta=16'h10c4;
7257: douta=16'h6bf4;
7258: douta=16'h4b10;
7259: douta=16'h1106;
7260: douta=16'h3a2a;
7261: douta=16'h52ad;
7262: douta=16'h52ac;
7263: douta=16'h5b0e;
7264: douta=16'h6b8f;
7265: douta=16'h3a2c;
7266: douta=16'h42ae;
7267: douta=16'h5b50;
7268: douta=16'h42ce;
7269: douta=16'h42ad;
7270: douta=16'h6bd1;
7271: douta=16'h21ca;
7272: douta=16'h5350;
7273: douta=16'h5b2f;
7274: douta=16'h42ad;
7275: douta=16'h320a;
7276: douta=16'h4a4b;
7277: douta=16'h6ac9;
7278: douta=16'h5207;
7279: douta=16'h2a8f;
7280: douta=16'h4985;
7281: douta=16'h51a5;
7282: douta=16'h5a07;
7283: douta=16'h49c6;
7284: douta=16'h41a6;
7285: douta=16'h4186;
7286: douta=16'h49e8;
7287: douta=16'h49e8;
7288: douta=16'h49e8;
7289: douta=16'h49e7;
7290: douta=16'h41a7;
7291: douta=16'h41c7;
7292: douta=16'h41a7;
7293: douta=16'h41c7;
7294: douta=16'h49c7;
7295: douta=16'h49e7;
7296: douta=16'h4165;
7297: douta=16'h5b2e;
7298: douta=16'h3124;
7299: douta=16'h2904;
7300: douta=16'h2a2b;
7301: douta=16'h29c9;
7302: douta=16'h2188;
7303: douta=16'ha3ed;
7304: douta=16'hac2e;
7305: douta=16'h9bed;
7306: douta=16'hac6e;
7307: douta=16'h52cd;
7308: douta=16'h6b6f;
7309: douta=16'h6baf;
7310: douta=16'h6b8f;
7311: douta=16'h6bb0;
7312: douta=16'h7411;
7313: douta=16'h636f;
7314: douta=16'h530d;
7315: douta=16'hbc8d;
7316: douta=16'hcd6f;
7317: douta=16'hde53;
7318: douta=16'he655;
7319: douta=16'heeb6;
7320: douta=16'he675;
7321: douta=16'he674;
7322: douta=16'hd5b2;
7323: douta=16'hbd11;
7324: douta=16'h9c72;
7325: douta=16'h9c92;
7326: douta=16'h8412;
7327: douta=16'h7b70;
7328: douta=16'h734e;
7329: douta=16'h5a6a;
7330: douta=16'hac2c;
7331: douta=16'he5d0;
7332: douta=16'hf6b6;
7333: douta=16'hf6f7;
7334: douta=16'h62ce;
7335: douta=16'he613;
7336: douta=16'hc552;
7337: douta=16'hacb2;
7338: douta=16'ha4b3;
7339: douta=16'h9452;
7340: douta=16'h9452;
7341: douta=16'h83d0;
7342: douta=16'h734d;
7343: douta=16'h732d;
7344: douta=16'h6b0d;
7345: douta=16'h51a5;
7346: douta=16'hac0a;
7347: douta=16'hd58f;
7348: douta=16'he613;
7349: douta=16'he675;
7350: douta=16'hddd2;
7351: douta=16'hddd2;
7352: douta=16'hc531;
7353: douta=16'hb4d2;
7354: douta=16'h9452;
7355: douta=16'h9452;
7356: douta=16'h7bf2;
7357: douta=16'h6b4f;
7358: douta=16'h6b70;
7359: douta=16'h6b91;
7360: douta=16'h6bb1;
7361: douta=16'h5b10;
7362: douta=16'h52ad;
7363: douta=16'h5aee;
7364: douta=16'hacf3;
7365: douta=16'h3a4d;
7366: douta=16'h6bd3;
7367: douta=16'h3aae;
7368: douta=16'h4b10;
7369: douta=16'h29cb;
7370: douta=16'h0863;
7371: douta=16'h322d;
7372: douta=16'h1947;
7373: douta=16'h1907;
7374: douta=16'h1947;
7375: douta=16'h1927;
7376: douta=16'h1106;
7377: douta=16'h10e5;
7378: douta=16'h1906;
7379: douta=16'h1105;
7380: douta=16'h1926;
7381: douta=16'h10e5;
7382: douta=16'h1905;
7383: douta=16'h1926;
7384: douta=16'h2187;
7385: douta=16'h2988;
7386: douta=16'h10c5;
7387: douta=16'h0000;
7388: douta=16'h0863;
7389: douta=16'h5373;
7390: douta=16'h422a;
7391: douta=16'h6b90;
7392: douta=16'h426b;
7393: douta=16'h5b0e;
7394: douta=16'h632e;
7395: douta=16'h5b70;
7396: douta=16'h5b50;
7397: douta=16'h5b50;
7398: douta=16'h428d;
7399: douta=16'h5330;
7400: douta=16'h530e;
7401: douta=16'h29a8;
7402: douta=16'ha48e;
7403: douta=16'h6268;
7404: douta=16'h6247;
7405: douta=16'h4aaf;
7406: douta=16'h4b94;
7407: douta=16'h6a66;
7408: douta=16'h6a68;
7409: douta=16'h51e6;
7410: douta=16'h5a29;
7411: douta=16'h49c8;
7412: douta=16'h41a7;
7413: douta=16'h49e8;
7414: douta=16'h49c7;
7415: douta=16'h41a7;
7416: douta=16'h41c7;
7417: douta=16'h49c7;
7418: douta=16'h49e7;
7419: douta=16'h49c7;
7420: douta=16'h49e8;
7421: douta=16'h49e8;
7422: douta=16'h41c7;
7423: douta=16'h41c7;
7424: douta=16'h4165;
7425: douta=16'h5b4f;
7426: douta=16'h3145;
7427: douta=16'h3145;
7428: douta=16'h2168;
7429: douta=16'h29a9;
7430: douta=16'h2188;
7431: douta=16'h6aab;
7432: douta=16'hac2e;
7433: douta=16'ha40e;
7434: douta=16'h9c0e;
7435: douta=16'h5aee;
7436: douta=16'h6b8f;
7437: douta=16'h6b6e;
7438: douta=16'h6bd0;
7439: douta=16'h6bb0;
7440: douta=16'h6bb0;
7441: douta=16'h638f;
7442: douta=16'h6baf;
7443: douta=16'h636e;
7444: douta=16'he654;
7445: douta=16'he674;
7446: douta=16'he675;
7447: douta=16'he696;
7448: douta=16'hd5d2;
7449: douta=16'hd5b2;
7450: douta=16'hbd11;
7451: douta=16'h9c71;
7452: douta=16'h9452;
7453: douta=16'h7bd0;
7454: douta=16'h736f;
7455: douta=16'h7b90;
7456: douta=16'h49e6;
7457: douta=16'hb44b;
7458: douta=16'hddf2;
7459: douta=16'heeb7;
7460: douta=16'hee95;
7461: douta=16'he674;
7462: douta=16'hddf4;
7463: douta=16'h8bce;
7464: douta=16'h7b6e;
7465: douta=16'ha493;
7466: douta=16'h9c94;
7467: douta=16'h8c32;
7468: douta=16'h8c11;
7469: douta=16'h7b8e;
7470: douta=16'h7b8f;
7471: douta=16'h49c7;
7472: douta=16'hbc6d;
7473: douta=16'hdd90;
7474: douta=16'hee95;
7475: douta=16'hee96;
7476: douta=16'heeb6;
7477: douta=16'he654;
7478: douta=16'hee74;
7479: douta=16'hddb2;
7480: douta=16'hbd11;
7481: douta=16'h9c93;
7482: douta=16'h83f1;
7483: douta=16'h7bb0;
7484: douta=16'h736f;
7485: douta=16'h630d;
7486: douta=16'h62cd;
7487: douta=16'h736f;
7488: douta=16'h6b70;
7489: douta=16'h62cd;
7490: douta=16'hee53;
7491: douta=16'hb4f1;
7492: douta=16'hacd2;
7493: douta=16'h6392;
7494: douta=16'h6392;
7495: douta=16'h5b72;
7496: douta=16'h42d0;
7497: douta=16'h42ae;
7498: douta=16'h4b10;
7499: douta=16'h2189;
7500: douta=16'h322d;
7501: douta=16'h320c;
7502: douta=16'h1967;
7503: douta=16'h10c5;
7504: douta=16'h10e6;
7505: douta=16'h10e6;
7506: douta=16'h1926;
7507: douta=16'h1105;
7508: douta=16'h18e5;
7509: douta=16'h10e5;
7510: douta=16'h1905;
7511: douta=16'h18e5;
7512: douta=16'h10e5;
7513: douta=16'h1905;
7514: douta=16'h10e4;
7515: douta=16'h1905;
7516: douta=16'h2167;
7517: douta=16'h0000;
7518: douta=16'h3a0a;
7519: douta=16'h1947;
7520: douta=16'h3a2b;
7521: douta=16'h6b90;
7522: douta=16'h632e;
7523: douta=16'h8c31;
7524: douta=16'h4ace;
7525: douta=16'h5b30;
7526: douta=16'h5b0e;
7527: douta=16'h1925;
7528: douta=16'ha513;
7529: douta=16'h93ab;
7530: douta=16'h6a67;
7531: douta=16'h3a6d;
7532: douta=16'h42ce;
7533: douta=16'h6c14;
7534: douta=16'h528d;
7535: douta=16'h6a47;
7536: douta=16'h5a48;
7537: douta=16'h5a29;
7538: douta=16'h5228;
7539: douta=16'h4a08;
7540: douta=16'h49e8;
7541: douta=16'h4a08;
7542: douta=16'h41a7;
7543: douta=16'h3987;
7544: douta=16'h49c7;
7545: douta=16'h49e8;
7546: douta=16'h41a7;
7547: douta=16'h49e8;
7548: douta=16'h5228;
7549: douta=16'h49c7;
7550: douta=16'h41a7;
7551: douta=16'h41a7;
7552: douta=16'h4165;
7553: douta=16'h4a09;
7554: douta=16'h3124;
7555: douta=16'h3124;
7556: douta=16'h29c9;
7557: douta=16'h29a9;
7558: douta=16'h2188;
7559: douta=16'h7b4c;
7560: douta=16'h93cd;
7561: douta=16'hac4e;
7562: douta=16'h9c0e;
7563: douta=16'h5aed;
7564: douta=16'h634e;
7565: douta=16'h636e;
7566: douta=16'h6bd0;
7567: douta=16'h73d0;
7568: douta=16'h638f;
7569: douta=16'h636f;
7570: douta=16'h6baf;
7571: douta=16'h6baf;
7572: douta=16'h5b4e;
7573: douta=16'hf6f6;
7574: douta=16'hee96;
7575: douta=16'hde34;
7576: douta=16'hcd92;
7577: douta=16'hb4d1;
7578: douta=16'ha471;
7579: douta=16'h9431;
7580: douta=16'h7bf1;
7581: douta=16'h6b4f;
7582: douta=16'h736f;
7583: douta=16'h51e5;
7584: douta=16'hbccc;
7585: douta=16'hd591;
7586: douta=16'heeb7;
7587: douta=16'hee95;
7588: douta=16'he675;
7589: douta=16'hd5d3;
7590: douta=16'hc552;
7591: douta=16'h9c93;
7592: douta=16'h9494;
7593: douta=16'h8c54;
7594: douta=16'h6b91;
7595: douta=16'h7bf2;
7596: douta=16'h6b70;
7597: douta=16'h5aef;
7598: douta=16'h6a48;
7599: douta=16'hcd0e;
7600: douta=16'hee95;
7601: douta=16'hd570;
7602: douta=16'he654;
7603: douta=16'hddf3;
7604: douta=16'hddd2;
7605: douta=16'hcd50;
7606: douta=16'hac91;
7607: douta=16'h9411;
7608: douta=16'h8c11;
7609: douta=16'h838f;
7610: douta=16'h734e;
7611: douta=16'h730d;
7612: douta=16'h7b4e;
7613: douta=16'h62cd;
7614: douta=16'h5acb;
7615: douta=16'h734d;
7616: douta=16'he5f2;
7617: douta=16'heeb7;
7618: douta=16'he655;
7619: douta=16'ha4b2;
7620: douta=16'h9cb4;
7621: douta=16'h5b50;
7622: douta=16'h6392;
7623: douta=16'h5b72;
7624: douta=16'h4b10;
7625: douta=16'h4acf;
7626: douta=16'h426d;
7627: douta=16'h42af;
7628: douta=16'h326f;
7629: douta=16'h21aa;
7630: douta=16'h2169;
7631: douta=16'h10a5;
7632: douta=16'h1927;
7633: douta=16'h29ca;
7634: douta=16'h1906;
7635: douta=16'h10e5;
7636: douta=16'h10e5;
7637: douta=16'h18e5;
7638: douta=16'h10e5;
7639: douta=16'h1905;
7640: douta=16'h10c4;
7641: douta=16'h1906;
7642: douta=16'h18e5;
7643: douta=16'h1905;
7644: douta=16'h18e5;
7645: douta=16'h18e5;
7646: douta=16'h1926;
7647: douta=16'h0884;
7648: douta=16'h29ca;
7649: douta=16'h3a8d;
7650: douta=16'h8452;
7651: douta=16'h5b0e;
7652: douta=16'h73d0;
7653: douta=16'h4a4a;
7654: douta=16'hb511;
7655: douta=16'h7aa8;
7656: douta=16'h7aa7;
7657: douta=16'h29a9;
7658: douta=16'h4acf;
7659: douta=16'h5b51;
7660: douta=16'h5b50;
7661: douta=16'h322d;
7662: douta=16'h4a6c;
7663: douta=16'h6a68;
7664: douta=16'h49e8;
7665: douta=16'h5a49;
7666: douta=16'h49e8;
7667: douta=16'h5249;
7668: douta=16'h49c7;
7669: douta=16'h49c7;
7670: douta=16'h41c7;
7671: douta=16'h41a7;
7672: douta=16'h3966;
7673: douta=16'h49e8;
7674: douta=16'h41a7;
7675: douta=16'h49e7;
7676: douta=16'h3986;
7677: douta=16'h41a7;
7678: douta=16'h49c7;
7679: douta=16'h41a7;
7680: douta=16'h28e5;
7681: douta=16'h30e2;
7682: douta=16'h28c2;
7683: douta=16'h3145;
7684: douta=16'h31ea;
7685: douta=16'h2988;
7686: douta=16'h1947;
7687: douta=16'h62ac;
7688: douta=16'h6aec;
7689: douta=16'h730c;
7690: douta=16'h528b;
7691: douta=16'h52cc;
7692: douta=16'h634f;
7693: douta=16'h6bb0;
7694: douta=16'h6b8f;
7695: douta=16'h6bb0;
7696: douta=16'h73f0;
7697: douta=16'h6baf;
7698: douta=16'h6baf;
7699: douta=16'h6bcf;
7700: douta=16'h6baf;
7701: douta=16'h534e;
7702: douta=16'hfeb5;
7703: douta=16'he634;
7704: douta=16'hb511;
7705: douta=16'hacb2;
7706: douta=16'ha492;
7707: douta=16'h83d1;
7708: douta=16'h7370;
7709: douta=16'h7370;
7710: douta=16'h8328;
7711: douta=16'hcd2f;
7712: douta=16'he675;
7713: douta=16'heeb7;
7714: douta=16'heeb7;
7715: douta=16'he675;
7716: douta=16'hd5f3;
7717: douta=16'hb4d2;
7718: douta=16'h8c94;
7719: douta=16'h8c74;
7720: douta=16'h8454;
7721: douta=16'h83f1;
7722: douta=16'h6b4e;
7723: douta=16'h6b0e;
7724: douta=16'h4a6b;
7725: douta=16'h9369;
7726: douta=16'hee74;
7727: douta=16'hf6f7;
7728: douta=16'hd550;
7729: douta=16'hee95;
7730: douta=16'h832b;
7731: douta=16'hbcf0;
7732: douta=16'hac90;
7733: douta=16'h9411;
7734: douta=16'h8bcf;
7735: douta=16'h83d0;
7736: douta=16'h7b6e;
7737: douta=16'h7b6e;
7738: douta=16'h7b2d;
7739: douta=16'h62cc;
7740: douta=16'h730c;
7741: douta=16'he613;
7742: douta=16'he656;
7743: douta=16'heeb7;
7744: douta=16'he656;
7745: douta=16'hd5d5;
7746: douta=16'hb554;
7747: douta=16'h9cd4;
7748: douta=16'h94b4;
7749: douta=16'h6371;
7750: douta=16'h6371;
7751: douta=16'h530f;
7752: douta=16'h4aaf;
7753: douta=16'h4acf;
7754: douta=16'h5b51;
7755: douta=16'h326f;
7756: douta=16'hbd54;
7757: douta=16'h2a2c;
7758: douta=16'h42af;
7759: douta=16'h42af;
7760: douta=16'h21ca;
7761: douta=16'h2168;
7762: douta=16'h10e5;
7763: douta=16'h1906;
7764: douta=16'h21a9;
7765: douta=16'h2147;
7766: douta=16'h10e5;
7767: douta=16'h10e5;
7768: douta=16'h10c5;
7769: douta=16'h10e5;
7770: douta=16'h10c5;
7771: douta=16'h10e5;
7772: douta=16'h10e5;
7773: douta=16'h1905;
7774: douta=16'h10c5;
7775: douta=16'h10c5;
7776: douta=16'h10e5;
7777: douta=16'h0000;
7778: douta=16'h10a4;
7779: douta=16'h2988;
7780: douta=16'had10;
7781: douta=16'h7a67;
7782: douta=16'h8b08;
7783: douta=16'h21cb;
7784: douta=16'h3a2d;
7785: douta=16'h322c;
7786: douta=16'h4b0f;
7787: douta=16'h6bb2;
7788: douta=16'h4b10;
7789: douta=16'h42f0;
7790: douta=16'h3aaf;
7791: douta=16'h6289;
7792: douta=16'h5249;
7793: douta=16'h5208;
7794: douta=16'h5228;
7795: douta=16'h49e8;
7796: douta=16'h49c7;
7797: douta=16'h41a7;
7798: douta=16'h41c7;
7799: douta=16'h49c7;
7800: douta=16'h49e7;
7801: douta=16'h3966;
7802: douta=16'h41a6;
7803: douta=16'h41a7;
7804: douta=16'h41c7;
7805: douta=16'h49c7;
7806: douta=16'h49c7;
7807: douta=16'h41a7;
7808: douta=16'h41a5;
7809: douta=16'h3944;
7810: douta=16'h41c7;
7811: douta=16'h3124;
7812: douta=16'h424b;
7813: douta=16'h29a8;
7814: douta=16'h2989;
7815: douta=16'h4a4a;
7816: douta=16'h5a8b;
7817: douta=16'h5aac;
7818: douta=16'h52cc;
7819: douta=16'h52cd;
7820: douta=16'h5b2e;
7821: douta=16'h636f;
7822: douta=16'h73f1;
7823: douta=16'h6bd0;
7824: douta=16'h6bf1;
7825: douta=16'h6bcf;
7826: douta=16'h638f;
7827: douta=16'h638f;
7828: douta=16'h6bef;
7829: douta=16'h6bd0;
7830: douta=16'h5b6e;
7831: douta=16'hc531;
7832: douta=16'ha490;
7833: douta=16'h8bcf;
7834: douta=16'h9431;
7835: douta=16'h7b6f;
7836: douta=16'h732e;
7837: douta=16'h9b6a;
7838: douta=16'hee76;
7839: douta=16'hee96;
7840: douta=16'hf6d7;
7841: douta=16'heeb7;
7842: douta=16'he675;
7843: douta=16'hd5b3;
7844: douta=16'ha4b3;
7845: douta=16'h9474;
7846: douta=16'h8453;
7847: douta=16'h7bd1;
7848: douta=16'h6b4f;
7849: douta=16'h6b2e;
7850: douta=16'h630d;
7851: douta=16'h49a7;
7852: douta=16'hac2c;
7853: douta=16'hee75;
7854: douta=16'hddf3;
7855: douta=16'hf6d7;
7856: douta=16'h730b;
7857: douta=16'he674;
7858: douta=16'hacd1;
7859: douta=16'ha471;
7860: douta=16'h7bd0;
7861: douta=16'h7baf;
7862: douta=16'h6b2d;
7863: douta=16'h7b6e;
7864: douta=16'h732d;
7865: douta=16'h5249;
7866: douta=16'h39a8;
7867: douta=16'hbc8f;
7868: douta=16'hac6d;
7869: douta=16'hd5d4;
7870: douta=16'hcd94;
7871: douta=16'hcdd5;
7872: douta=16'hc575;
7873: douta=16'hb535;
7874: douta=16'h9cb5;
7875: douta=16'h9494;
7876: douta=16'h9494;
7877: douta=16'h73d1;
7878: douta=16'h6350;
7879: douta=16'h5b30;
7880: douta=16'h4aae;
7881: douta=16'h4ace;
7882: douta=16'h632f;
7883: douta=16'hddd3;
7884: douta=16'h7c74;
7885: douta=16'h5350;
7886: douta=16'h5b72;
7887: douta=16'h4af0;
7888: douta=16'h322c;
7889: douta=16'h29ca;
7890: douta=16'h2189;
7891: douta=16'h1927;
7892: douta=16'h21aa;
7893: douta=16'h42d0;
7894: douta=16'h1968;
7895: douta=16'h2147;
7896: douta=16'h2128;
7897: douta=16'h2169;
7898: douta=16'h29eb;
7899: douta=16'h29aa;
7900: douta=16'h0863;
7901: douta=16'h10e5;
7902: douta=16'h10c5;
7903: douta=16'h10e5;
7904: douta=16'h10c5;
7905: douta=16'h10c4;
7906: douta=16'h2126;
7907: douta=16'h10e5;
7908: douta=16'h10e6;
7909: douta=16'h3a4d;
7910: douta=16'h532f;
7911: douta=16'h428e;
7912: douta=16'h3a4d;
7913: douta=16'h7c13;
7914: douta=16'h5b50;
7915: douta=16'h5330;
7916: douta=16'h42d0;
7917: douta=16'h73f4;
7918: douta=16'h3aaf;
7919: douta=16'had34;
7920: douta=16'h6269;
7921: douta=16'h5249;
7922: douta=16'h49e8;
7923: douta=16'h49c7;
7924: douta=16'h41a7;
7925: douta=16'h49c7;
7926: douta=16'h41a7;
7927: douta=16'h39a6;
7928: douta=16'h41a7;
7929: douta=16'h4186;
7930: douta=16'h39a6;
7931: douta=16'h3986;
7932: douta=16'h41a6;
7933: douta=16'h41a7;
7934: douta=16'h49c8;
7935: douta=16'h49e8;
7936: douta=16'hb468;
7937: douta=16'h4165;
7938: douta=16'h5b2e;
7939: douta=16'h3945;
7940: douta=16'h3167;
7941: douta=16'h29a8;
7942: douta=16'h3a2b;
7943: douta=16'h422a;
7944: douta=16'h4a2b;
7945: douta=16'h4a8c;
7946: douta=16'h426c;
7947: douta=16'h52cd;
7948: douta=16'h5b0e;
7949: douta=16'h638f;
7950: douta=16'h6bb0;
7951: douta=16'h6bb0;
7952: douta=16'h6bd1;
7953: douta=16'h638f;
7954: douta=16'h63af;
7955: douta=16'h6baf;
7956: douta=16'h6bf0;
7957: douta=16'h6bd0;
7958: douta=16'h6baf;
7959: douta=16'h5b4e;
7960: douta=16'h9430;
7961: douta=16'h940f;
7962: douta=16'h7b6e;
7963: douta=16'h6b0e;
7964: douta=16'h3168;
7965: douta=16'hde12;
7966: douta=16'he676;
7967: douta=16'heeb6;
7968: douta=16'hf6f8;
7969: douta=16'he675;
7970: douta=16'hcdb4;
7971: douta=16'hc573;
7972: douta=16'h9494;
7973: douta=16'h8c74;
7974: douta=16'h8413;
7975: douta=16'h6b70;
7976: douta=16'h632e;
7977: douta=16'h6aed;
7978: douta=16'h3945;
7979: douta=16'habe9;
7980: douta=16'hddf2;
7981: douta=16'hee73;
7982: douta=16'he654;
7983: douta=16'hb4af;
7984: douta=16'hb4b1;
7985: douta=16'hac91;
7986: douta=16'h62cc;
7987: douta=16'h8bf0;
7988: douta=16'h83d0;
7989: douta=16'h83f0;
7990: douta=16'h734d;
7991: douta=16'h6aec;
7992: douta=16'h526a;
7993: douta=16'hb44d;
7994: douta=16'he634;
7995: douta=16'hf6f8;
7996: douta=16'he675;
7997: douta=16'hde15;
7998: douta=16'hd5b4;
7999: douta=16'hddf4;
8000: douta=16'hbd34;
8001: douta=16'h8c32;
8002: douta=16'h83f1;
8003: douta=16'h8411;
8004: douta=16'h8412;
8005: douta=16'h7370;
8006: douta=16'h6b4f;
8007: douta=16'h7370;
8008: douta=16'h836f;
8009: douta=16'hddb2;
8010: douta=16'hd5d4;
8011: douta=16'h8c95;
8012: douta=16'h6bb1;
8013: douta=16'h4ace;
8014: douta=16'h52ef;
8015: douta=16'h4ace;
8016: douta=16'h322c;
8017: douta=16'h39eb;
8018: douta=16'h31ca;
8019: douta=16'h1127;
8020: douta=16'h8453;
8021: douta=16'h6bf3;
8022: douta=16'h3a6d;
8023: douta=16'h21eb;
8024: douta=16'h322c;
8025: douta=16'h29eb;
8026: douta=16'h324d;
8027: douta=16'h1969;
8028: douta=16'h1927;
8029: douta=16'h1947;
8030: douta=16'h2168;
8031: douta=16'h10e5;
8032: douta=16'h18e5;
8033: douta=16'h18e6;
8034: douta=16'h10e5;
8035: douta=16'h10c5;
8036: douta=16'h1906;
8037: douta=16'h73f3;
8038: douta=16'h4aef;
8039: douta=16'h5b50;
8040: douta=16'h7413;
8041: douta=16'h5b91;
8042: douta=16'h4aef;
8043: douta=16'h6bd3;
8044: douta=16'h5352;
8045: douta=16'h5352;
8046: douta=16'h4b31;
8047: douta=16'h42ee;
8048: douta=16'h9d78;
8049: douta=16'h6269;
8050: douta=16'h49e8;
8051: douta=16'h49c8;
8052: douta=16'h41a7;
8053: douta=16'h41a7;
8054: douta=16'h41a6;
8055: douta=16'h49c7;
8056: douta=16'h39a6;
8057: douta=16'h4186;
8058: douta=16'h41c7;
8059: douta=16'h3966;
8060: douta=16'h49c8;
8061: douta=16'h49e8;
8062: douta=16'h49e7;
8063: douta=16'h5209;
8064: douta=16'hf5ab;
8065: douta=16'h3965;
8066: douta=16'h630d;
8067: douta=16'h3124;
8068: douta=16'h2924;
8069: douta=16'h2187;
8070: douta=16'h3a2b;
8071: douta=16'h3a0a;
8072: douta=16'h31c9;
8073: douta=16'h422a;
8074: douta=16'h3a4b;
8075: douta=16'h4aac;
8076: douta=16'h52ed;
8077: douta=16'h6390;
8078: douta=16'h6370;
8079: douta=16'h6bd0;
8080: douta=16'h6bb1;
8081: douta=16'h5b2e;
8082: douta=16'h5b6e;
8083: douta=16'h5b6e;
8084: douta=16'h638f;
8085: douta=16'h638e;
8086: douta=16'h530d;
8087: douta=16'h530c;
8088: douta=16'h4acc;
8089: douta=16'h4acb;
8090: douta=16'h632d;
8091: douta=16'h4a8c;
8092: douta=16'hde34;
8093: douta=16'heeb6;
8094: douta=16'heeb6;
8095: douta=16'heed7;
8096: douta=16'hd5b3;
8097: douta=16'hc573;
8098: douta=16'hacd4;
8099: douta=16'had14;
8100: douta=16'h9cb4;
8101: douta=16'h8412;
8102: douta=16'h73b0;
8103: douta=16'h6b2e;
8104: douta=16'h6b2e;
8105: douta=16'h72ca;
8106: douta=16'hc4ee;
8107: douta=16'hddf2;
8108: douta=16'he655;
8109: douta=16'h83d0;
8110: douta=16'hd571;
8111: douta=16'h9c91;
8112: douta=16'h73b0;
8113: douta=16'h83d1;
8114: douta=16'h83d0;
8115: douta=16'h7b8f;
8116: douta=16'h6b0d;
8117: douta=16'h62ed;
8118: douta=16'h31a9;
8119: douta=16'h9bec;
8120: douta=16'he5f3;
8121: douta=16'hf6d7;
8122: douta=16'hd5d2;
8123: douta=16'hde13;
8124: douta=16'hb514;
8125: douta=16'h9453;
8126: douta=16'h9432;
8127: douta=16'h9452;
8128: douta=16'h8c31;
8129: douta=16'h9472;
8130: douta=16'h9492;
8131: douta=16'h8432;
8132: douta=16'h8412;
8133: douta=16'h736e;
8134: douta=16'h9c0f;
8135: douta=16'heeb5;
8136: douta=16'hddf4;
8137: douta=16'hacd4;
8138: douta=16'h9c94;
8139: douta=16'h8433;
8140: douta=16'h6b6f;
8141: douta=16'h630e;
8142: douta=16'h630f;
8143: douta=16'h4a8d;
8144: douta=16'h424c;
8145: douta=16'h29a9;
8146: douta=16'hb491;
8147: douta=16'h7bd2;
8148: douta=16'h5b0f;
8149: douta=16'h5b50;
8150: douta=16'h42ae;
8151: douta=16'h3a4c;
8152: douta=16'h42ae;
8153: douta=16'h21cb;
8154: douta=16'ha4f5;
8155: douta=16'h3a4d;
8156: douta=16'h42cf;
8157: douta=16'h320c;
8158: douta=16'h31eb;
8159: douta=16'h10e5;
8160: douta=16'h4af1;
8161: douta=16'h10c4;
8162: douta=16'h10e5;
8163: douta=16'h10e5;
8164: douta=16'h1906;
8165: douta=16'h0884;
8166: douta=16'h0000;
8167: douta=16'h6bb1;
8168: douta=16'h5b71;
8169: douta=16'h5b72;
8170: douta=16'h8495;
8171: douta=16'h5b72;
8172: douta=16'h5351;
8173: douta=16'h4b31;
8174: douta=16'h63f4;
8175: douta=16'h6c56;
8176: douta=16'h4b73;
8177: douta=16'hadda;
8178: douta=16'h5394;
8179: douta=16'h5227;
8180: douta=16'h49e7;
8181: douta=16'h49c7;
8182: douta=16'h41a6;
8183: douta=16'h41a7;
8184: douta=16'h41a7;
8185: douta=16'h41a7;
8186: douta=16'h49e7;
8187: douta=16'h4a08;
8188: douta=16'h49e8;
8189: douta=16'h49e8;
8190: douta=16'h49e8;
8191: douta=16'h5208;
8192: douta=16'he54a;
8193: douta=16'h28c4;
8194: douta=16'h3945;
8195: douta=16'h3103;
8196: douta=16'h3124;
8197: douta=16'h2147;
8198: douta=16'h1926;
8199: douta=16'h31c9;
8200: douta=16'h31a8;
8201: douta=16'h2987;
8202: douta=16'h3a2a;
8203: douta=16'h4a8c;
8204: douta=16'h4a8c;
8205: douta=16'h530e;
8206: douta=16'h6390;
8207: douta=16'h6bb1;
8208: douta=16'h6bd1;
8209: douta=16'h5b4e;
8210: douta=16'h5b6f;
8211: douta=16'h5b6e;
8212: douta=16'h5b4e;
8213: douta=16'h5b4e;
8214: douta=16'h4acb;
8215: douta=16'h4acc;
8216: douta=16'h532d;
8217: douta=16'h530d;
8218: douta=16'h52ec;
8219: douta=16'h5b2e;
8220: douta=16'h734c;
8221: douta=16'heeb7;
8222: douta=16'he696;
8223: douta=16'he655;
8224: douta=16'hbd12;
8225: douta=16'hc554;
8226: douta=16'hb535;
8227: douta=16'h9cb4;
8228: douta=16'h8412;
8229: douta=16'h738f;
8230: douta=16'h83f2;
8231: douta=16'h6b4e;
8232: douta=16'h9b2a;
8233: douta=16'hddf3;
8234: douta=16'hee96;
8235: douta=16'hee95;
8236: douta=16'he655;
8237: douta=16'ha492;
8238: douta=16'h426d;
8239: douta=16'ha4b3;
8240: douta=16'h7bb0;
8241: douta=16'h734e;
8242: douta=16'h7b8f;
8243: douta=16'h732c;
8244: douta=16'h6acc;
8245: douta=16'h5a8c;
8246: douta=16'hd50e;
8247: douta=16'heed7;
8248: douta=16'heeb7;
8249: douta=16'hb533;
8250: douta=16'hcd93;
8251: douta=16'hb513;
8252: douta=16'h9452;
8253: douta=16'h8432;
8254: douta=16'h52ef;
8255: douta=16'h6b6f;
8256: douta=16'h8c30;
8257: douta=16'h83af;
8258: douta=16'h8c10;
8259: douta=16'h836e;
8260: douta=16'hc552;
8261: douta=16'hd5b3;
8262: douta=16'hacd3;
8263: douta=16'hacd4;
8264: douta=16'had15;
8265: douta=16'h8433;
8266: douta=16'h7bd1;
8267: douta=16'h7bb0;
8268: douta=16'h6b0e;
8269: douta=16'h630e;
8270: douta=16'h630e;
8271: douta=16'h52ad;
8272: douta=16'h9451;
8273: douta=16'hacd3;
8274: douta=16'h8412;
8275: douta=16'h6b6f;
8276: douta=16'h630e;
8277: douta=16'h52cd;
8278: douta=16'h424c;
8279: douta=16'h324c;
8280: douta=16'h52ae;
8281: douta=16'h9453;
8282: douta=16'h7bf3;
8283: douta=16'h530f;
8284: douta=16'h42ae;
8285: douta=16'h426d;
8286: douta=16'h29ca;
8287: douta=16'h2168;
8288: douta=16'h320b;
8289: douta=16'h29ca;
8290: douta=16'h1906;
8291: douta=16'h1906;
8292: douta=16'h10c5;
8293: douta=16'h10a4;
8294: douta=16'h1926;
8295: douta=16'h0083;
8296: douta=16'h84b5;
8297: douta=16'h73f3;
8298: douta=16'h8cd6;
8299: douta=16'h5331;
8300: douta=16'h63f5;
8301: douta=16'h63f4;
8302: douta=16'h4332;
8303: douta=16'h5bf5;
8304: douta=16'h7cb8;
8305: douta=16'h53b4;
8306: douta=16'h8518;
8307: douta=16'h755b;
8308: douta=16'h49e8;
8309: douta=16'h41a7;
8310: douta=16'h41a6;
8311: douta=16'h41a6;
8312: douta=16'h49c7;
8313: douta=16'h49e7;
8314: douta=16'h5228;
8315: douta=16'h5208;
8316: douta=16'h5249;
8317: douta=16'h5208;
8318: douta=16'h5228;
8319: douta=16'h5228;
8320: douta=16'hdd2b;
8321: douta=16'h41c5;
8322: douta=16'h30e3;
8323: douta=16'h3124;
8324: douta=16'h3924;
8325: douta=16'h2168;
8326: douta=16'h1926;
8327: douta=16'h29a9;
8328: douta=16'h2988;
8329: douta=16'h320b;
8330: douta=16'h3a2b;
8331: douta=16'h3a4b;
8332: douta=16'h4aad;
8333: douta=16'h5b2f;
8334: douta=16'h5b4f;
8335: douta=16'h4aed;
8336: douta=16'h5b4f;
8337: douta=16'h532e;
8338: douta=16'h5b4e;
8339: douta=16'h5b4e;
8340: douta=16'h5b6f;
8341: douta=16'h638f;
8342: douta=16'h5b6e;
8343: douta=16'h4acc;
8344: douta=16'h530d;
8345: douta=16'h530d;
8346: douta=16'h4aac;
8347: douta=16'h530c;
8348: douta=16'h532d;
8349: douta=16'hacb1;
8350: douta=16'hd5f5;
8351: douta=16'hd5f4;
8352: douta=16'hbd53;
8353: douta=16'ha4d4;
8354: douta=16'ha4f5;
8355: douta=16'h9cd4;
8356: douta=16'h8411;
8357: douta=16'h734e;
8358: douta=16'h6b2e;
8359: douta=16'he5d1;
8360: douta=16'heeb5;
8361: douta=16'heed7;
8362: douta=16'heeb7;
8363: douta=16'he635;
8364: douta=16'hcd73;
8365: douta=16'h9cb3;
8366: douta=16'h8453;
8367: douta=16'h6bd3;
8368: douta=16'h5acd;
8369: douta=16'h6b0d;
8370: douta=16'h6acc;
8371: douta=16'h5a8b;
8372: douta=16'h72ea;
8373: douta=16'he612;
8374: douta=16'hf6f8;
8375: douta=16'hee96;
8376: douta=16'hcdb4;
8377: douta=16'hb514;
8378: douta=16'h8c94;
8379: douta=16'hacd4;
8380: douta=16'h9452;
8381: douta=16'h8412;
8382: douta=16'h83f1;
8383: douta=16'h7baf;
8384: douta=16'h734e;
8385: douta=16'h93ee;
8386: douta=16'he613;
8387: douta=16'hc553;
8388: douta=16'hc553;
8389: douta=16'h9c53;
8390: douta=16'h9452;
8391: douta=16'ha4d4;
8392: douta=16'h8c53;
8393: douta=16'h8432;
8394: douta=16'h736e;
8395: douta=16'h734e;
8396: douta=16'h6b2e;
8397: douta=16'h62ac;
8398: douta=16'h83d0;
8399: douta=16'ha493;
8400: douta=16'h9c94;
8401: douta=16'h83d1;
8402: douta=16'h734f;
8403: douta=16'h630e;
8404: douta=16'h5b0d;
8405: douta=16'h52ad;
8406: douta=16'h424c;
8407: douta=16'hacd4;
8408: douta=16'h8c73;
8409: douta=16'h8452;
8410: douta=16'h7bf2;
8411: douta=16'h4a8d;
8412: douta=16'h52ce;
8413: douta=16'h3a4d;
8414: douta=16'h320b;
8415: douta=16'h5b72;
8416: douta=16'h6bf3;
8417: douta=16'h530f;
8418: douta=16'h2189;
8419: douta=16'h29aa;
8420: douta=16'h0884;
8421: douta=16'h08c4;
8422: douta=16'h18e5;
8423: douta=16'h10e6;
8424: douta=16'h6371;
8425: douta=16'h6bf3;
8426: douta=16'h6c35;
8427: douta=16'h7435;
8428: douta=16'h7456;
8429: douta=16'h6c56;
8430: douta=16'h5bb4;
8431: douta=16'h7497;
8432: douta=16'h5394;
8433: douta=16'h5bd4;
8434: douta=16'h4b93;
8435: douta=16'h74b8;
8436: douta=16'h8d7a;
8437: douta=16'h959c;
8438: douta=16'h3924;
8439: douta=16'h49e7;
8440: douta=16'h49e8;
8441: douta=16'h5208;
8442: douta=16'h5249;
8443: douta=16'h5208;
8444: douta=16'h5208;
8445: douta=16'h5208;
8446: douta=16'h5228;
8447: douta=16'h5228;
8448: douta=16'hdd4b;
8449: douta=16'hac29;
8450: douta=16'h3945;
8451: douta=16'h630d;
8452: douta=16'h3924;
8453: douta=16'h10e4;
8454: douta=16'h10a4;
8455: douta=16'h2125;
8456: douta=16'h1905;
8457: douta=16'h31eb;
8458: douta=16'h322b;
8459: douta=16'h320b;
8460: douta=16'h3a2b;
8461: douta=16'h4ace;
8462: douta=16'h532f;
8463: douta=16'h532f;
8464: douta=16'h5b4f;
8465: douta=16'h4acd;
8466: douta=16'h4aed;
8467: douta=16'h530d;
8468: douta=16'h4b0d;
8469: douta=16'h534e;
8470: douta=16'h5b6f;
8471: douta=16'h4aac;
8472: douta=16'h532d;
8473: douta=16'h636f;
8474: douta=16'h5b2d;
8475: douta=16'h5b4e;
8476: douta=16'h6bd0;
8477: douta=16'h6bf1;
8478: douta=16'h4b2f;
8479: douta=16'hacd2;
8480: douta=16'hacb2;
8481: douta=16'hacd3;
8482: douta=16'h8c73;
8483: douta=16'h736e;
8484: douta=16'h62cd;
8485: douta=16'h4a2b;
8486: douta=16'hbc6b;
8487: douta=16'hd571;
8488: douta=16'hbd10;
8489: douta=16'heeb7;
8490: douta=16'hddd2;
8491: douta=16'hcdb4;
8492: douta=16'hacf4;
8493: douta=16'h9493;
8494: douta=16'h7bd1;
8495: douta=16'h734e;
8496: douta=16'h6b2e;
8497: douta=16'h422b;
8498: douta=16'h2189;
8499: douta=16'hac0c;
8500: douta=16'he654;
8501: douta=16'hee75;
8502: douta=16'hc533;
8503: douta=16'ha4d4;
8504: douta=16'h8432;
8505: douta=16'h9473;
8506: douta=16'h8433;
8507: douta=16'h8432;
8508: douta=16'h83f0;
8509: douta=16'h83b0;
8510: douta=16'h7b6f;
8511: douta=16'h6b0c;
8512: douta=16'he5d4;
8513: douta=16'hbd12;
8514: douta=16'h9495;
8515: douta=16'ha4b3;
8516: douta=16'h9c74;
8517: douta=16'h8c12;
8518: douta=16'h9452;
8519: douta=16'h83f0;
8520: douta=16'h7b6e;
8521: douta=16'h7b4d;
8522: douta=16'h730c;
8523: douta=16'h732d;
8524: douta=16'hb535;
8525: douta=16'ha4b4;
8526: douta=16'h9453;
8527: douta=16'h8bf1;
8528: douta=16'h83d0;
8529: douta=16'h83d0;
8530: douta=16'h7b6f;
8531: douta=16'h6b2f;
8532: douta=16'h52cc;
8533: douta=16'h73d0;
8534: douta=16'h8412;
8535: douta=16'h83f1;
8536: douta=16'h7bd1;
8537: douta=16'h7390;
8538: douta=16'h6b4f;
8539: douta=16'h52cd;
8540: douta=16'h4aad;
8541: douta=16'h4a8d;
8542: douta=16'h5aee;
8543: douta=16'hc575;
8544: douta=16'h6bb2;
8545: douta=16'h63b2;
8546: douta=16'h4aae;
8547: douta=16'h2189;
8548: douta=16'h1906;
8549: douta=16'h1906;
8550: douta=16'h10e5;
8551: douta=16'h10c5;
8552: douta=16'h10e5;
8553: douta=16'h5312;
8554: douta=16'h5bf3;
8555: douta=16'h8cf7;
8556: douta=16'h63f4;
8557: douta=16'h5393;
8558: douta=16'h8d39;
8559: douta=16'h7cb7;
8560: douta=16'h6c35;
8561: douta=16'h6c37;
8562: douta=16'h6c57;
8563: douta=16'h855b;
8564: douta=16'h21c9;
8565: douta=16'h29ca;
8566: douta=16'h1947;
8567: douta=16'h5a69;
8568: douta=16'h4a28;
8569: douta=16'h5228;
8570: douta=16'h5229;
8571: douta=16'h5228;
8572: douta=16'h5208;
8573: douta=16'h49e8;
8574: douta=16'h4a08;
8575: douta=16'h49c7;
8576: douta=16'hdd4b;
8577: douta=16'hedec;
8578: douta=16'h4165;
8579: douta=16'h7bd1;
8580: douta=16'h4165;
8581: douta=16'h10a3;
8582: douta=16'h1905;
8583: douta=16'h2146;
8584: douta=16'h2105;
8585: douta=16'h29ea;
8586: douta=16'h322b;
8587: douta=16'h29ea;
8588: douta=16'h428d;
8589: douta=16'h4ace;
8590: douta=16'h4ace;
8591: douta=16'h530e;
8592: douta=16'h530e;
8593: douta=16'h3a6b;
8594: douta=16'h4aad;
8595: douta=16'h530e;
8596: douta=16'h530e;
8597: douta=16'h4aed;
8598: douta=16'h4aed;
8599: douta=16'h4acc;
8600: douta=16'h4aac;
8601: douta=16'h4aac;
8602: douta=16'h5b2e;
8603: douta=16'h636f;
8604: douta=16'h5b6f;
8605: douta=16'h63d0;
8606: douta=16'h63d0;
8607: douta=16'h63d0;
8608: douta=16'h536f;
8609: douta=16'h7bd0;
8610: douta=16'h9411;
8611: douta=16'h6b2d;
8612: douta=16'h39c8;
8613: douta=16'hbcae;
8614: douta=16'he614;
8615: douta=16'hf759;
8616: douta=16'hb4f1;
8617: douta=16'he675;
8618: douta=16'hb4d3;
8619: douta=16'h9c93;
8620: douta=16'h83f1;
8621: douta=16'h7bd1;
8622: douta=16'h734e;
8623: douta=16'h6b2d;
8624: douta=16'h62cc;
8625: douta=16'h4a4b;
8626: douta=16'he613;
8627: douta=16'he674;
8628: douta=16'hd5f5;
8629: douta=16'hbd54;
8630: douta=16'ha515;
8631: douta=16'h8c94;
8632: douta=16'h9453;
8633: douta=16'h632f;
8634: douta=16'h5b0e;
8635: douta=16'h838f;
8636: douta=16'h838f;
8637: douta=16'h5a6c;
8638: douta=16'hf6b6;
8639: douta=16'he655;
8640: douta=16'hb514;
8641: douta=16'h8453;
8642: douta=16'h94b5;
8643: douta=16'h6b91;
8644: douta=16'h6371;
8645: douta=16'h9430;
8646: douta=16'h732d;
8647: douta=16'h6aec;
8648: douta=16'h5249;
8649: douta=16'h8c11;
8650: douta=16'h6b70;
8651: douta=16'h8412;
8652: douta=16'h7baf;
8653: douta=16'h736f;
8654: douta=16'h736f;
8655: douta=16'h7b8f;
8656: douta=16'h62ee;
8657: douta=16'h6b4e;
8658: douta=16'ha493;
8659: douta=16'hcdd4;
8660: douta=16'ha4d4;
8661: douta=16'h8c53;
8662: douta=16'h8c53;
8663: douta=16'h8c52;
8664: douta=16'h73b0;
8665: douta=16'h7390;
8666: douta=16'h73b0;
8667: douta=16'h632e;
8668: douta=16'h7b6e;
8669: douta=16'hd5d5;
8670: douta=16'hc554;
8671: douta=16'h9cf5;
8672: douta=16'h8474;
8673: douta=16'h6bb2;
8674: douta=16'h4b10;
8675: douta=16'h3a2c;
8676: douta=16'h3a8d;
8677: douta=16'h2168;
8678: douta=16'h5b31;
8679: douta=16'h2126;
8680: douta=16'h2168;
8681: douta=16'h1905;
8682: douta=16'h5b93;
8683: douta=16'h8cf6;
8684: douta=16'h6c14;
8685: douta=16'h8cf8;
8686: douta=16'h84d8;
8687: douta=16'h7c75;
8688: douta=16'h5bb4;
8689: douta=16'h5bf5;
8690: douta=16'h84f9;
8691: douta=16'h1926;
8692: douta=16'h29ca;
8693: douta=16'h21a9;
8694: douta=16'h31c9;
8695: douta=16'h29c9;
8696: douta=16'h320a;
8697: douta=16'h49c7;
8698: douta=16'h5249;
8699: douta=16'h5229;
8700: douta=16'h5228;
8701: douta=16'h49e8;
8702: douta=16'h49e8;
8703: douta=16'h49e8;
8704: douta=16'he56c;
8705: douta=16'he54b;
8706: douta=16'h3924;
8707: douta=16'h628a;
8708: douta=16'h1861;
8709: douta=16'h52ac;
8710: douta=16'h31c8;
8711: douta=16'h7b0c;
8712: douta=16'h9d16;
8713: douta=16'h29c9;
8714: douta=16'h320b;
8715: douta=16'h29ca;
8716: douta=16'h3a4c;
8717: douta=16'h3a6d;
8718: douta=16'h4aee;
8719: douta=16'h4aee;
8720: douta=16'h4ace;
8721: douta=16'h322a;
8722: douta=16'h3a6b;
8723: douta=16'h428c;
8724: douta=16'h4acd;
8725: douta=16'h4b0e;
8726: douta=16'h4aed;
8727: douta=16'h428b;
8728: douta=16'h4aac;
8729: douta=16'h52ed;
8730: douta=16'h4acc;
8731: douta=16'h530d;
8732: douta=16'h534e;
8733: douta=16'h5b8f;
8734: douta=16'h5b8f;
8735: douta=16'h5b8f;
8736: douta=16'h63b0;
8737: douta=16'h63d0;
8738: douta=16'h5b8f;
8739: douta=16'h634f;
8740: douta=16'hbcd1;
8741: douta=16'hc4f0;
8742: douta=16'hf6b6;
8743: douta=16'hc511;
8744: douta=16'hcd52;
8745: douta=16'hacb2;
8746: douta=16'h9c92;
8747: douta=16'h8c53;
8748: douta=16'h6b2e;
8749: douta=16'h62ec;
8750: douta=16'h62cc;
8751: douta=16'h5a6a;
8752: douta=16'h524a;
8753: douta=16'he635;
8754: douta=16'h7414;
8755: douta=16'hbd75;
8756: douta=16'h94d5;
8757: douta=16'h94d5;
8758: douta=16'h94b5;
8759: douta=16'h8432;
8760: douta=16'h736f;
8761: douta=16'h7b90;
8762: douta=16'h7b6f;
8763: douta=16'h62cd;
8764: douta=16'hd52f;
8765: douta=16'hcd93;
8766: douta=16'ha4d4;
8767: douta=16'h8c33;
8768: douta=16'h8434;
8769: douta=16'h73f1;
8770: douta=16'h4a8d;
8771: douta=16'h7b8f;
8772: douta=16'h6acc;
8773: douta=16'h732e;
8774: douta=16'h5aab;
8775: douta=16'h8bf1;
8776: douta=16'h7bf1;
8777: douta=16'h7b8f;
8778: douta=16'h5aed;
8779: douta=16'h73b0;
8780: douta=16'h7bb0;
8781: douta=16'h734e;
8782: douta=16'h52ac;
8783: douta=16'h9410;
8784: douta=16'hac93;
8785: douta=16'hb4d3;
8786: douta=16'h8c53;
8787: douta=16'h8412;
8788: douta=16'h8412;
8789: douta=16'h7bd1;
8790: douta=16'h7b90;
8791: douta=16'h6b2e;
8792: douta=16'h6b6f;
8793: douta=16'h630e;
8794: douta=16'h9410;
8795: douta=16'he676;
8796: douta=16'he677;
8797: douta=16'hde36;
8798: douta=16'ha515;
8799: douta=16'h8c74;
8800: douta=16'h73f2;
8801: douta=16'h6391;
8802: douta=16'h5b30;
8803: douta=16'h5b30;
8804: douta=16'h324d;
8805: douta=16'h428e;
8806: douta=16'h52ee;
8807: douta=16'h2146;
8808: douta=16'h18e4;
8809: douta=16'h10c4;
8810: douta=16'h2168;
8811: douta=16'h84d7;
8812: douta=16'h8495;
8813: douta=16'h7435;
8814: douta=16'h63f4;
8815: douta=16'h7456;
8816: douta=16'h7476;
8817: douta=16'h9d9a;
8818: douta=16'h29a8;
8819: douta=16'h29a9;
8820: douta=16'h39eb;
8821: douta=16'h3a0b;
8822: douta=16'h3a4c;
8823: douta=16'h3a8d;
8824: douta=16'h4b31;
8825: douta=16'h6477;
8826: douta=16'h51e7;
8827: douta=16'h3987;
8828: douta=16'h3987;
8829: douta=16'h49c7;
8830: douta=16'h4a08;
8831: douta=16'h49e8;
8832: douta=16'he56c;
8833: douta=16'hdd4b;
8834: douta=16'h49c5;
8835: douta=16'h5164;
8836: douta=16'h9432;
8837: douta=16'h83f2;
8838: douta=16'h734f;
8839: douta=16'ha410;
8840: douta=16'had78;
8841: douta=16'h21ca;
8842: douta=16'h322c;
8843: douta=16'h2189;
8844: douta=16'h3a4c;
8845: douta=16'h3a6d;
8846: douta=16'h3a6c;
8847: douta=16'h42ae;
8848: douta=16'h4ace;
8849: douta=16'h324b;
8850: douta=16'h322b;
8851: douta=16'h3a6b;
8852: douta=16'h3a6b;
8853: douta=16'h3a6b;
8854: douta=16'h42cd;
8855: douta=16'h4b0e;
8856: douta=16'h31e9;
8857: douta=16'h4a8c;
8858: douta=16'h424b;
8859: douta=16'h530e;
8860: douta=16'h5b4f;
8861: douta=16'h5b6f;
8862: douta=16'h42ac;
8863: douta=16'h5b6f;
8864: douta=16'h5b8f;
8865: douta=16'h6390;
8866: douta=16'h63d1;
8867: douta=16'h5b70;
8868: douta=16'h4b2e;
8869: douta=16'hc510;
8870: douta=16'hbcf2;
8871: douta=16'hacb2;
8872: douta=16'hc533;
8873: douta=16'h8432;
8874: douta=16'h9473;
8875: douta=16'h83d0;
8876: douta=16'h7b90;
8877: douta=16'h6b0d;
8878: douta=16'h62cc;
8879: douta=16'h8b29;
8880: douta=16'hde55;
8881: douta=16'hde35;
8882: douta=16'h9d16;
8883: douta=16'h8c74;
8884: douta=16'h94b5;
8885: douta=16'h8c94;
8886: douta=16'h8c53;
8887: douta=16'h734e;
8888: douta=16'h734f;
8889: douta=16'h8390;
8890: douta=16'h730d;
8891: douta=16'hd5b3;
8892: douta=16'hbd75;
8893: douta=16'hbd55;
8894: douta=16'had35;
8895: douta=16'h8434;
8896: douta=16'h6bb1;
8897: douta=16'h736f;
8898: douta=16'h39eb;
8899: douta=16'h420a;
8900: douta=16'h31a8;
8901: douta=16'h7bb0;
8902: douta=16'h7bd1;
8903: douta=16'h732e;
8904: douta=16'h5a8b;
8905: douta=16'h732d;
8906: douta=16'h730c;
8907: douta=16'h31c9;
8908: douta=16'h39c9;
8909: douta=16'hcdb4;
8910: douta=16'hb514;
8911: douta=16'h9cb5;
8912: douta=16'h9494;
8913: douta=16'h7bd1;
8914: douta=16'h734e;
8915: douta=16'h6b0e;
8916: douta=16'h62ed;
8917: douta=16'h5aed;
8918: douta=16'h31ca;
8919: douta=16'h62ac;
8920: douta=16'hee75;
8921: douta=16'he697;
8922: douta=16'hcdf7;
8923: douta=16'hc5b6;
8924: douta=16'had15;
8925: douta=16'had15;
8926: douta=16'h8452;
8927: douta=16'h6b91;
8928: douta=16'h6b90;
8929: douta=16'h6b91;
8930: douta=16'h5b30;
8931: douta=16'h4ace;
8932: douta=16'h3a2c;
8933: douta=16'hc574;
8934: douta=16'h21aa;
8935: douta=16'h18c5;
8936: douta=16'h31c9;
8937: douta=16'h10c4;
8938: douta=16'h18e5;
8939: douta=16'h0083;
8940: douta=16'h63b2;
8941: douta=16'h9d58;
8942: douta=16'h84b5;
8943: douta=16'h9d58;
8944: douta=16'h7c76;
8945: douta=16'h5330;
8946: douta=16'h6414;
8947: douta=16'h6c14;
8948: douta=16'h6c77;
8949: douta=16'h6bf3;
8950: douta=16'h630c;
8951: douta=16'h6247;
8952: douta=16'h6a46;
8953: douta=16'h61e4;
8954: douta=16'h59e5;
8955: douta=16'h5a28;
8956: douta=16'h49e8;
8957: douta=16'h41a7;
8958: douta=16'h49c7;
8959: douta=16'h41c7;
8960: douta=16'he58e;
8961: douta=16'he56c;
8962: douta=16'hac48;
8963: douta=16'h6226;
8964: douta=16'hcdb7;
8965: douta=16'h9c53;
8966: douta=16'h83b0;
8967: douta=16'hcd96;
8968: douta=16'hb577;
8969: douta=16'h1906;
8970: douta=16'h08a4;
8971: douta=16'h21a9;
8972: douta=16'h2188;
8973: douta=16'h31eb;
8974: douta=16'h3a6d;
8975: douta=16'h3a6c;
8976: douta=16'h29eb;
8977: douta=16'h3a4b;
8978: douta=16'h3a6c;
8979: douta=16'h322b;
8980: douta=16'h322b;
8981: douta=16'h324b;
8982: douta=16'h428c;
8983: douta=16'h42ac;
8984: douta=16'h4aed;
8985: douta=16'h52ee;
8986: douta=16'h4acd;
8987: douta=16'h42ac;
8988: douta=16'h428c;
8989: douta=16'h532e;
8990: douta=16'h5b6f;
8991: douta=16'h534f;
8992: douta=16'h5b6f;
8993: douta=16'h5b6f;
8994: douta=16'h63b0;
8995: douta=16'h5b8f;
8996: douta=16'h636f;
8997: douta=16'h6bb0;
8998: douta=16'h736f;
8999: douta=16'h9c50;
9000: douta=16'h9430;
9001: douta=16'h7bcf;
9002: douta=16'h7b8f;
9003: douta=16'h7bb0;
9004: douta=16'h732d;
9005: douta=16'h528c;
9006: douta=16'hf694;
9007: douta=16'hee97;
9008: douta=16'he696;
9009: douta=16'had36;
9010: douta=16'h9cf6;
9011: douta=16'h7c13;
9012: douta=16'h9cd4;
9013: douta=16'h7c11;
9014: douta=16'h632f;
9015: douta=16'h630d;
9016: douta=16'h5ace;
9017: douta=16'hbc8f;
9018: douta=16'hddd4;
9019: douta=16'hd5d4;
9020: douta=16'h94b4;
9021: douta=16'h73f2;
9022: douta=16'h52ae;
9023: douta=16'h83ae;
9024: douta=16'h732e;
9025: douta=16'h6b0c;
9026: douta=16'h5a6a;
9027: douta=16'h8bf1;
9028: douta=16'h9473;
9029: douta=16'h632f;
9030: douta=16'h62ac;
9031: douta=16'h6acb;
9032: douta=16'h62cb;
9033: douta=16'h5a8a;
9034: douta=16'h3987;
9035: douta=16'he5f5;
9036: douta=16'h8c55;
9037: douta=16'h9454;
9038: douta=16'h9473;
9039: douta=16'h7bf2;
9040: douta=16'h8433;
9041: douta=16'h736f;
9042: douta=16'h6b0d;
9043: douta=16'h734f;
9044: douta=16'h52ad;
9045: douta=16'hbd52;
9046: douta=16'hee96;
9047: douta=16'hde36;
9048: douta=16'hbd53;
9049: douta=16'had14;
9050: douta=16'hb556;
9051: douta=16'h9494;
9052: douta=16'h94b4;
9053: douta=16'h8c73;
9054: douta=16'h8433;
9055: douta=16'h8412;
9056: douta=16'h6b70;
9057: douta=16'h632f;
9058: douta=16'h4ace;
9059: douta=16'h7b2c;
9060: douta=16'he635;
9061: douta=16'h6bb1;
9062: douta=16'h52cd;
9063: douta=16'h320b;
9064: douta=16'h1905;
9065: douta=16'h31ea;
9066: douta=16'h2125;
9067: douta=16'h1084;
9068: douta=16'h63d3;
9069: douta=16'h9d7a;
9070: douta=16'h8d18;
9071: douta=16'h63d2;
9072: douta=16'h3187;
9073: douta=16'h5162;
9074: douta=16'h7203;
9075: douta=16'h7244;
9076: douta=16'h7265;
9077: douta=16'h6a25;
9078: douta=16'h6a25;
9079: douta=16'h6a25;
9080: douta=16'h6a05;
9081: douta=16'h61e5;
9082: douta=16'h59e5;
9083: douta=16'h49a6;
9084: douta=16'h41c7;
9085: douta=16'h49e8;
9086: douta=16'h5228;
9087: douta=16'h3987;
9088: douta=16'he58d;
9089: douta=16'he56c;
9090: douta=16'hedcc;
9091: douta=16'h7aa8;
9092: douta=16'hcd54;
9093: douta=16'hac92;
9094: douta=16'hc4b0;
9095: douta=16'he676;
9096: douta=16'hb536;
9097: douta=16'h7c55;
9098: douta=16'h8d18;
9099: douta=16'h1927;
9100: douta=16'h320a;
9101: douta=16'h326d;
9102: douta=16'h3a8d;
9103: douta=16'h3a8d;
9104: douta=16'h3a4c;
9105: douta=16'h3a4c;
9106: douta=16'h29ea;
9107: douta=16'h3a6c;
9108: douta=16'h3a6c;
9109: douta=16'h3a8c;
9110: douta=16'h3a4c;
9111: douta=16'h3a6b;
9112: douta=16'h530f;
9113: douta=16'h636f;
9114: douta=16'h636f;
9115: douta=16'h634f;
9116: douta=16'h532e;
9117: douta=16'h532e;
9118: douta=16'h5b4f;
9119: douta=16'h534f;
9120: douta=16'h534f;
9121: douta=16'h5b4f;
9122: douta=16'h63d1;
9123: douta=16'h5b6f;
9124: douta=16'h6390;
9125: douta=16'h638f;
9126: douta=16'h634e;
9127: douta=16'h6bd0;
9128: douta=16'h6baf;
9129: douta=16'h736e;
9130: douta=16'h732d;
9131: douta=16'h72cb;
9132: douta=16'h62ab;
9133: douta=16'hde55;
9134: douta=16'hb514;
9135: douta=16'hc574;
9136: douta=16'hbd76;
9137: douta=16'h9d17;
9138: douta=16'h94b6;
9139: douta=16'h7bf2;
9140: douta=16'h7bf1;
9141: douta=16'h7bf1;
9142: douta=16'h6b6f;
9143: douta=16'h4a6c;
9144: douta=16'he614;
9145: douta=16'hd593;
9146: douta=16'hb4f4;
9147: douta=16'h9cd5;
9148: douta=16'h8433;
9149: douta=16'h6b90;
9150: douta=16'h736e;
9151: douta=16'h3a2b;
9152: douta=16'h29ca;
9153: douta=16'h93f0;
9154: douta=16'h8412;
9155: douta=16'h424c;
9156: douta=16'h732d;
9157: douta=16'h6b0c;
9158: douta=16'h72ec;
9159: douta=16'h522a;
9160: douta=16'h3987;
9161: douta=16'hc511;
9162: douta=16'hb4d3;
9163: douta=16'h73d2;
9164: douta=16'h8c53;
9165: douta=16'h7bf2;
9166: douta=16'h9493;
9167: douta=16'h3a6d;
9168: douta=16'h7390;
9169: douta=16'h6b4e;
9170: douta=16'h734f;
9171: douta=16'hd5d4;
9172: douta=16'hde56;
9173: douta=16'hde15;
9174: douta=16'hb555;
9175: douta=16'h8c51;
9176: douta=16'h8c11;
9177: douta=16'h9c93;
9178: douta=16'ha4f5;
9179: douta=16'h9474;
9180: douta=16'h8433;
9181: douta=16'h83f2;
9182: douta=16'h736f;
9183: douta=16'h6b90;
9184: douta=16'h62ed;
9185: douta=16'h6aeb;
9186: douta=16'had10;
9187: douta=16'hde34;
9188: douta=16'hcd94;
9189: douta=16'h7c13;
9190: douta=16'h6b90;
9191: douta=16'h4aef;
9192: douta=16'h428e;
9193: douta=16'h29ca;
9194: douta=16'h2126;
9195: douta=16'h2988;
9196: douta=16'h1906;
9197: douta=16'h9d59;
9198: douta=16'h7cd8;
9199: douta=16'h2904;
9200: douta=16'h8264;
9201: douta=16'h7a44;
9202: douta=16'h7a45;
9203: douta=16'h7245;
9204: douta=16'h6a25;
9205: douta=16'h6a24;
9206: douta=16'h6a05;
9207: douta=16'h6205;
9208: douta=16'h61e5;
9209: douta=16'h61e5;
9210: douta=16'h59e5;
9211: douta=16'h51c6;
9212: douta=16'h4144;
9213: douta=16'h5208;
9214: douta=16'h49e7;
9215: douta=16'h41c8;
9216: douta=16'he58d;
9217: douta=16'he56c;
9218: douta=16'hedad;
9219: douta=16'h7a66;
9220: douta=16'hc512;
9221: douta=16'hbcb1;
9222: douta=16'hff18;
9223: douta=16'he697;
9224: douta=16'h8434;
9225: douta=16'h8496;
9226: douta=16'h2147;
9227: douta=16'h10e5;
9228: douta=16'h29ca;
9229: douta=16'h2a0c;
9230: douta=16'h324d;
9231: douta=16'h3a6d;
9232: douta=16'h3a8d;
9233: douta=16'h3a6d;
9234: douta=16'h29ea;
9235: douta=16'h2a0b;
9236: douta=16'h324c;
9237: douta=16'h3a8d;
9238: douta=16'h3a6c;
9239: douta=16'h2125;
9240: douta=16'h2125;
9241: douta=16'h31a7;
9242: douta=16'h31c8;
9243: douta=16'h2987;
9244: douta=16'h2146;
9245: douta=16'h2967;
9246: douta=16'h42ac;
9247: douta=16'h5350;
9248: douta=16'h42cd;
9249: douta=16'h530e;
9250: douta=16'h5b4f;
9251: douta=16'h5b4e;
9252: douta=16'h5b4f;
9253: douta=16'h5b4e;
9254: douta=16'h6b90;
9255: douta=16'h638f;
9256: douta=16'h638f;
9257: douta=16'h6b8f;
9258: douta=16'h6b90;
9259: douta=16'h6b90;
9260: douta=16'h532e;
9261: douta=16'hcdb6;
9262: douta=16'hb556;
9263: douta=16'hbd96;
9264: douta=16'ha4f5;
9265: douta=16'h9cd6;
9266: douta=16'h7390;
9267: douta=16'h7bd1;
9268: douta=16'h7bd0;
9269: douta=16'h732e;
9270: douta=16'h5a8c;
9271: douta=16'hf6b4;
9272: douta=16'hacf4;
9273: douta=16'h9cd6;
9274: douta=16'h8453;
9275: douta=16'h8413;
9276: douta=16'h6b70;
9277: douta=16'h62cc;
9278: douta=16'h62ec;
9279: douta=16'h5a49;
9280: douta=16'h62cd;
9281: douta=16'h8c94;
9282: douta=16'h6b4f;
9283: douta=16'h62cd;
9284: douta=16'h424b;
9285: douta=16'h29a8;
9286: douta=16'h524a;
9287: douta=16'h730c;
9288: douta=16'h94b4;
9289: douta=16'h94b5;
9290: douta=16'h94b5;
9291: douta=16'h7c13;
9292: douta=16'h52ef;
9293: douta=16'h52ce;
9294: douta=16'h83b0;
9295: douta=16'h632e;
9296: douta=16'h8bef;
9297: douta=16'he656;
9298: douta=16'hd616;
9299: douta=16'hbd74;
9300: douta=16'hc5b6;
9301: douta=16'had15;
9302: douta=16'ha515;
9303: douta=16'ha4f5;
9304: douta=16'h9cd3;
9305: douta=16'h8c52;
9306: douta=16'h8411;
9307: douta=16'h7bf1;
9308: douta=16'h8412;
9309: douta=16'h7bf2;
9310: douta=16'h62cc;
9311: douta=16'h1061;
9312: douta=16'hcdb2;
9313: douta=16'hd5f5;
9314: douta=16'hcdb5;
9315: douta=16'hb535;
9316: douta=16'ha515;
9317: douta=16'h7c34;
9318: douta=16'h7c55;
9319: douta=16'h5b31;
9320: douta=16'h42cf;
9321: douta=16'h3a4d;
9322: douta=16'h4aae;
9323: douta=16'h29a8;
9324: douta=16'h0884;
9325: douta=16'h2968;
9326: douta=16'h42ae;
9327: douta=16'h8284;
9328: douta=16'h7a64;
9329: douta=16'h7a44;
9330: douta=16'h7245;
9331: douta=16'h7224;
9332: douta=16'h6a24;
9333: douta=16'h6204;
9334: douta=16'h61e4;
9335: douta=16'h61e5;
9336: douta=16'h61e5;
9337: douta=16'h61e5;
9338: douta=16'h59c5;
9339: douta=16'h51a5;
9340: douta=16'h4964;
9341: douta=16'h4123;
9342: douta=16'h4165;
9343: douta=16'h630c;
9344: douta=16'hed6b;
9345: douta=16'he54b;
9346: douta=16'hdd09;
9347: douta=16'h92c8;
9348: douta=16'hd573;
9349: douta=16'hcd92;
9350: douta=16'hf77a;
9351: douta=16'hddf6;
9352: douta=16'h6bd3;
9353: douta=16'h84b7;
9354: douta=16'h73b2;
9355: douta=16'h8496;
9356: douta=16'h9579;
9357: douta=16'h326d;
9358: douta=16'h3aae;
9359: douta=16'h3aae;
9360: douta=16'h3a8e;
9361: douta=16'h3a8d;
9362: douta=16'h21a9;
9363: douta=16'h29ea;
9364: douta=16'h2167;
9365: douta=16'h10a3;
9366: douta=16'h1905;
9367: douta=16'h2967;
9368: douta=16'h39ea;
9369: douta=16'h422a;
9370: douta=16'h422a;
9371: douta=16'h39ea;
9372: douta=16'h31a9;
9373: douta=16'h2146;
9374: douta=16'h10e5;
9375: douta=16'h10e5;
9376: douta=16'h10a4;
9377: douta=16'h42ee;
9378: douta=16'h4b0d;
9379: douta=16'h52ed;
9380: douta=16'h5b4e;
9381: douta=16'h5b0e;
9382: douta=16'h6b90;
9383: douta=16'h638f;
9384: douta=16'h6bd0;
9385: douta=16'h6bb0;
9386: douta=16'h634e;
9387: douta=16'h6bb0;
9388: douta=16'h636e;
9389: douta=16'h638f;
9390: douta=16'h73af;
9391: douta=16'h9cb3;
9392: douta=16'had14;
9393: douta=16'h9493;
9394: douta=16'h8412;
9395: douta=16'h7bf1;
9396: douta=16'h526b;
9397: douta=16'h93ee;
9398: douta=16'he655;
9399: douta=16'hacf5;
9400: douta=16'h8c95;
9401: douta=16'h8c95;
9402: douta=16'h736f;
9403: douta=16'h7b90;
9404: douta=16'h5aab;
9405: douta=16'h62cc;
9406: douta=16'h62cb;
9407: douta=16'hacd3;
9408: douta=16'h4a2a;
9409: douta=16'h6b4f;
9410: douta=16'h524a;
9411: douta=16'h2988;
9412: douta=16'h41e8;
9413: douta=16'h2968;
9414: douta=16'hd5b2;
9415: douta=16'hbd13;
9416: douta=16'h7c13;
9417: douta=16'h6370;
9418: douta=16'h83f2;
9419: douta=16'h6b2f;
9420: douta=16'h62ed;
9421: douta=16'h736f;
9422: douta=16'h7bb0;
9423: douta=16'hd5f4;
9424: douta=16'hde77;
9425: douta=16'hcdf7;
9426: douta=16'hc5d7;
9427: douta=16'hc5b6;
9428: douta=16'had56;
9429: douta=16'ha515;
9430: douta=16'h7c34;
9431: douta=16'h9472;
9432: douta=16'h9473;
9433: douta=16'h8432;
9434: douta=16'h83f1;
9435: douta=16'h62ee;
9436: douta=16'h6aeb;
9437: douta=16'ha46f;
9438: douta=16'hde13;
9439: douta=16'he634;
9440: douta=16'he655;
9441: douta=16'hde34;
9442: douta=16'hbd33;
9443: douta=16'had14;
9444: douta=16'h9cf6;
9445: douta=16'h7c34;
9446: douta=16'h7455;
9447: douta=16'h63f4;
9448: douta=16'h4b10;
9449: douta=16'h42ae;
9450: douta=16'h2989;
9451: douta=16'h7c54;
9452: douta=16'h1907;
9453: douta=16'h18e5;
9454: douta=16'h1949;
9455: douta=16'h7aa5;
9456: douta=16'h7a85;
9457: douta=16'h7a65;
9458: douta=16'h7a65;
9459: douta=16'h7224;
9460: douta=16'h61e4;
9461: douta=16'h61c4;
9462: douta=16'h59a4;
9463: douta=16'h59e5;
9464: douta=16'h72ea;
9465: douta=16'h8c51;
9466: douta=16'h9d13;
9467: douta=16'h9d13;
9468: douta=16'h8c50;
9469: douta=16'h7b8d;
9470: douta=16'h5a69;
9471: douta=16'h4a27;
9472: douta=16'he507;
9473: douta=16'he4e7;
9474: douta=16'hdcc6;
9475: douta=16'hf73b;
9476: douta=16'hee96;
9477: douta=16'hee56;
9478: douta=16'hf6f8;
9479: douta=16'hbd95;
9480: douta=16'h8454;
9481: douta=16'h7c54;
9482: douta=16'h8c75;
9483: douta=16'h94f8;
9484: douta=16'h3a8d;
9485: douta=16'h2a0c;
9486: douta=16'h326d;
9487: douta=16'h42af;
9488: douta=16'h3a8e;
9489: douta=16'h326d;
9490: douta=16'h1967;
9491: douta=16'h2147;
9492: douta=16'h18e5;
9493: douta=16'h2146;
9494: douta=16'h31ea;
9495: douta=16'h31c9;
9496: douta=16'h39ea;
9497: douta=16'h424b;
9498: douta=16'h4a8c;
9499: douta=16'h424c;
9500: douta=16'h426d;
9501: douta=16'h4acf;
9502: douta=16'h3a4c;
9503: douta=16'h420b;
9504: douta=16'h10e5;
9505: douta=16'h10c5;
9506: douta=16'h29c9;
9507: douta=16'h4acd;
9508: douta=16'h530d;
9509: douta=16'h530d;
9510: douta=16'h5b4e;
9511: douta=16'h5b4f;
9512: douta=16'h636f;
9513: douta=16'h6b8f;
9514: douta=16'h634f;
9515: douta=16'h6bb0;
9516: douta=16'h6bb0;
9517: douta=16'h73d0;
9518: douta=16'h73cf;
9519: douta=16'h6b8f;
9520: douta=16'h73cf;
9521: douta=16'h6b6d;
9522: douta=16'h7bef;
9523: douta=16'h738e;
9524: douta=16'hcd33;
9525: douta=16'h94d5;
9526: douta=16'ha4f6;
9527: douta=16'h8c53;
9528: douta=16'h73b0;
9529: douta=16'h7b90;
9530: douta=16'h732e;
9531: douta=16'h736e;
9532: douta=16'h62ab;
9533: douta=16'hacb2;
9534: douta=16'h73f2;
9535: douta=16'h8433;
9536: douta=16'h3a0a;
9537: douta=16'h62ac;
9538: douta=16'h62ab;
9539: douta=16'h6289;
9540: douta=16'h6aab;
9541: douta=16'h7c34;
9542: douta=16'ha515;
9543: douta=16'h8474;
9544: douta=16'h632f;
9545: douta=16'h52ae;
9546: douta=16'h736f;
9547: douta=16'h62ed;
9548: douta=16'h4a6c;
9549: douta=16'hde35;
9550: douta=16'hde56;
9551: douta=16'hde56;
9552: douta=16'hc5b6;
9553: douta=16'hb577;
9554: douta=16'h8c94;
9555: douta=16'h9d16;
9556: douta=16'ha557;
9557: douta=16'h9494;
9558: douta=16'h8432;
9559: douta=16'h6b90;
9560: douta=16'h6b70;
9561: douta=16'h524a;
9562: douta=16'h62c9;
9563: douta=16'h49e7;
9564: douta=16'hac90;
9565: douta=16'hbd12;
9566: douta=16'he676;
9567: douta=16'hc574;
9568: douta=16'hbd34;
9569: douta=16'ha4d5;
9570: douta=16'h9cd5;
9571: douta=16'h94d5;
9572: douta=16'h8c75;
9573: douta=16'h7433;
9574: douta=16'h73f3;
9575: douta=16'h7434;
9576: douta=16'h4b10;
9577: douta=16'h29eb;
9578: douta=16'h5b0f;
9579: douta=16'h4b0f;
9580: douta=16'h31ea;
9581: douta=16'h2127;
9582: douta=16'h10e5;
9583: douta=16'h7a24;
9584: douta=16'h7a86;
9585: douta=16'h936a;
9586: douta=16'ha44d;
9587: douta=16'hbd51;
9588: douta=16'hc592;
9589: douta=16'had0f;
9590: douta=16'h942d;
9591: douta=16'h7b4a;
9592: douta=16'h6267;
9593: douta=16'h5184;
9594: douta=16'h5164;
9595: douta=16'h51a5;
9596: douta=16'h5185;
9597: douta=16'h4985;
9598: douta=16'h49a5;
9599: douta=16'h4185;
9600: douta=16'hd484;
9601: douta=16'hd484;
9602: douta=16'hee55;
9603: douta=16'hff3a;
9604: douta=16'heeb8;
9605: douta=16'hff3a;
9606: douta=16'hee98;
9607: douta=16'h8433;
9608: douta=16'h8c75;
9609: douta=16'h6b2f;
9610: douta=16'h8496;
9611: douta=16'h9518;
9612: douta=16'h08e6;
9613: douta=16'h21ca;
9614: douta=16'h324d;
9615: douta=16'h3a6d;
9616: douta=16'h324d;
9617: douta=16'h42af;
9618: douta=16'h1948;
9619: douta=16'h1947;
9620: douta=16'h18e5;
9621: douta=16'h1927;
9622: douta=16'h29a8;
9623: douta=16'h31c9;
9624: douta=16'h422c;
9625: douta=16'h426c;
9626: douta=16'h424c;
9627: douta=16'h4a8c;
9628: douta=16'h426c;
9629: douta=16'h424c;
9630: douta=16'h39eb;
9631: douta=16'h31c9;
9632: douta=16'h31a9;
9633: douta=16'h29a8;
9634: douta=16'h10a4;
9635: douta=16'h320a;
9636: douta=16'h52cd;
9637: douta=16'h52cd;
9638: douta=16'h4acd;
9639: douta=16'h5b2e;
9640: douta=16'h530e;
9641: douta=16'h5b2e;
9642: douta=16'h634e;
9643: douta=16'h636f;
9644: douta=16'h6b8f;
9645: douta=16'h73f0;
9646: douta=16'h6b6e;
9647: douta=16'h634d;
9648: douta=16'h632d;
9649: douta=16'h6b6e;
9650: douta=16'h738f;
9651: douta=16'h7baf;
9652: douta=16'h7baf;
9653: douta=16'h736d;
9654: douta=16'h8bef;
9655: douta=16'h8bcf;
9656: douta=16'h83af;
9657: douta=16'h736d;
9658: douta=16'h732c;
9659: douta=16'h836d;
9660: douta=16'h9c92;
9661: douta=16'h8c32;
9662: douta=16'h734e;
9663: douta=16'h732d;
9664: douta=16'h6aeb;
9665: douta=16'h6acb;
9666: douta=16'h6269;
9667: douta=16'hc574;
9668: douta=16'h7bf1;
9669: douta=16'h9495;
9670: douta=16'h94b5;
9671: douta=16'h7bf1;
9672: douta=16'h7390;
9673: douta=16'h734f;
9674: douta=16'h52ad;
9675: douta=16'hb535;
9676: douta=16'hde77;
9677: douta=16'hd5f6;
9678: douta=16'h9cd5;
9679: douta=16'had56;
9680: douta=16'h94b5;
9681: douta=16'h7bf1;
9682: douta=16'h8412;
9683: douta=16'h7bf2;
9684: douta=16'h94d5;
9685: douta=16'h7c12;
9686: douta=16'h6b91;
9687: douta=16'h524a;
9688: douta=16'hcdb4;
9689: douta=16'hddf4;
9690: douta=16'he656;
9691: douta=16'hde35;
9692: douta=16'hf6b7;
9693: douta=16'hacd1;
9694: douta=16'ha451;
9695: douta=16'hacb4;
9696: douta=16'hbd54;
9697: douta=16'h9cb4;
9698: douta=16'h94b4;
9699: douta=16'h8453;
9700: douta=16'h73f2;
9701: douta=16'h73b2;
9702: douta=16'h5b50;
9703: douta=16'h5b51;
9704: douta=16'h4aee;
9705: douta=16'h6b2d;
9706: douta=16'h3a4c;
9707: douta=16'h52cc;
9708: douta=16'h29ca;
9709: douta=16'h1926;
9710: douta=16'h18e5;
9711: douta=16'h83cc;
9712: douta=16'h9bca;
9713: douta=16'h82c7;
9714: douta=16'h7225;
9715: douta=16'h61c4;
9716: douta=16'h61e5;
9717: douta=16'h61e5;
9718: douta=16'h61e4;
9719: douta=16'h59e5;
9720: douta=16'h59e5;
9721: douta=16'h51a5;
9722: douta=16'h51a5;
9723: douta=16'h4985;
9724: douta=16'h4985;
9725: douta=16'h49a5;
9726: douta=16'h4985;
9727: douta=16'h4186;
9728: douta=16'hcd4c;
9729: douta=16'haae0;
9730: douta=16'hff1a;
9731: douta=16'hff3b;
9732: douta=16'hf6d8;
9733: douta=16'hff9c;
9734: douta=16'hde17;
9735: douta=16'h8c34;
9736: douta=16'h8c95;
9737: douta=16'h7bd2;
9738: douta=16'h94d6;
9739: douta=16'h9d18;
9740: douta=16'h2147;
9741: douta=16'h2189;
9742: douta=16'h29ca;
9743: douta=16'h21ca;
9744: douta=16'h29ea;
9745: douta=16'h29ca;
9746: douta=16'h2168;
9747: douta=16'h1106;
9748: douta=16'h2168;
9749: douta=16'h2168;
9750: douta=16'h2147;
9751: douta=16'h31a9;
9752: douta=16'h428d;
9753: douta=16'h3a0b;
9754: douta=16'h4a6c;
9755: douta=16'h426c;
9756: douta=16'h3a2b;
9757: douta=16'h424c;
9758: douta=16'h4a8d;
9759: douta=16'h31c9;
9760: douta=16'h31a8;
9761: douta=16'h2967;
9762: douta=16'h2126;
9763: douta=16'h2167;
9764: douta=16'h4aad;
9765: douta=16'h4aed;
9766: douta=16'h4aac;
9767: douta=16'h530d;
9768: douta=16'h530d;
9769: douta=16'h4aac;
9770: douta=16'h4aac;
9771: douta=16'h5aed;
9772: douta=16'h634e;
9773: douta=16'h6b8f;
9774: douta=16'h73d0;
9775: douta=16'h6b8f;
9776: douta=16'h632d;
9777: douta=16'h5acb;
9778: douta=16'h6b2d;
9779: douta=16'h6b6d;
9780: douta=16'h6b4d;
9781: douta=16'h6aeb;
9782: douta=16'h738e;
9783: douta=16'h736e;
9784: douta=16'h732d;
9785: douta=16'h734d;
9786: douta=16'h7b6e;
9787: douta=16'h7b4d;
9788: douta=16'h7b8e;
9789: douta=16'h8bcf;
9790: douta=16'h834d;
9791: douta=16'h7b0b;
9792: douta=16'h834b;
9793: douta=16'h9471;
9794: douta=16'h836f;
9795: douta=16'h734e;
9796: douta=16'h7bb0;
9797: douta=16'h630e;
9798: douta=16'h736f;
9799: douta=16'h732d;
9800: douta=16'h6aed;
9801: douta=16'h734e;
9802: douta=16'hd5d4;
9803: douta=16'hb535;
9804: douta=16'hc5b6;
9805: douta=16'hb557;
9806: douta=16'h9cd6;
9807: douta=16'h8453;
9808: douta=16'h7bf2;
9809: douta=16'h6b70;
9810: douta=16'h6b6f;
9811: douta=16'h7370;
9812: douta=16'h734f;
9813: douta=16'h49e8;
9814: douta=16'he615;
9815: douta=16'hbd13;
9816: douta=16'he676;
9817: douta=16'hde35;
9818: douta=16'hcd93;
9819: douta=16'hacf4;
9820: douta=16'h8c52;
9821: douta=16'h8c12;
9822: douta=16'ha4b3;
9823: douta=16'h9cb3;
9824: douta=16'h8c73;
9825: douta=16'h83f1;
9826: douta=16'h7390;
9827: douta=16'h7390;
9828: douta=16'h6b70;
9829: douta=16'h6bb2;
9830: douta=16'h4a49;
9831: douta=16'h5a88;
9832: douta=16'hbd11;
9833: douta=16'h9451;
9834: douta=16'h630d;
9835: douta=16'h5b4f;
9836: douta=16'h29a8;
9837: douta=16'h52ad;
9838: douta=16'h2147;
9839: douta=16'h10c5;
9840: douta=16'h8286;
9841: douta=16'h7a45;
9842: douta=16'h7225;
9843: douta=16'h7225;
9844: douta=16'h6a05;
9845: douta=16'h6205;
9846: douta=16'h61e5;
9847: douta=16'h59e5;
9848: douta=16'h59c5;
9849: douta=16'h51c5;
9850: douta=16'h51a5;
9851: douta=16'h51a5;
9852: douta=16'h49a6;
9853: douta=16'h49a5;
9854: douta=16'h4185;
9855: douta=16'h4165;
9856: douta=16'hcd2b;
9857: douta=16'hf6b7;
9858: douta=16'hf6d8;
9859: douta=16'hff3a;
9860: douta=16'hf6f9;
9861: douta=16'hf718;
9862: douta=16'h9cb4;
9863: douta=16'h8c94;
9864: douta=16'h8cb6;
9865: douta=16'h8c74;
9866: douta=16'h94d6;
9867: douta=16'h31e9;
9868: douta=16'h18e4;
9869: douta=16'h18e5;
9870: douta=16'h2168;
9871: douta=16'h1926;
9872: douta=16'h1906;
9873: douta=16'h1967;
9874: douta=16'h1947;
9875: douta=16'h1148;
9876: douta=16'h2189;
9877: douta=16'h1906;
9878: douta=16'h29ca;
9879: douta=16'h18e5;
9880: douta=16'h31ea;
9881: douta=16'h2148;
9882: douta=16'h3a0a;
9883: douta=16'h5b30;
9884: douta=16'h322c;
9885: douta=16'h2988;
9886: douta=16'h3a2b;
9887: douta=16'h31a9;
9888: douta=16'h41ea;
9889: douta=16'h31c9;
9890: douta=16'h31c8;
9891: douta=16'h29ea;
9892: douta=16'h3a6b;
9893: douta=16'h4aad;
9894: douta=16'h52cd;
9895: douta=16'h52ed;
9896: douta=16'h530d;
9897: douta=16'h634e;
9898: douta=16'h5b0d;
9899: douta=16'h5b2d;
9900: douta=16'h632d;
9901: douta=16'h52ab;
9902: douta=16'h5aab;
9903: douta=16'h528a;
9904: douta=16'h632d;
9905: douta=16'h5acb;
9906: douta=16'h62cb;
9907: douta=16'h630c;
9908: douta=16'h62cb;
9909: douta=16'h62cb;
9910: douta=16'h6b0c;
9911: douta=16'h734d;
9912: douta=16'h7b8e;
9913: douta=16'h7baf;
9914: douta=16'h8c51;
9915: douta=16'h83cf;
9916: douta=16'h83cf;
9917: douta=16'h8431;
9918: douta=16'ha557;
9919: douta=16'hb533;
9920: douta=16'hcdb3;
9921: douta=16'hccaa;
9922: douta=16'hdca7;
9923: douta=16'hc468;
9924: douta=16'h940e;
9925: douta=16'h7b6f;
9926: douta=16'h6b2e;
9927: douta=16'h7b4d;
9928: douta=16'hee97;
9929: douta=16'he697;
9930: douta=16'hcdf6;
9931: douta=16'hbd96;
9932: douta=16'ha517;
9933: douta=16'h94d5;
9934: douta=16'h8412;
9935: douta=16'h736f;
9936: douta=16'h736f;
9937: douta=16'h6b2e;
9938: douta=16'h5acd;
9939: douta=16'h8bee;
9940: douta=16'hcd91;
9941: douta=16'he656;
9942: douta=16'hde35;
9943: douta=16'hddf5;
9944: douta=16'had14;
9945: douta=16'hbd95;
9946: douta=16'ha4f5;
9947: douta=16'h8c74;
9948: douta=16'h73b0;
9949: douta=16'h7bd1;
9950: douta=16'h7390;
9951: douta=16'h6b4f;
9952: douta=16'h6b2d;
9953: douta=16'h5acc;
9954: douta=16'h632e;
9955: douta=16'h5a8a;
9956: douta=16'h62cb;
9957: douta=16'h942e;
9958: douta=16'haccf;
9959: douta=16'hd5d3;
9960: douta=16'hde14;
9961: douta=16'hacf4;
9962: douta=16'h7c12;
9963: douta=16'h5b30;
9964: douta=16'h3a4c;
9965: douta=16'h31ea;
9966: douta=16'h3a2b;
9967: douta=16'h1906;
9968: douta=16'h1106;
9969: douta=16'h8286;
9970: douta=16'h7225;
9971: douta=16'h6a04;
9972: douta=16'h61e5;
9973: douta=16'h61e4;
9974: douta=16'h59e5;
9975: douta=16'h59c5;
9976: douta=16'h59c5;
9977: douta=16'h51c5;
9978: douta=16'h51c6;
9979: douta=16'h51c5;
9980: douta=16'h49a6;
9981: douta=16'h49a6;
9982: douta=16'h4185;
9983: douta=16'h41a6;
9984: douta=16'he674;
9985: douta=16'hf71a;
9986: douta=16'hf71a;
9987: douta=16'hf739;
9988: douta=16'hff3a;
9989: douta=16'hde57;
9990: douta=16'ha4f5;
9991: douta=16'h94b5;
9992: douta=16'h9494;
9993: douta=16'h94d5;
9994: douta=16'h94d6;
9995: douta=16'h63b3;
9996: douta=16'h7436;
9997: douta=16'h42ae;
9998: douta=16'h10c4;
9999: douta=16'h1926;
10000: douta=16'h1927;
10001: douta=16'h1947;
10002: douta=16'h1948;
10003: douta=16'h1948;
10004: douta=16'h2168;
10005: douta=16'h1926;
10006: douta=16'h10c5;
10007: douta=16'h2188;
10008: douta=16'h29ca;
10009: douta=16'h1906;
10010: douta=16'h2967;
10011: douta=16'h2988;
10012: douta=16'h2147;
10013: douta=16'h3189;
10014: douta=16'h2988;
10015: douta=16'h3188;
10016: douta=16'h2988;
10017: douta=16'h31e9;
10018: douta=16'h31e9;
10019: douta=16'h322a;
10020: douta=16'h3a4b;
10021: douta=16'h426b;
10022: douta=16'h428c;
10023: douta=16'h4a8c;
10024: douta=16'h52cd;
10025: douta=16'h52ed;
10026: douta=16'h5b2e;
10027: douta=16'h5acc;
10028: douta=16'h632d;
10029: douta=16'h5aec;
10030: douta=16'h5aab;
10031: douta=16'h630c;
10032: douta=16'h4a48;
10033: douta=16'h5a8a;
10034: douta=16'h734d;
10035: douta=16'h62ec;
10036: douta=16'h736d;
10037: douta=16'h83ef;
10038: douta=16'h8c31;
10039: douta=16'h8411;
10040: douta=16'ha555;
10041: douta=16'hce38;
10042: douta=16'hcd6f;
10043: douta=16'he5b0;
10044: douta=16'hd467;
10045: douta=16'hc3e1;
10046: douta=16'hcc24;
10047: douta=16'hcc25;
10048: douta=16'hcc65;
10049: douta=16'hcc66;
10050: douta=16'hd467;
10051: douta=16'hd466;
10052: douta=16'hd466;
10053: douta=16'hd466;
10054: douta=16'hd465;
10055: douta=16'hb4d2;
10056: douta=16'hbd97;
10057: douta=16'had16;
10058: douta=16'had57;
10059: douta=16'hb596;
10060: douta=16'h8c53;
10061: douta=16'h7bf2;
10062: douta=16'h8411;
10063: douta=16'h6b2e;
10064: douta=16'h5acc;
10065: douta=16'hacd2;
10066: douta=16'ha4b0;
10067: douta=16'hcdf4;
10068: douta=16'hcd94;
10069: douta=16'hd5f4;
10070: douta=16'hc576;
10071: douta=16'hb556;
10072: douta=16'hb535;
10073: douta=16'h9cf5;
10074: douta=16'h9cb5;
10075: douta=16'h6b4f;
10076: douta=16'h7bd1;
10077: douta=16'h83f1;
10078: douta=16'h632f;
10079: douta=16'h630e;
10080: douta=16'h4a29;
10081: douta=16'h3123;
10082: douta=16'h5248;
10083: douta=16'h5a89;
10084: douta=16'h732b;
10085: douta=16'hcdd3;
10086: douta=16'he656;
10087: douta=16'hde35;
10088: douta=16'hcd73;
10089: douta=16'ha514;
10090: douta=16'h8495;
10091: douta=16'h5b50;
10092: douta=16'h4ace;
10093: douta=16'h3a6c;
10094: douta=16'h2168;
10095: douta=16'h2988;
10096: douta=16'h10c5;
10097: douta=16'h3965;
10098: douta=16'h7245;
10099: douta=16'h6a25;
10100: douta=16'h6205;
10101: douta=16'h61e4;
10102: douta=16'h59e5;
10103: douta=16'h59c5;
10104: douta=16'h51a5;
10105: douta=16'h59e6;
10106: douta=16'h51c5;
10107: douta=16'h51c5;
10108: douta=16'h49a6;
10109: douta=16'h49a6;
10110: douta=16'h4185;
10111: douta=16'h4165;
10112: douta=16'hf6f7;
10113: douta=16'hf6f9;
10114: douta=16'hff3a;
10115: douta=16'hf6f9;
10116: douta=16'hff9c;
10117: douta=16'hc5b6;
10118: douta=16'h8c53;
10119: douta=16'h94b5;
10120: douta=16'h9473;
10121: douta=16'ha517;
10122: douta=16'h94b6;
10123: douta=16'h7435;
10124: douta=16'h6c34;
10125: douta=16'h8497;
10126: douta=16'h2a2a;
10127: douta=16'h1105;
10128: douta=16'h1926;
10129: douta=16'h1947;
10130: douta=16'h1127;
10131: douta=16'h1927;
10132: douta=16'h1947;
10133: douta=16'h1926;
10134: douta=16'h2189;
10135: douta=16'h1082;
10136: douta=16'h1968;
10137: douta=16'h2168;
10138: douta=16'h1946;
10139: douta=16'h18e4;
10140: douta=16'h322b;
10141: douta=16'h18a1;
10142: douta=16'h0000;
10143: douta=16'h0821;
10144: douta=16'h18e4;
10145: douta=16'h1905;
10146: douta=16'h31ea;
10147: douta=16'h3a0a;
10148: douta=16'h3a2a;
10149: douta=16'h31e9;
10150: douta=16'h31a8;
10151: douta=16'h39c8;
10152: douta=16'h4a6b;
10153: douta=16'h3a09;
10154: douta=16'h4a8b;
10155: douta=16'h4a4a;
10156: douta=16'h4a6a;
10157: douta=16'h638e;
10158: douta=16'h7390;
10159: douta=16'h8473;
10160: douta=16'h6b8f;
10161: douta=16'h6b8f;
10162: douta=16'h93cd;
10163: douta=16'hcd70;
10164: douta=16'hbbc4;
10165: douta=16'hcbe3;
10166: douta=16'hc3c3;
10167: douta=16'hc3e2;
10168: douta=16'hcc25;
10169: douta=16'hcc25;
10170: douta=16'hcc25;
10171: douta=16'hcc45;
10172: douta=16'hcc45;
10173: douta=16'hcc45;
10174: douta=16'hcc45;
10175: douta=16'hcc46;
10176: douta=16'hcc66;
10177: douta=16'hcc46;
10178: douta=16'hcc45;
10179: douta=16'hd466;
10180: douta=16'hd466;
10181: douta=16'hd466;
10182: douta=16'hd465;
10183: douta=16'hd486;
10184: douta=16'hbcaf;
10185: douta=16'h9c51;
10186: douta=16'h9451;
10187: douta=16'ha4f5;
10188: douta=16'h8c11;
10189: douta=16'h73d0;
10190: douta=16'h6b4f;
10191: douta=16'h732e;
10192: douta=16'he677;
10193: douta=16'hbd52;
10194: douta=16'he6b7;
10195: douta=16'hde15;
10196: douta=16'hd5d5;
10197: douta=16'hb535;
10198: douta=16'h9494;
10199: douta=16'h8412;
10200: douta=16'h8c33;
10201: douta=16'h9494;
10202: douta=16'h8c74;
10203: douta=16'h630e;
10204: douta=16'h632e;
10205: douta=16'h632f;
10206: douta=16'h41e8;
10207: douta=16'h5228;
10208: douta=16'hcd52;
10209: douta=16'hc550;
10210: douta=16'hde14;
10211: douta=16'he676;
10212: douta=16'he676;
10213: douta=16'he656;
10214: douta=16'hde35;
10215: douta=16'hcdb5;
10216: douta=16'h9cf5;
10217: douta=16'h94d5;
10218: douta=16'h8475;
10219: douta=16'h6bf3;
10220: douta=16'h6bb2;
10221: douta=16'h4b10;
10222: douta=16'h530f;
10223: douta=16'h1106;
10224: douta=16'h2168;
10225: douta=16'h10c6;
10226: douta=16'h7226;
10227: douta=16'h6a24;
10228: douta=16'h6a05;
10229: douta=16'h6205;
10230: douta=16'h59e5;
10231: douta=16'h59c5;
10232: douta=16'h59c5;
10233: douta=16'h51c6;
10234: douta=16'h51c5;
10235: douta=16'h49c6;
10236: douta=16'h49a6;
10237: douta=16'h4985;
10238: douta=16'h4186;
10239: douta=16'h4165;
10240: douta=16'hff1a;
10241: douta=16'hf6f9;
10242: douta=16'hf6f9;
10243: douta=16'hff19;
10244: douta=16'heeb7;
10245: douta=16'had16;
10246: douta=16'ha516;
10247: douta=16'ha516;
10248: douta=16'ha4d5;
10249: douta=16'h9cd6;
10250: douta=16'h6bf3;
10251: douta=16'h7414;
10252: douta=16'h7c96;
10253: douta=16'h8497;
10254: douta=16'h8497;
10255: douta=16'h84f8;
10256: douta=16'h29ca;
10257: douta=16'h1105;
10258: douta=16'h1106;
10259: douta=16'h1126;
10260: douta=16'h10e5;
10261: douta=16'h1126;
10262: douta=16'h2147;
10263: douta=16'h2188;
10264: douta=16'h10c4;
10265: douta=16'h2126;
10266: douta=16'h3186;
10267: douta=16'h10c5;
10268: douta=16'h2126;
10269: douta=16'h18a3;
10270: douta=16'h1061;
10271: douta=16'h18c4;
10272: douta=16'h29a9;
10273: douta=16'h31ea;
10274: douta=16'h2968;
10275: douta=16'h3a2a;
10276: douta=16'h3209;
10277: douta=16'h424b;
10278: douta=16'h422b;
10279: douta=16'h422a;
10280: douta=16'h4acd;
10281: douta=16'h4a8c;
10282: douta=16'h52ab;
10283: douta=16'h6acb;
10284: douta=16'h7ac8;
10285: douta=16'h92c3;
10286: douta=16'hab23;
10287: douta=16'hb384;
10288: douta=16'hb385;
10289: douta=16'hb3a5;
10290: douta=16'hbba6;
10291: douta=16'hbbc4;
10292: douta=16'hbbc5;
10293: douta=16'hbbe5;
10294: douta=16'hc405;
10295: douta=16'hc404;
10296: douta=16'hc404;
10297: douta=16'hcc46;
10298: douta=16'hcc25;
10299: douta=16'hcc45;
10300: douta=16'hcc25;
10301: douta=16'hcc45;
10302: douta=16'hcc45;
10303: douta=16'hcc45;
10304: douta=16'hcc46;
10305: douta=16'hd466;
10306: douta=16'hcc46;
10307: douta=16'hd445;
10308: douta=16'hd421;
10309: douta=16'hcc22;
10310: douta=16'hd4a9;
10311: douta=16'hddaf;
10312: douta=16'heeb5;
10313: douta=16'hff9a;
10314: douta=16'hc5f5;
10315: douta=16'h836e;
10316: douta=16'h730c;
10317: douta=16'ha490;
10318: douta=16'he656;
10319: douta=16'hcdb3;
10320: douta=16'h9cd6;
10321: douta=16'hcdd6;
10322: douta=16'hb597;
10323: douta=16'h9cd6;
10324: douta=16'h9cd5;
10325: douta=16'h9cb4;
10326: douta=16'h8c33;
10327: douta=16'h7390;
10328: douta=16'h7390;
10329: douta=16'h7bd0;
10330: douta=16'h73b0;
10331: douta=16'h5aac;
10332: douta=16'h49e7;
10333: douta=16'h9c4f;
10334: douta=16'hc550;
10335: douta=16'he635;
10336: douta=16'hcdb2;
10337: douta=16'hd5d4;
10338: douta=16'hd5f4;
10339: douta=16'hddf5;
10340: douta=16'hcdb5;
10341: douta=16'hacd4;
10342: douta=16'ha4d5;
10343: douta=16'h9cf5;
10344: douta=16'h9cf5;
10345: douta=16'h94d5;
10346: douta=16'h7c34;
10347: douta=16'h7434;
10348: douta=16'h6bf3;
10349: douta=16'h5330;
10350: douta=16'h3a2b;
10351: douta=16'h73f1;
10352: douta=16'h2147;
10353: douta=16'h2948;
10354: douta=16'h6a46;
10355: douta=16'h6a25;
10356: douta=16'h6a25;
10357: douta=16'h61e5;
10358: douta=16'h61e5;
10359: douta=16'h59e5;
10360: douta=16'h59e6;
10361: douta=16'h51a5;
10362: douta=16'h51c6;
10363: douta=16'h49c6;
10364: douta=16'h49a6;
10365: douta=16'h4185;
10366: douta=16'h4186;
10367: douta=16'h4186;
10368: douta=16'hf6d8;
10369: douta=16'hff19;
10370: douta=16'hf739;
10371: douta=16'hff19;
10372: douta=16'hd593;
10373: douta=16'ha4d5;
10374: douta=16'ha536;
10375: douta=16'ha4f5;
10376: douta=16'h9cb4;
10377: douta=16'h9cd5;
10378: douta=16'h7414;
10379: douta=16'h7434;
10380: douta=16'h7435;
10381: douta=16'h7c76;
10382: douta=16'h8497;
10383: douta=16'h73f3;
10384: douta=16'h6c35;
10385: douta=16'h10c5;
10386: douta=16'h10e5;
10387: douta=16'h10e5;
10388: douta=16'h10e5;
10389: douta=16'h10e5;
10390: douta=16'h10c4;
10391: douta=16'h1906;
10392: douta=16'h10e5;
10393: douta=16'h18e5;
10394: douta=16'h18e4;
10395: douta=16'h10e4;
10396: douta=16'h1926;
10397: douta=16'h2125;
10398: douta=16'h29a9;
10399: douta=16'h31ea;
10400: douta=16'h322b;
10401: douta=16'h3a2c;
10402: douta=16'h322b;
10403: douta=16'h42ce;
10404: douta=16'h4a4a;
10405: douta=16'h51a5;
10406: douta=16'h61e4;
10407: douta=16'h69e3;
10408: douta=16'h7a24;
10409: douta=16'h8aa4;
10410: douta=16'h92c4;
10411: douta=16'h92e4;
10412: douta=16'h9b05;
10413: douta=16'ha345;
10414: douta=16'hab65;
10415: douta=16'hab85;
10416: douta=16'hb385;
10417: douta=16'hb384;
10418: douta=16'hbba5;
10419: douta=16'hbbc5;
10420: douta=16'hbbe5;
10421: douta=16'hc3e5;
10422: douta=16'hc425;
10423: douta=16'hc426;
10424: douta=16'hd467;
10425: douta=16'hcc25;
10426: douta=16'hcc45;
10427: douta=16'hcc25;
10428: douta=16'hcc24;
10429: douta=16'hc3e2;
10430: douta=16'hcc24;
10431: douta=16'hcca8;
10432: douta=16'hddae;
10433: douta=16'heed7;
10434: douta=16'hf7bc;
10435: douta=16'hf7bb;
10436: douta=16'heed6;
10437: douta=16'hddaf;
10438: douta=16'hd487;
10439: douta=16'hcc22;
10440: douta=16'hd425;
10441: douta=16'hd466;
10442: douta=16'hd466;
10443: douta=16'hd466;
10444: douta=16'hbd95;
10445: douta=16'hd5d5;
10446: douta=16'hcdb5;
10447: douta=16'hde35;
10448: douta=16'ha537;
10449: douta=16'hbd98;
10450: douta=16'h94b5;
10451: douta=16'h7bf2;
10452: douta=16'h7bd1;
10453: douta=16'h7b90;
10454: douta=16'h7b70;
10455: douta=16'h630e;
10456: douta=16'h6b6f;
10457: douta=16'h4a49;
10458: douta=16'h49e7;
10459: douta=16'hc571;
10460: douta=16'hd5d3;
10461: douta=16'hde56;
10462: douta=16'hde55;
10463: douta=16'hde55;
10464: douta=16'ha4b3;
10465: douta=16'hde56;
10466: douta=16'hbd34;
10467: douta=16'hbd14;
10468: douta=16'h9493;
10469: douta=16'h8c93;
10470: douta=16'h8c93;
10471: douta=16'h7c32;
10472: douta=16'h7c13;
10473: douta=16'h7c33;
10474: douta=16'h7c13;
10475: douta=16'h6bf2;
10476: douta=16'h6b91;
10477: douta=16'h6b91;
10478: douta=16'h41a7;
10479: douta=16'h428d;
10480: douta=16'h5b0f;
10481: douta=16'h10e5;
10482: douta=16'h08a5;
10483: douta=16'h7245;
10484: douta=16'h6205;
10485: douta=16'h6205;
10486: douta=16'h59e5;
10487: douta=16'h5a05;
10488: douta=16'h51c5;
10489: douta=16'h51c6;
10490: douta=16'h49a5;
10491: douta=16'h49a6;
10492: douta=16'h49a5;
10493: douta=16'h4185;
10494: douta=16'h4186;
10495: douta=16'h4166;
10496: douta=16'heeb7;
10497: douta=16'hff7b;
10498: douta=16'hf6d8;
10499: douta=16'hff7b;
10500: douta=16'hcdb5;
10501: douta=16'h9453;
10502: douta=16'had56;
10503: douta=16'hb515;
10504: douta=16'ha4f5;
10505: douta=16'h8c95;
10506: douta=16'h7414;
10507: douta=16'h8475;
10508: douta=16'h8476;
10509: douta=16'h8496;
10510: douta=16'h7c54;
10511: douta=16'h8cb7;
10512: douta=16'h0042;
10513: douta=16'h10e5;
10514: douta=16'h10e5;
10515: douta=16'h10c4;
10516: douta=16'h1106;
10517: douta=16'h10e5;
10518: douta=16'h10e6;
10519: douta=16'h10c4;
10520: douta=16'h10e5;
10521: douta=16'h18e4;
10522: douta=16'h2947;
10523: douta=16'h18e5;
10524: douta=16'h29ca;
10525: douta=16'h2168;
10526: douta=16'h3209;
10527: douta=16'h39c8;
10528: douta=16'h4963;
10529: douta=16'h4901;
10530: douta=16'h5183;
10531: douta=16'h59c4;
10532: douta=16'h69e4;
10533: douta=16'h7224;
10534: douta=16'h7224;
10535: douta=16'h7a44;
10536: douta=16'h7a44;
10537: douta=16'h8aa4;
10538: douta=16'h8ac4;
10539: douta=16'h92e4;
10540: douta=16'h9b05;
10541: douta=16'ha344;
10542: douta=16'hab86;
10543: douta=16'hb385;
10544: douta=16'hb385;
10545: douta=16'hb3c5;
10546: douta=16'hbbc5;
10547: douta=16'hbbc6;
10548: douta=16'hbbe5;
10549: douta=16'hbbc3;
10550: douta=16'hbb83;
10551: douta=16'hc3e3;
10552: douta=16'hccaa;
10553: douta=16'hd590;
10554: douta=16'he6d7;
10555: douta=16'hf79b;
10556: douta=16'hef58;
10557: douta=16'he672;
10558: douta=16'hdd6d;
10559: douta=16'hd4a7;
10560: douta=16'hc420;
10561: douta=16'hcc22;
10562: douta=16'hcc45;
10563: douta=16'hd466;
10564: douta=16'hd487;
10565: douta=16'hd486;
10566: douta=16'hd466;
10567: douta=16'hd466;
10568: douta=16'hd466;
10569: douta=16'hd466;
10570: douta=16'hd466;
10571: douta=16'hd486;
10572: douta=16'hd465;
10573: douta=16'ha492;
10574: douta=16'had56;
10575: douta=16'ha537;
10576: douta=16'h9cd6;
10577: douta=16'hb577;
10578: douta=16'h73b1;
10579: douta=16'h7bb1;
10580: douta=16'h6b70;
10581: douta=16'h7370;
10582: douta=16'h5aac;
10583: douta=16'h39a7;
10584: douta=16'h7bae;
10585: douta=16'h9c4f;
10586: douta=16'hd614;
10587: douta=16'hde35;
10588: douta=16'hee97;
10589: douta=16'hde15;
10590: douta=16'hd5f5;
10591: douta=16'hcd94;
10592: douta=16'h9cd4;
10593: douta=16'h8432;
10594: douta=16'ha4d5;
10595: douta=16'h8c52;
10596: douta=16'h8c53;
10597: douta=16'h7bd1;
10598: douta=16'h73b0;
10599: douta=16'h632e;
10600: douta=16'h632e;
10601: douta=16'h630e;
10602: douta=16'h632e;
10603: douta=16'h28e4;
10604: douta=16'h62ca;
10605: douta=16'h83ee;
10606: douta=16'h630e;
10607: douta=16'h52cf;
10608: douta=16'h3a4a;
10609: douta=16'h29a9;
10610: douta=16'h29a9;
10611: douta=16'h10e5;
10612: douta=16'h6226;
10613: douta=16'h6226;
10614: douta=16'h59e5;
10615: douta=16'h59e6;
10616: douta=16'h51c6;
10617: douta=16'h51a5;
10618: douta=16'h51a6;
10619: douta=16'h49a6;
10620: douta=16'h49a6;
10621: douta=16'h41a6;
10622: douta=16'h4186;
10623: douta=16'h3965;
10624: douta=16'hff19;
10625: douta=16'hff7b;
10626: douta=16'hff5a;
10627: douta=16'heeb9;
10628: douta=16'hacf5;
10629: douta=16'ha4d5;
10630: douta=16'had36;
10631: douta=16'hb514;
10632: douta=16'had16;
10633: douta=16'h73f3;
10634: douta=16'h7c34;
10635: douta=16'h7c55;
10636: douta=16'h8476;
10637: douta=16'h8476;
10638: douta=16'h7c54;
10639: douta=16'h322a;
10640: douta=16'h10c4;
10641: douta=16'h0883;
10642: douta=16'h08a4;
10643: douta=16'h10a5;
10644: douta=16'h1967;
10645: douta=16'h2188;
10646: douta=16'h29ca;
10647: douta=16'h29ca;
10648: douta=16'h29c9;
10649: douta=16'h20e4;
10650: douta=16'h2967;
10651: douta=16'h28a1;
10652: douta=16'h30c2;
10653: douta=16'h4143;
10654: douta=16'h4963;
10655: douta=16'h3102;
10656: douta=16'h59c4;
10657: douta=16'h59c4;
10658: douta=16'h6203;
10659: douta=16'h61e4;
10660: douta=16'h7224;
10661: douta=16'h7224;
10662: douta=16'h7224;
10663: douta=16'h7a64;
10664: douta=16'h8284;
10665: douta=16'h8aa4;
10666: douta=16'h8ae4;
10667: douta=16'h9b05;
10668: douta=16'h9b25;
10669: douta=16'ha345;
10670: douta=16'ha303;
10671: douta=16'hab22;
10672: douta=16'hab65;
10673: douta=16'hbc48;
10674: douta=16'hde13;
10675: douta=16'hef18;
10676: douta=16'hf79a;
10677: douta=16'hef17;
10678: douta=16'hde31;
10679: douta=16'hcce9;
10680: douta=16'hc403;
10681: douta=16'hc3e2;
10682: douta=16'hc404;
10683: douta=16'hcc25;
10684: douta=16'hcc46;
10685: douta=16'hcc66;
10686: douta=16'hcc46;
10687: douta=16'hcc45;
10688: douta=16'hcc65;
10689: douta=16'hcc66;
10690: douta=16'hd466;
10691: douta=16'hd466;
10692: douta=16'hd466;
10693: douta=16'hd466;
10694: douta=16'hd466;
10695: douta=16'hd466;
10696: douta=16'hd466;
10697: douta=16'hd467;
10698: douta=16'hd466;
10699: douta=16'hd467;
10700: douta=16'hd466;
10701: douta=16'hd465;
10702: douta=16'h9451;
10703: douta=16'h9453;
10704: douta=16'h9473;
10705: douta=16'h83f1;
10706: douta=16'h7bd1;
10707: douta=16'h7391;
10708: douta=16'h630e;
10709: douta=16'h49e7;
10710: douta=16'h7b4b;
10711: douta=16'hc592;
10712: douta=16'hde55;
10713: douta=16'he6b7;
10714: douta=16'he696;
10715: douta=16'he656;
10716: douta=16'hd616;
10717: douta=16'hcd95;
10718: douta=16'hb555;
10719: douta=16'h9cd5;
10720: douta=16'h9474;
10721: douta=16'h8c53;
10722: douta=16'h8433;
10723: douta=16'h7bf1;
10724: douta=16'h6b4f;
10725: douta=16'h8411;
10726: douta=16'h6b2e;
10727: douta=16'h630c;
10728: douta=16'h5a48;
10729: douta=16'h940d;
10730: douta=16'h8bcd;
10731: douta=16'ha46e;
10732: douta=16'hacb0;
10733: douta=16'hb4d1;
10734: douta=16'h3a2a;
10735: douta=16'h31a8;
10736: douta=16'h2948;
10737: douta=16'h10e6;
10738: douta=16'h10c5;
10739: douta=16'h18e5;
10740: douta=16'h6206;
10741: douta=16'h6205;
10742: douta=16'h59e5;
10743: douta=16'h59e6;
10744: douta=16'h51c5;
10745: douta=16'h49a5;
10746: douta=16'h49a6;
10747: douta=16'h49a6;
10748: douta=16'h4185;
10749: douta=16'h4185;
10750: douta=16'h4186;
10751: douta=16'h4166;
10752: douta=16'hff7b;
10753: douta=16'hffbd;
10754: douta=16'hffdd;
10755: douta=16'he657;
10756: douta=16'ha4b4;
10757: douta=16'hb556;
10758: douta=16'hb535;
10759: douta=16'hbd76;
10760: douta=16'ha4f5;
10761: douta=16'h7413;
10762: douta=16'h8455;
10763: douta=16'h8475;
10764: douta=16'h8475;
10765: douta=16'h7c34;
10766: douta=16'h8c96;
10767: douta=16'h326e;
10768: douta=16'h21cb;
10769: douta=16'h2a2d;
10770: douta=16'h21cb;
10771: douta=16'h18a3;
10772: douta=16'h1881;
10773: douta=16'h1861;
10774: douta=16'h1881;
10775: douta=16'h20a2;
10776: douta=16'h28c2;
10777: douta=16'h2903;
10778: douta=16'h2126;
10779: douta=16'h4123;
10780: douta=16'h3923;
10781: douta=16'h4144;
10782: douta=16'h4964;
10783: douta=16'h51a4;
10784: douta=16'h61c4;
10785: douta=16'h59c4;
10786: douta=16'h61e4;
10787: douta=16'h6a04;
10788: douta=16'h7224;
10789: douta=16'h7204;
10790: douta=16'h7224;
10791: douta=16'h7203;
10792: douta=16'h7223;
10793: douta=16'h8ac6;
10794: douta=16'ha40a;
10795: douta=16'hc591;
10796: douta=16'hde95;
10797: douta=16'he6f6;
10798: douta=16'hde32;
10799: douta=16'hcd4e;
10800: douta=16'hbc27;
10801: douta=16'hb3a2;
10802: douta=16'hbb83;
10803: douta=16'hbbc4;
10804: douta=16'hc3e5;
10805: douta=16'hc405;
10806: douta=16'hc405;
10807: douta=16'hc425;
10808: douta=16'hcc25;
10809: douta=16'hcc26;
10810: douta=16'hcc26;
10811: douta=16'hcc46;
10812: douta=16'hcc45;
10813: douta=16'hcc45;
10814: douta=16'hcc45;
10815: douta=16'hd467;
10816: douta=16'hd466;
10817: douta=16'hcc46;
10818: douta=16'hcc66;
10819: douta=16'hd466;
10820: douta=16'hcc66;
10821: douta=16'hd466;
10822: douta=16'hd466;
10823: douta=16'hd466;
10824: douta=16'hd466;
10825: douta=16'hd466;
10826: douta=16'hd466;
10827: douta=16'hd466;
10828: douta=16'hd467;
10829: douta=16'hd488;
10830: douta=16'hdc84;
10831: douta=16'h8c52;
10832: douta=16'h8411;
10833: douta=16'h7b90;
10834: douta=16'h5a69;
10835: douta=16'h734b;
10836: douta=16'h940d;
10837: douta=16'hc552;
10838: douta=16'hde35;
10839: douta=16'hd635;
10840: douta=16'hbd33;
10841: douta=16'hcdd5;
10842: douta=16'hc595;
10843: douta=16'hacf5;
10844: douta=16'ha4f4;
10845: douta=16'h94b4;
10846: douta=16'h7c12;
10847: douta=16'h8c94;
10848: douta=16'h8c33;
10849: douta=16'h632f;
10850: douta=16'h8c32;
10851: douta=16'h73f1;
10852: douta=16'h6b4e;
10853: douta=16'h1060;
10854: douta=16'h7b2b;
10855: douta=16'hbd53;
10856: douta=16'h8c0d;
10857: douta=16'h5248;
10858: douta=16'hac8f;
10859: douta=16'hd5d4;
10860: douta=16'hc553;
10861: douta=16'ha470;
10862: douta=16'h62ed;
10863: douta=16'h31e9;
10864: douta=16'h18e5;
10865: douta=16'h420a;
10866: douta=16'h29a9;
10867: douta=16'h29a8;
10868: douta=16'h6a46;
10869: douta=16'h59e5;
10870: douta=16'h59e5;
10871: douta=16'h59e6;
10872: douta=16'h51c6;
10873: douta=16'h49a5;
10874: douta=16'h49a6;
10875: douta=16'h49a6;
10876: douta=16'h4186;
10877: douta=16'h4186;
10878: douta=16'h3965;
10879: douta=16'h3986;
10880: douta=16'hff9c;
10881: douta=16'hffbc;
10882: douta=16'hffdd;
10883: douta=16'hd5b3;
10884: douta=16'h9c73;
10885: douta=16'hb556;
10886: douta=16'hbd95;
10887: douta=16'hb555;
10888: douta=16'h8c74;
10889: douta=16'h8454;
10890: douta=16'h8475;
10891: douta=16'h7c34;
10892: douta=16'h7c55;
10893: douta=16'h8454;
10894: douta=16'h1020;
10895: douta=16'h18c3;
10896: douta=16'h1041;
10897: douta=16'h1861;
10898: douta=16'h1882;
10899: douta=16'h1883;
10900: douta=16'h1882;
10901: douta=16'h20a2;
10902: douta=16'h20a2;
10903: douta=16'h28c3;
10904: douta=16'h28e2;
10905: douta=16'h2904;
10906: douta=16'h18e5;
10907: douta=16'h3903;
10908: douta=16'h4143;
10909: douta=16'h4964;
10910: douta=16'h4984;
10911: douta=16'h5984;
10912: douta=16'h5163;
10913: douta=16'h5983;
10914: douta=16'h6a46;
10915: douta=16'h8329;
10916: douta=16'hacae;
10917: douta=16'hbd91;
10918: douta=16'hc5d1;
10919: douta=16'hb4ee;
10920: douta=16'ha40a;
10921: douta=16'h9306;
10922: douta=16'h8aa2;
10923: douta=16'h9282;
10924: douta=16'h9b04;
10925: douta=16'hab85;
10926: douta=16'hab85;
10927: douta=16'hb3a5;
10928: douta=16'hb3a4;
10929: douta=16'hc405;
10930: douta=16'hc405;
10931: douta=16'hc405;
10932: douta=16'hc425;
10933: douta=16'hc425;
10934: douta=16'hc445;
10935: douta=16'hc425;
10936: douta=16'hc425;
10937: douta=16'hcc25;
10938: douta=16'hcc26;
10939: douta=16'hcc26;
10940: douta=16'hcc45;
10941: douta=16'hcc46;
10942: douta=16'hcc46;
10943: douta=16'hcc46;
10944: douta=16'hcc47;
10945: douta=16'hcc66;
10946: douta=16'hcc66;
10947: douta=16'hcc66;
10948: douta=16'hd467;
10949: douta=16'hcc66;
10950: douta=16'hd467;
10951: douta=16'hd467;
10952: douta=16'hcc66;
10953: douta=16'hd466;
10954: douta=16'hd466;
10955: douta=16'hd467;
10956: douta=16'hd466;
10957: douta=16'hd467;
10958: douta=16'hcc66;
10959: douta=16'hd487;
10960: douta=16'h9c4f;
10961: douta=16'h9c4e;
10962: douta=16'hbd31;
10963: douta=16'hc573;
10964: douta=16'heeb7;
10965: douta=16'hde16;
10966: douta=16'hd615;
10967: douta=16'hcdd5;
10968: douta=16'hcdb5;
10969: douta=16'ha4d3;
10970: douta=16'h9cd5;
10971: douta=16'h9494;
10972: douta=16'h7bd1;
10973: douta=16'h7bf2;
10974: douta=16'h7bd1;
10975: douta=16'h73d1;
10976: douta=16'h73d1;
10977: douta=16'h4a28;
10978: douta=16'h3964;
10979: douta=16'h83cd;
10980: douta=16'h7bac;
10981: douta=16'hb4f1;
10982: douta=16'hb531;
10983: douta=16'h83ac;
10984: douta=16'h83ad;
10985: douta=16'hd5d4;
10986: douta=16'hcdb2;
10987: douta=16'h9c6f;
10988: douta=16'hb512;
10989: douta=16'hacd2;
10990: douta=16'h7bd1;
10991: douta=16'h4ace;
10992: douta=16'h3a0a;
10993: douta=16'h18e5;
10994: douta=16'h2968;
10995: douta=16'h1926;
10996: douta=16'h6a26;
10997: douta=16'h59e6;
10998: douta=16'h59e6;
10999: douta=16'h51c5;
11000: douta=16'h51c5;
11001: douta=16'h49a5;
11002: douta=16'h49a5;
11003: douta=16'h4986;
11004: douta=16'h4186;
11005: douta=16'h4186;
11006: douta=16'h4186;
11007: douta=16'h3986;
11008: douta=16'hff9c;
11009: douta=16'hff9c;
11010: douta=16'he6b8;
11011: douta=16'he657;
11012: douta=16'had36;
11013: douta=16'hb556;
11014: douta=16'hc596;
11015: douta=16'had55;
11016: douta=16'h8cb6;
11017: douta=16'h8475;
11018: douta=16'h8454;
11019: douta=16'h8495;
11020: douta=16'h8433;
11021: douta=16'h94f7;
11022: douta=16'h18a3;
11023: douta=16'h18a3;
11024: douta=16'h1061;
11025: douta=16'h18a2;
11026: douta=16'h1882;
11027: douta=16'h1882;
11028: douta=16'h20a2;
11029: douta=16'h20a2;
11030: douta=16'h2082;
11031: douta=16'h28c2;
11032: douta=16'h28c2;
11033: douta=16'h2925;
11034: douta=16'h18c4;
11035: douta=16'h49a5;
11036: douta=16'h62ca;
11037: douta=16'h8c2f;
11038: douta=16'h9490;
11039: douta=16'h8c2e;
11040: douta=16'h6a87;
11041: douta=16'h72a7;
11042: douta=16'h61e4;
11043: douta=16'h61a3;
11044: douta=16'h6a04;
11045: douta=16'h7203;
11046: douta=16'h7244;
11047: douta=16'h7a63;
11048: douta=16'h82a4;
11049: douta=16'h8ac4;
11050: douta=16'h92e5;
11051: douta=16'h9b25;
11052: douta=16'ha325;
11053: douta=16'hab64;
11054: douta=16'hab65;
11055: douta=16'hab84;
11056: douta=16'hbbc6;
11057: douta=16'hc406;
11058: douta=16'hc405;
11059: douta=16'hc426;
11060: douta=16'hc425;
11061: douta=16'hc425;
11062: douta=16'hc405;
11063: douta=16'hc425;
11064: douta=16'hcc26;
11065: douta=16'hcc26;
11066: douta=16'hcc25;
11067: douta=16'hcc46;
11068: douta=16'hcc46;
11069: douta=16'hcc46;
11070: douta=16'hcc46;
11071: douta=16'hcc46;
11072: douta=16'hcc46;
11073: douta=16'hd467;
11074: douta=16'hcc66;
11075: douta=16'hd467;
11076: douta=16'hd467;
11077: douta=16'hcc66;
11078: douta=16'hd466;
11079: douta=16'hd467;
11080: douta=16'hd467;
11081: douta=16'hd467;
11082: douta=16'hd467;
11083: douta=16'hd467;
11084: douta=16'hd467;
11085: douta=16'hd467;
11086: douta=16'hd467;
11087: douta=16'hd467;
11088: douta=16'hc448;
11089: douta=16'hacb1;
11090: douta=16'hd5d4;
11091: douta=16'hcdb4;
11092: douta=16'hc574;
11093: douta=16'hc555;
11094: douta=16'hc576;
11095: douta=16'hb536;
11096: douta=16'h9cf6;
11097: douta=16'h7c12;
11098: douta=16'h8432;
11099: douta=16'h73b0;
11100: douta=16'h7bd1;
11101: douta=16'h6b90;
11102: douta=16'h630e;
11103: douta=16'h41c6;
11104: douta=16'h732c;
11105: douta=16'h8bed;
11106: douta=16'hb530;
11107: douta=16'h9c4f;
11108: douta=16'hc531;
11109: douta=16'hbd51;
11110: douta=16'hb4f0;
11111: douta=16'hd635;
11112: douta=16'hde56;
11113: douta=16'hd5f4;
11114: douta=16'hd5b3;
11115: douta=16'hc553;
11116: douta=16'hacf3;
11117: douta=16'h9493;
11118: douta=16'h8412;
11119: douta=16'h5b4f;
11120: douta=16'h52ce;
11121: douta=16'h424c;
11122: douta=16'h5aac;
11123: douta=16'h18e5;
11124: douta=16'h2127;
11125: douta=16'h6205;
11126: douta=16'h59e6;
11127: douta=16'h51e5;
11128: douta=16'h51a5;
11129: douta=16'h49a5;
11130: douta=16'h49a6;
11131: douta=16'h49a6;
11132: douta=16'h49a6;
11133: douta=16'h4186;
11134: douta=16'h4186;
11135: douta=16'h3966;
11136: douta=16'hffdd;
11137: douta=16'hfffe;
11138: douta=16'he677;
11139: douta=16'hb555;
11140: douta=16'hbdb7;
11141: douta=16'hbd75;
11142: douta=16'hc595;
11143: douta=16'ha516;
11144: douta=16'h8c95;
11145: douta=16'h8c75;
11146: douta=16'h8454;
11147: douta=16'h8475;
11148: douta=16'h7c33;
11149: douta=16'h324b;
11150: douta=16'h1881;
11151: douta=16'h18a2;
11152: douta=16'h1062;
11153: douta=16'h1040;
11154: douta=16'h1061;
11155: douta=16'h20c3;
11156: douta=16'h2924;
11157: douta=16'h39a6;
11158: douta=16'h4a28;
11159: douta=16'h5269;
11160: douta=16'h4a27;
11161: douta=16'h2967;
11162: douta=16'h20e3;
11163: douta=16'h3902;
11164: douta=16'h4122;
11165: douta=16'h4963;
11166: douta=16'h51a4;
11167: douta=16'h6aea;
11168: douta=16'h3102;
11169: douta=16'h61e4;
11170: douta=16'h6a04;
11171: douta=16'h7224;
11172: douta=16'h7244;
11173: douta=16'h7244;
11174: douta=16'h7a44;
11175: douta=16'h7a63;
11176: douta=16'h8aa4;
11177: douta=16'h8ac5;
11178: douta=16'h9305;
11179: douta=16'h9b05;
11180: douta=16'h9b25;
11181: douta=16'hab65;
11182: douta=16'hab65;
11183: douta=16'hb3a5;
11184: douta=16'hb3c5;
11185: douta=16'hbbc5;
11186: douta=16'hbbe5;
11187: douta=16'hc405;
11188: douta=16'hbbe5;
11189: douta=16'hc405;
11190: douta=16'hc426;
11191: douta=16'hc405;
11192: douta=16'hc425;
11193: douta=16'hc425;
11194: douta=16'hcc26;
11195: douta=16'hcc26;
11196: douta=16'hcc46;
11197: douta=16'hcc46;
11198: douta=16'hcc46;
11199: douta=16'hcc46;
11200: douta=16'hcc66;
11201: douta=16'hd467;
11202: douta=16'hd467;
11203: douta=16'hd466;
11204: douta=16'hd467;
11205: douta=16'hd466;
11206: douta=16'hd466;
11207: douta=16'hd466;
11208: douta=16'hd467;
11209: douta=16'hd467;
11210: douta=16'hd467;
11211: douta=16'hd467;
11212: douta=16'hd467;
11213: douta=16'hd467;
11214: douta=16'hd467;
11215: douta=16'hd487;
11216: douta=16'hd466;
11217: douta=16'h942f;
11218: douta=16'ha492;
11219: douta=16'ha4d3;
11220: douta=16'hc575;
11221: douta=16'h94b5;
11222: douta=16'h8c74;
11223: douta=16'h7bf2;
11224: douta=16'h7bd1;
11225: douta=16'h6bb1;
11226: douta=16'h8432;
11227: douta=16'h5acb;
11228: douta=16'h39a6;
11229: douta=16'h5a8a;
11230: douta=16'h942e;
11231: douta=16'hb4d0;
11232: douta=16'hbd10;
11233: douta=16'hbd10;
11234: douta=16'hbd31;
11235: douta=16'hbd52;
11236: douta=16'hcdd4;
11237: douta=16'hd635;
11238: douta=16'hde15;
11239: douta=16'hde35;
11240: douta=16'hcdb4;
11241: douta=16'hc573;
11242: douta=16'hb514;
11243: douta=16'h9cb4;
11244: douta=16'h9cb4;
11245: douta=16'h8c93;
11246: douta=16'h8c74;
11247: douta=16'h6b6f;
11248: douta=16'h4acd;
11249: douta=16'h424b;
11250: douta=16'h2167;
11251: douta=16'h3189;
11252: douta=16'h1905;
11253: douta=16'h1905;
11254: douta=16'h59e6;
11255: douta=16'h51c5;
11256: douta=16'h51c5;
11257: douta=16'h49a6;
11258: douta=16'h49a6;
11259: douta=16'h49a6;
11260: douta=16'h41a6;
11261: douta=16'h4166;
11262: douta=16'h3966;
11263: douta=16'h3986;
11264: douta=16'hff9d;
11265: douta=16'hffbd;
11266: douta=16'heeb8;
11267: douta=16'ha4f4;
11268: douta=16'hbd96;
11269: douta=16'hc5b5;
11270: douta=16'hbd55;
11271: douta=16'h8c53;
11272: douta=16'h8454;
11273: douta=16'h8c75;
11274: douta=16'h8474;
11275: douta=16'h7bf3;
11276: douta=16'h94f7;
11277: douta=16'h18a3;
11278: douta=16'h18e3;
11279: douta=16'h29a8;
11280: douta=16'h2946;
11281: douta=16'h1904;
11282: douta=16'h20e3;
11283: douta=16'h2082;
11284: douta=16'h1881;
11285: douta=16'h2082;
11286: douta=16'h20c2;
11287: douta=16'h28e2;
11288: douta=16'h30e3;
11289: douta=16'h29a8;
11290: douta=16'h30e3;
11291: douta=16'h4143;
11292: douta=16'h4963;
11293: douta=16'h4964;
11294: douta=16'h51a4;
11295: douta=16'h83ef;
11296: douta=16'h59a3;
11297: douta=16'h69e4;
11298: douta=16'h7224;
11299: douta=16'h7224;
11300: douta=16'h7244;
11301: douta=16'h7244;
11302: douta=16'h7224;
11303: douta=16'h8285;
11304: douta=16'h8aa4;
11305: douta=16'h92e5;
11306: douta=16'h9305;
11307: douta=16'h9b05;
11308: douta=16'ha345;
11309: douta=16'hab64;
11310: douta=16'hb385;
11311: douta=16'hb3a5;
11312: douta=16'hb3c5;
11313: douta=16'hbbe6;
11314: douta=16'hbbc6;
11315: douta=16'hbbe5;
11316: douta=16'hc405;
11317: douta=16'hc406;
11318: douta=16'hc406;
11319: douta=16'hc425;
11320: douta=16'hc425;
11321: douta=16'hc425;
11322: douta=16'hcc26;
11323: douta=16'hcc46;
11324: douta=16'hcc46;
11325: douta=16'hcc46;
11326: douta=16'hd467;
11327: douta=16'hd467;
11328: douta=16'hcc46;
11329: douta=16'hd467;
11330: douta=16'hcc46;
11331: douta=16'hd467;
11332: douta=16'hd467;
11333: douta=16'hd467;
11334: douta=16'hd466;
11335: douta=16'hd467;
11336: douta=16'hd467;
11337: douta=16'hd467;
11338: douta=16'hd467;
11339: douta=16'hd467;
11340: douta=16'hd467;
11341: douta=16'hd467;
11342: douta=16'hd487;
11343: douta=16'hd487;
11344: douta=16'hcc87;
11345: douta=16'hcd6f;
11346: douta=16'hacd3;
11347: douta=16'h9452;
11348: douta=16'h9473;
11349: douta=16'h83f1;
11350: douta=16'h7bd0;
11351: douta=16'h6b4f;
11352: douta=16'h6b4f;
11353: douta=16'h5acd;
11354: douta=16'h5a68;
11355: douta=16'h8bcd;
11356: douta=16'ha4b0;
11357: douta=16'hc573;
11358: douta=16'hc572;
11359: douta=16'hc573;
11360: douta=16'hddf4;
11361: douta=16'hd5d3;
11362: douta=16'hde35;
11363: douta=16'hc5b4;
11364: douta=16'hc594;
11365: douta=16'hcdf4;
11366: douta=16'hc5b4;
11367: douta=16'hcdb4;
11368: douta=16'hc574;
11369: douta=16'hb514;
11370: douta=16'ha4f4;
11371: douta=16'h94b4;
11372: douta=16'h8c93;
11373: douta=16'h8412;
11374: douta=16'h73b1;
11375: douta=16'h73d1;
11376: douta=16'h6b90;
11377: douta=16'h632d;
11378: douta=16'h18a3;
11379: douta=16'h732e;
11380: douta=16'h29c9;
11381: douta=16'h18e5;
11382: douta=16'h61e6;
11383: douta=16'h59e6;
11384: douta=16'h51c6;
11385: douta=16'h49a6;
11386: douta=16'h49a5;
11387: douta=16'h4185;
11388: douta=16'h4185;
11389: douta=16'h4186;
11390: douta=16'h3966;
11391: douta=16'h3966;
11392: douta=16'hffbd;
11393: douta=16'hde77;
11394: douta=16'he697;
11395: douta=16'ha4b4;
11396: douta=16'hb535;
11397: douta=16'hc595;
11398: douta=16'hbd76;
11399: douta=16'h8c74;
11400: douta=16'h8c74;
11401: douta=16'h8454;
11402: douta=16'h73f3;
11403: douta=16'h8454;
11404: douta=16'h2145;
11405: douta=16'h18c3;
11406: douta=16'h18a3;
11407: douta=16'h1082;
11408: douta=16'h1882;
11409: douta=16'h1882;
11410: douta=16'h1881;
11411: douta=16'h20a2;
11412: douta=16'h20a2;
11413: douta=16'h20a2;
11414: douta=16'h20c2;
11415: douta=16'h28e2;
11416: douta=16'h30e2;
11417: douta=16'h2988;
11418: douta=16'h4123;
11419: douta=16'h4143;
11420: douta=16'h4963;
11421: douta=16'h51a4;
11422: douta=16'h59a4;
11423: douta=16'h9d13;
11424: douta=16'h6a04;
11425: douta=16'h7224;
11426: douta=16'h7224;
11427: douta=16'h7244;
11428: douta=16'h7244;
11429: douta=16'h7224;
11430: douta=16'h7a44;
11431: douta=16'h8284;
11432: douta=16'h8ac5;
11433: douta=16'h92c4;
11434: douta=16'h9304;
11435: douta=16'ha325;
11436: douta=16'ha345;
11437: douta=16'hab85;
11438: douta=16'hb385;
11439: douta=16'hb385;
11440: douta=16'hb3c5;
11441: douta=16'hbbe5;
11442: douta=16'hbbe5;
11443: douta=16'hbc06;
11444: douta=16'hc406;
11445: douta=16'hc426;
11446: douta=16'hc426;
11447: douta=16'hc425;
11448: douta=16'hc425;
11449: douta=16'hc425;
11450: douta=16'hcc46;
11451: douta=16'hcc46;
11452: douta=16'hcc46;
11453: douta=16'hcc47;
11454: douta=16'hd467;
11455: douta=16'hd466;
11456: douta=16'hcc46;
11457: douta=16'hd467;
11458: douta=16'hcc66;
11459: douta=16'hd467;
11460: douta=16'hd467;
11461: douta=16'hd466;
11462: douta=16'hd467;
11463: douta=16'hd467;
11464: douta=16'hd488;
11465: douta=16'hd467;
11466: douta=16'hd467;
11467: douta=16'hd467;
11468: douta=16'hd468;
11469: douta=16'hd467;
11470: douta=16'hd467;
11471: douta=16'hd487;
11472: douta=16'hd487;
11473: douta=16'hbccd;
11474: douta=16'hb44b;
11475: douta=16'h9410;
11476: douta=16'h83b0;
11477: douta=16'h734e;
11478: douta=16'h62cd;
11479: douta=16'h49e6;
11480: douta=16'h5a8a;
11481: douta=16'hd614;
11482: douta=16'h8bed;
11483: douta=16'hbd30;
11484: douta=16'hcdb4;
11485: douta=16'hbd52;
11486: douta=16'hde35;
11487: douta=16'he676;
11488: douta=16'hde15;
11489: douta=16'hde35;
11490: douta=16'hd615;
11491: douta=16'ha4d3;
11492: douta=16'hc595;
11493: douta=16'hb534;
11494: douta=16'hacf4;
11495: douta=16'hb514;
11496: douta=16'h9cb4;
11497: douta=16'h8432;
11498: douta=16'h7bb1;
11499: douta=16'h73b1;
11500: douta=16'h736f;
11501: douta=16'h5a69;
11502: douta=16'h2903;
11503: douta=16'h62ca;
11504: douta=16'h5269;
11505: douta=16'h5b50;
11506: douta=16'h4aef;
11507: douta=16'h736f;
11508: douta=16'h1083;
11509: douta=16'h2126;
11510: douta=16'h4186;
11511: douta=16'h51e6;
11512: douta=16'h49c5;
11513: douta=16'h49a6;
11514: douta=16'h4186;
11515: douta=16'h4186;
11516: douta=16'h4185;
11517: douta=16'h3966;
11518: douta=16'h4166;
11519: douta=16'h4166;
11520: douta=16'hffdd;
11521: douta=16'hde16;
11522: douta=16'hd5f6;
11523: douta=16'h9c93;
11524: douta=16'hc595;
11525: douta=16'hbd55;
11526: douta=16'h9cd5;
11527: douta=16'h94b5;
11528: douta=16'h8c74;
11529: douta=16'h8454;
11530: douta=16'h8454;
11531: douta=16'h94f7;
11532: douta=16'h1861;
11533: douta=16'h20c2;
11534: douta=16'h18a3;
11535: douta=16'h1082;
11536: douta=16'h1882;
11537: douta=16'h1882;
11538: douta=16'h2082;
11539: douta=16'h1881;
11540: douta=16'h20a2;
11541: douta=16'h20a2;
11542: douta=16'h28c2;
11543: douta=16'h28e2;
11544: douta=16'h3103;
11545: douta=16'h2126;
11546: douta=16'h4163;
11547: douta=16'h4163;
11548: douta=16'h4984;
11549: douta=16'h51a4;
11550: douta=16'h5163;
11551: douta=16'h9cd1;
11552: douta=16'h6204;
11553: douta=16'h61c4;
11554: douta=16'h7224;
11555: douta=16'h7244;
11556: douta=16'h7a65;
11557: douta=16'h7244;
11558: douta=16'h7a64;
11559: douta=16'h82a4;
11560: douta=16'h8ac4;
11561: douta=16'h9304;
11562: douta=16'h9305;
11563: douta=16'h9b25;
11564: douta=16'ha345;
11565: douta=16'hab85;
11566: douta=16'hb385;
11567: douta=16'hb3a5;
11568: douta=16'hbbc5;
11569: douta=16'hbbe6;
11570: douta=16'hbbe5;
11571: douta=16'hbc06;
11572: douta=16'hc406;
11573: douta=16'hc405;
11574: douta=16'hcc26;
11575: douta=16'hc425;
11576: douta=16'hc425;
11577: douta=16'hc425;
11578: douta=16'hcc26;
11579: douta=16'hcc46;
11580: douta=16'hcc47;
11581: douta=16'hcc46;
11582: douta=16'hcc46;
11583: douta=16'hcc67;
11584: douta=16'hd467;
11585: douta=16'hd467;
11586: douta=16'hd467;
11587: douta=16'hd467;
11588: douta=16'hcc47;
11589: douta=16'hd467;
11590: douta=16'hd467;
11591: douta=16'hd468;
11592: douta=16'hd467;
11593: douta=16'hd487;
11594: douta=16'hd467;
11595: douta=16'hd467;
11596: douta=16'hd467;
11597: douta=16'hd467;
11598: douta=16'hd487;
11599: douta=16'hd468;
11600: douta=16'hd467;
11601: douta=16'hb4cd;
11602: douta=16'hcc46;
11603: douta=16'ha44e;
11604: douta=16'h62ec;
11605: douta=16'h4a28;
11606: douta=16'h9c4f;
11607: douta=16'ha490;
11608: douta=16'hd614;
11609: douta=16'h8bee;
11610: douta=16'hd5f3;
11611: douta=16'hd5d3;
11612: douta=16'hd5d4;
11613: douta=16'he677;
11614: douta=16'hd5d4;
11615: douta=16'hbd74;
11616: douta=16'hc574;
11617: douta=16'hb554;
11618: douta=16'ha4d4;
11619: douta=16'had14;
11620: douta=16'h9cd5;
11621: douta=16'h8c53;
11622: douta=16'h8432;
11623: douta=16'h8c33;
11624: douta=16'h7bf1;
11625: douta=16'h7bf1;
11626: douta=16'h5248;
11627: douta=16'h3944;
11628: douta=16'h5a88;
11629: douta=16'h5a89;
11630: douta=16'h734b;
11631: douta=16'h83ad;
11632: douta=16'h524a;
11633: douta=16'h2126;
11634: douta=16'h2146;
11635: douta=16'h5249;
11636: douta=16'h3a2b;
11637: douta=16'h18e5;
11638: douta=16'h5a06;
11639: douta=16'h51c6;
11640: douta=16'h49c6;
11641: douta=16'h49a6;
11642: douta=16'h49a6;
11643: douta=16'h4186;
11644: douta=16'h4185;
11645: douta=16'h4185;
11646: douta=16'h4166;
11647: douta=16'h4166;
11648: douta=16'hffbc;
11649: douta=16'he698;
11650: douta=16'ha4f4;
11651: douta=16'had15;
11652: douta=16'hcdb5;
11653: douta=16'hbd55;
11654: douta=16'h8c53;
11655: douta=16'h9494;
11656: douta=16'h8c74;
11657: douta=16'h8434;
11658: douta=16'h8454;
11659: douta=16'h73f2;
11660: douta=16'h20e3;
11661: douta=16'h20c3;
11662: douta=16'h20e3;
11663: douta=16'h1882;
11664: douta=16'h1882;
11665: douta=16'h18a2;
11666: douta=16'h1881;
11667: douta=16'h20a2;
11668: douta=16'h20a2;
11669: douta=16'h20c2;
11670: douta=16'h28e2;
11671: douta=16'h28e2;
11672: douta=16'h3146;
11673: douta=16'h18e5;
11674: douta=16'h4143;
11675: douta=16'h4963;
11676: douta=16'h5184;
11677: douta=16'h59a4;
11678: douta=16'h5183;
11679: douta=16'h8bec;
11680: douta=16'h6204;
11681: douta=16'h59a4;
11682: douta=16'h7224;
11683: douta=16'h7a64;
11684: douta=16'h7a44;
11685: douta=16'h7a44;
11686: douta=16'h7a64;
11687: douta=16'h82a5;
11688: douta=16'h8ac4;
11689: douta=16'h9304;
11690: douta=16'h9b05;
11691: douta=16'ha325;
11692: douta=16'ha365;
11693: douta=16'hab85;
11694: douta=16'hb3a5;
11695: douta=16'hb3a6;
11696: douta=16'hbbe6;
11697: douta=16'hbbe6;
11698: douta=16'hc406;
11699: douta=16'hbc06;
11700: douta=16'hc406;
11701: douta=16'hc406;
11702: douta=16'hc426;
11703: douta=16'hcc47;
11704: douta=16'hc426;
11705: douta=16'hcc46;
11706: douta=16'hcc46;
11707: douta=16'hcc47;
11708: douta=16'hcc46;
11709: douta=16'hcc46;
11710: douta=16'hcc46;
11711: douta=16'hcc46;
11712: douta=16'hcc47;
11713: douta=16'hd467;
11714: douta=16'hd467;
11715: douta=16'hcc67;
11716: douta=16'hd467;
11717: douta=16'hd467;
11718: douta=16'hd467;
11719: douta=16'hd467;
11720: douta=16'hd467;
11721: douta=16'hd467;
11722: douta=16'hd467;
11723: douta=16'hd487;
11724: douta=16'hd467;
11725: douta=16'hd467;
11726: douta=16'hd487;
11727: douta=16'hd487;
11728: douta=16'hd467;
11729: douta=16'hbcce;
11730: douta=16'hcc46;
11731: douta=16'hd486;
11732: douta=16'h940f;
11733: douta=16'h9c2e;
11734: douta=16'hc571;
11735: douta=16'hbd73;
11736: douta=16'hcdd5;
11737: douta=16'hcdd6;
11738: douta=16'hde56;
11739: douta=16'hd5f4;
11740: douta=16'hd5d3;
11741: douta=16'hbd33;
11742: douta=16'hb513;
11743: douta=16'hb513;
11744: douta=16'hacf4;
11745: douta=16'h9cb4;
11746: douta=16'h9cb4;
11747: douta=16'h8c73;
11748: douta=16'h7c32;
11749: douta=16'h7bb0;
11750: douta=16'h7b8f;
11751: douta=16'h51e6;
11752: douta=16'h41a5;
11753: douta=16'h5226;
11754: douta=16'h732c;
11755: douta=16'h62c9;
11756: douta=16'h6b0a;
11757: douta=16'h83cd;
11758: douta=16'h942e;
11759: douta=16'h9c4f;
11760: douta=16'h7b8e;
11761: douta=16'h2967;
11762: douta=16'h10e3;
11763: douta=16'h0883;
11764: douta=16'h0042;
11765: douta=16'h2126;
11766: douta=16'h5249;
11767: douta=16'h51c6;
11768: douta=16'h49a6;
11769: douta=16'h4986;
11770: douta=16'h49a6;
11771: douta=16'h4185;
11772: douta=16'h4185;
11773: douta=16'h4186;
11774: douta=16'h4186;
11775: douta=16'h4186;
11776: douta=16'hd5d5;
11777: douta=16'he677;
11778: douta=16'ha4b3;
11779: douta=16'hb556;
11780: douta=16'hc595;
11781: douta=16'hb556;
11782: douta=16'h9494;
11783: douta=16'h94b5;
11784: douta=16'h8c74;
11785: douta=16'h8454;
11786: douta=16'h8454;
11787: douta=16'h1020;
11788: douta=16'h20c3;
11789: douta=16'h20a3;
11790: douta=16'h20e3;
11791: douta=16'h1882;
11792: douta=16'h1882;
11793: douta=16'h20a2;
11794: douta=16'h1881;
11795: douta=16'h20a2;
11796: douta=16'h20a2;
11797: douta=16'h28e2;
11798: douta=16'h28e2;
11799: douta=16'h30e2;
11800: douta=16'h39a8;
11801: douta=16'h18c5;
11802: douta=16'h4143;
11803: douta=16'h4963;
11804: douta=16'h5184;
11805: douta=16'h59c4;
11806: douta=16'h6206;
11807: douta=16'h72a7;
11808: douta=16'h6a24;
11809: douta=16'h59a4;
11810: douta=16'h7244;
11811: douta=16'h7a64;
11812: douta=16'h7a64;
11813: douta=16'h7a44;
11814: douta=16'h7a84;
11815: douta=16'h82a4;
11816: douta=16'h8ae5;
11817: douta=16'h9304;
11818: douta=16'h9b05;
11819: douta=16'ha345;
11820: douta=16'hab65;
11821: douta=16'hb385;
11822: douta=16'hb3a5;
11823: douta=16'hbbc6;
11824: douta=16'hbbe6;
11825: douta=16'hbbe6;
11826: douta=16'hc406;
11827: douta=16'hc406;
11828: douta=16'hc406;
11829: douta=16'hc426;
11830: douta=16'hc426;
11831: douta=16'hc426;
11832: douta=16'hcc26;
11833: douta=16'hcc47;
11834: douta=16'hcc47;
11835: douta=16'hcc47;
11836: douta=16'hcc46;
11837: douta=16'hcc46;
11838: douta=16'hcc46;
11839: douta=16'hcc46;
11840: douta=16'hd467;
11841: douta=16'hcc47;
11842: douta=16'hcc67;
11843: douta=16'hd467;
11844: douta=16'hd467;
11845: douta=16'hd467;
11846: douta=16'hd467;
11847: douta=16'hd467;
11848: douta=16'hd467;
11849: douta=16'hd467;
11850: douta=16'hd467;
11851: douta=16'hd467;
11852: douta=16'hd487;
11853: douta=16'hd467;
11854: douta=16'hd487;
11855: douta=16'hd468;
11856: douta=16'hd488;
11857: douta=16'hb4ce;
11858: douta=16'hcc45;
11859: douta=16'hd487;
11860: douta=16'habec;
11861: douta=16'hacd0;
11862: douta=16'hcdd4;
11863: douta=16'hd615;
11864: douta=16'hb513;
11865: douta=16'hde36;
11866: douta=16'hcdb5;
11867: douta=16'hacf3;
11868: douta=16'ha4b2;
11869: douta=16'h9c93;
11870: douta=16'h9c94;
11871: douta=16'h8c11;
11872: douta=16'h9452;
11873: douta=16'h8412;
11874: douta=16'h7390;
11875: douta=16'h62aa;
11876: douta=16'h3944;
11877: douta=16'h41a5;
11878: douta=16'h6ac9;
11879: douta=16'h5a88;
11880: douta=16'h732a;
11881: douta=16'h7b8c;
11882: douta=16'h9c6f;
11883: douta=16'hacf0;
11884: douta=16'hb4f0;
11885: douta=16'hb511;
11886: douta=16'hb511;
11887: douta=16'hacd1;
11888: douta=16'h8c30;
11889: douta=16'h6b6f;
11890: douta=16'h424b;
11891: douta=16'h2967;
11892: douta=16'h31c9;
11893: douta=16'h2988;
11894: douta=16'h0863;
11895: douta=16'h51a5;
11896: douta=16'h4965;
11897: douta=16'h4124;
11898: douta=16'h4165;
11899: douta=16'h5208;
11900: douta=16'h630c;
11901: douta=16'h73d1;
11902: douta=16'h84b5;
11903: douta=16'h84b4;
11904: douta=16'hcdb5;
11905: douta=16'hde37;
11906: douta=16'ha4d3;
11907: douta=16'hb514;
11908: douta=16'hb535;
11909: douta=16'h9494;
11910: douta=16'h9474;
11911: douta=16'h94b5;
11912: douta=16'h8c74;
11913: douta=16'h8c95;
11914: douta=16'h9d38;
11915: douta=16'h20c3;
11916: douta=16'h20c3;
11917: douta=16'h20c3;
11918: douta=16'h18c3;
11919: douta=16'h1882;
11920: douta=16'h1882;
11921: douta=16'h2082;
11922: douta=16'h20a2;
11923: douta=16'h2082;
11924: douta=16'h20c2;
11925: douta=16'h28e2;
11926: douta=16'h28c2;
11927: douta=16'h30e3;
11928: douta=16'h39e9;
11929: douta=16'h28e4;
11930: douta=16'h4143;
11931: douta=16'h4963;
11932: douta=16'h5184;
11933: douta=16'h59a4;
11934: douta=16'h6b0a;
11935: douta=16'h61a3;
11936: douta=16'h6a24;
11937: douta=16'h51a4;
11938: douta=16'h7a64;
11939: douta=16'h7a64;
11940: douta=16'h7a44;
11941: douta=16'h7a84;
11942: douta=16'h8284;
11943: douta=16'h8ac5;
11944: douta=16'h8ae4;
11945: douta=16'h9305;
11946: douta=16'h9b26;
11947: douta=16'ha345;
11948: douta=16'hab65;
11949: douta=16'hb3a5;
11950: douta=16'hb3a5;
11951: douta=16'hbbc5;
11952: douta=16'hbbe6;
11953: douta=16'hbbe6;
11954: douta=16'hc406;
11955: douta=16'hc406;
11956: douta=16'hc426;
11957: douta=16'hc426;
11958: douta=16'hc426;
11959: douta=16'hcc26;
11960: douta=16'hc426;
11961: douta=16'hcc46;
11962: douta=16'hcc46;
11963: douta=16'hcc46;
11964: douta=16'hcc46;
11965: douta=16'hcc46;
11966: douta=16'hcc67;
11967: douta=16'hcc47;
11968: douta=16'hcc67;
11969: douta=16'hcc46;
11970: douta=16'hd467;
11971: douta=16'hd467;
11972: douta=16'hd467;
11973: douta=16'hcc67;
11974: douta=16'hd467;
11975: douta=16'hd468;
11976: douta=16'hd487;
11977: douta=16'hd467;
11978: douta=16'hd487;
11979: douta=16'hd467;
11980: douta=16'hd467;
11981: douta=16'hd487;
11982: douta=16'hd467;
11983: douta=16'hd488;
11984: douta=16'hd487;
11985: douta=16'hb4ce;
11986: douta=16'hcc45;
11987: douta=16'hd487;
11988: douta=16'hcc87;
11989: douta=16'ha4b1;
11990: douta=16'hc553;
11991: douta=16'hcdf5;
11992: douta=16'hbd54;
11993: douta=16'hbd96;
11994: douta=16'hb556;
11995: douta=16'h9493;
11996: douta=16'h8411;
11997: douta=16'h83f1;
11998: douta=16'h7bb0;
11999: douta=16'h83f0;
12000: douta=16'h5248;
12001: douta=16'h2903;
12002: douta=16'h6aea;
12003: douta=16'h62ca;
12004: douta=16'h732a;
12005: douta=16'h730a;
12006: douta=16'h8bcc;
12007: douta=16'h8c0e;
12008: douta=16'h944f;
12009: douta=16'h9c6f;
12010: douta=16'hb510;
12011: douta=16'hc572;
12012: douta=16'hcd92;
12013: douta=16'hd5d4;
12014: douta=16'hcd93;
12015: douta=16'hacd2;
12016: douta=16'h8c10;
12017: douta=16'h632e;
12018: douta=16'h52cd;
12019: douta=16'h426c;
12020: douta=16'h2106;
12021: douta=16'h1905;
12022: douta=16'h2127;
12023: douta=16'h10e5;
12024: douta=16'h8471;
12025: douta=16'h632c;
12026: douta=16'h52aa;
12027: douta=16'h5228;
12028: douta=16'h49c6;
12029: douta=16'h4985;
12030: douta=16'h4985;
12031: douta=16'h5185;
12032: douta=16'hde37;
12033: douta=16'had14;
12034: douta=16'hacf4;
12035: douta=16'hd5f6;
12036: douta=16'hb555;
12037: douta=16'h9c73;
12038: douta=16'h94b5;
12039: douta=16'h94b5;
12040: douta=16'h8454;
12041: douta=16'h8c95;
12042: douta=16'h2124;
12043: douta=16'h20a3;
12044: douta=16'h20c3;
12045: douta=16'h20c3;
12046: douta=16'h1882;
12047: douta=16'h1882;
12048: douta=16'h1861;
12049: douta=16'h20a2;
12050: douta=16'h20a2;
12051: douta=16'h20a2;
12052: douta=16'h20c2;
12053: douta=16'h28e2;
12054: douta=16'h30e2;
12055: douta=16'h3103;
12056: douta=16'h31a8;
12057: douta=16'h3944;
12058: douta=16'h4963;
12059: douta=16'h4984;
12060: douta=16'h5184;
12061: douta=16'h61c4;
12062: douta=16'h8c50;
12063: douta=16'h69e3;
12064: douta=16'h6a24;
12065: douta=16'h4164;
12066: douta=16'h7244;
12067: douta=16'h7a84;
12068: douta=16'h7a64;
12069: douta=16'h7a64;
12070: douta=16'h8285;
12071: douta=16'h8aa4;
12072: douta=16'h8ae4;
12073: douta=16'h9b25;
12074: douta=16'ha346;
12075: douta=16'ha345;
12076: douta=16'hab85;
12077: douta=16'hb3a5;
12078: douta=16'hb3a6;
12079: douta=16'hbbc5;
12080: douta=16'hbbe6;
12081: douta=16'hbbe6;
12082: douta=16'hc406;
12083: douta=16'hc406;
12084: douta=16'hc405;
12085: douta=16'hc426;
12086: douta=16'hc426;
12087: douta=16'hc426;
12088: douta=16'hcc26;
12089: douta=16'hcc47;
12090: douta=16'hcc46;
12091: douta=16'hcc45;
12092: douta=16'hcc46;
12093: douta=16'hcc47;
12094: douta=16'hcc47;
12095: douta=16'hcc67;
12096: douta=16'hcc47;
12097: douta=16'hd467;
12098: douta=16'hd467;
12099: douta=16'hd467;
12100: douta=16'hd467;
12101: douta=16'hcc67;
12102: douta=16'hd467;
12103: douta=16'hd468;
12104: douta=16'hd467;
12105: douta=16'hd467;
12106: douta=16'hd467;
12107: douta=16'hd467;
12108: douta=16'hd488;
12109: douta=16'hd488;
12110: douta=16'hd488;
12111: douta=16'hd467;
12112: douta=16'hd488;
12113: douta=16'hb4ee;
12114: douta=16'hcc25;
12115: douta=16'hd488;
12116: douta=16'hd487;
12117: douta=16'h9430;
12118: douta=16'h9c92;
12119: douta=16'had15;
12120: douta=16'hb515;
12121: douta=16'h9493;
12122: douta=16'h8c53;
12123: douta=16'h73b0;
12124: douta=16'h736f;
12125: douta=16'h6acc;
12126: douta=16'h3964;
12127: douta=16'h62a9;
12128: douta=16'h62c9;
12129: douta=16'h6b2a;
12130: douta=16'h5a68;
12131: douta=16'ha4b0;
12132: douta=16'h940e;
12133: douta=16'h93ed;
12134: douta=16'h9c4e;
12135: douta=16'hb4f0;
12136: douta=16'hc551;
12137: douta=16'hcd93;
12138: douta=16'hd5f4;
12139: douta=16'hd5d4;
12140: douta=16'hd5f4;
12141: douta=16'hcdd4;
12142: douta=16'hcd93;
12143: douta=16'hbd53;
12144: douta=16'h9c51;
12145: douta=16'h83f0;
12146: douta=16'h52ed;
12147: douta=16'h52ee;
12148: douta=16'h31c9;
12149: douta=16'h10c3;
12150: douta=16'h2126;
12151: douta=16'h08a4;
12152: douta=16'h2904;
12153: douta=16'h51a6;
12154: douta=16'h49a5;
12155: douta=16'h49a5;
12156: douta=16'h51c6;
12157: douta=16'h51c6;
12158: douta=16'h59c6;
12159: douta=16'h51c5;
12160: douta=16'he698;
12161: douta=16'hb535;
12162: douta=16'had15;
12163: douta=16'hc595;
12164: douta=16'ha536;
12165: douta=16'h9474;
12166: douta=16'h9494;
12167: douta=16'h9495;
12168: douta=16'h8433;
12169: douta=16'h9d59;
12170: douta=16'h20a3;
12171: douta=16'h20a3;
12172: douta=16'h20c3;
12173: douta=16'h20c3;
12174: douta=16'h18a2;
12175: douta=16'h20a2;
12176: douta=16'h20a2;
12177: douta=16'h20a2;
12178: douta=16'h20a2;
12179: douta=16'h20c2;
12180: douta=16'h28c2;
12181: douta=16'h28e3;
12182: douta=16'h3103;
12183: douta=16'h3103;
12184: douta=16'h2967;
12185: douta=16'h4963;
12186: douta=16'h4984;
12187: douta=16'h5184;
12188: douta=16'h59a4;
12189: douta=16'h61e4;
12190: douta=16'ha573;
12191: douta=16'h6a24;
12192: douta=16'h7224;
12193: douta=16'h6204;
12194: douta=16'h7a64;
12195: douta=16'h7a84;
12196: douta=16'h7a84;
12197: douta=16'h8285;
12198: douta=16'h82a4;
12199: douta=16'h8ac4;
12200: douta=16'h8ac4;
12201: douta=16'h9325;
12202: douta=16'ha325;
12203: douta=16'ha345;
12204: douta=16'hab85;
12205: douta=16'hb3a6;
12206: douta=16'hb3a6;
12207: douta=16'hbbc6;
12208: douta=16'hbc06;
12209: douta=16'hbbe5;
12210: douta=16'hc406;
12211: douta=16'hc405;
12212: douta=16'hc426;
12213: douta=16'hc426;
12214: douta=16'hc426;
12215: douta=16'hcc46;
12216: douta=16'hcc26;
12217: douta=16'hcc46;
12218: douta=16'hcc47;
12219: douta=16'hcc47;
12220: douta=16'hcc46;
12221: douta=16'hcc46;
12222: douta=16'hcc47;
12223: douta=16'hcc67;
12224: douta=16'hcc46;
12225: douta=16'hd467;
12226: douta=16'hd467;
12227: douta=16'hd467;
12228: douta=16'hcc67;
12229: douta=16'hd467;
12230: douta=16'hd468;
12231: douta=16'hd487;
12232: douta=16'hd467;
12233: douta=16'hd467;
12234: douta=16'hd467;
12235: douta=16'hd467;
12236: douta=16'hd487;
12237: douta=16'hd487;
12238: douta=16'hd488;
12239: douta=16'hd488;
12240: douta=16'hcc68;
12241: douta=16'haccd;
12242: douta=16'hcc25;
12243: douta=16'hcc68;
12244: douta=16'hcc88;
12245: douta=16'hc468;
12246: douta=16'h9431;
12247: douta=16'h83f1;
12248: douta=16'h7bb0;
12249: douta=16'h738f;
12250: douta=16'h9432;
12251: douta=16'h49e6;
12252: douta=16'h39a4;
12253: douta=16'h5a68;
12254: douta=16'h7b8d;
12255: douta=16'h6b0a;
12256: douta=16'h838c;
12257: douta=16'h83cd;
12258: douta=16'ha470;
12259: douta=16'h942f;
12260: douta=16'hbd10;
12261: douta=16'hb4f0;
12262: douta=16'hc552;
12263: douta=16'hd5d3;
12264: douta=16'hcdb3;
12265: douta=16'hd615;
12266: douta=16'hd5f4;
12267: douta=16'hd5b3;
12268: douta=16'hc533;
12269: douta=16'hb4f3;
12270: douta=16'hacd3;
12271: douta=16'ha4b3;
12272: douta=16'hacf4;
12273: douta=16'h8c93;
12274: douta=16'h7412;
12275: douta=16'h422a;
12276: douta=16'h1927;
12277: douta=16'h1927;
12278: douta=16'h08a3;
12279: douta=16'h18c5;
12280: douta=16'h08c6;
12281: douta=16'h59e6;
12282: douta=16'h51c5;
12283: douta=16'h59e6;
12284: douta=16'h51c6;
12285: douta=16'h59e6;
12286: douta=16'h59e6;
12287: douta=16'h59e6;
12288: douta=16'hcdb5;
12289: douta=16'hb534;
12290: douta=16'hcdd5;
12291: douta=16'hbd55;
12292: douta=16'h9453;
12293: douta=16'h9cb4;
12294: douta=16'h94d5;
12295: douta=16'h8c74;
12296: douta=16'h8454;
12297: douta=16'h2945;
12298: douta=16'h20c3;
12299: douta=16'h20a3;
12300: douta=16'h20c3;
12301: douta=16'h20a2;
12302: douta=16'h18a1;
12303: douta=16'h1881;
12304: douta=16'h20a2;
12305: douta=16'h20a2;
12306: douta=16'h20a2;
12307: douta=16'h20c2;
12308: douta=16'h28e2;
12309: douta=16'h30e3;
12310: douta=16'h30e3;
12311: douta=16'h3903;
12312: douta=16'h1906;
12313: douta=16'h4963;
12314: douta=16'h4983;
12315: douta=16'h51a4;
12316: douta=16'h59a4;
12317: douta=16'h59c3;
12318: douta=16'ha4f2;
12319: douta=16'h6a24;
12320: douta=16'h7244;
12321: douta=16'h8285;
12322: douta=16'h7a64;
12323: douta=16'h8284;
12324: douta=16'h7a64;
12325: douta=16'h7a64;
12326: douta=16'h82a4;
12327: douta=16'h8aa4;
12328: douta=16'h92c4;
12329: douta=16'h9b26;
12330: douta=16'ha346;
12331: douta=16'ha365;
12332: douta=16'hab85;
12333: douta=16'hb3a5;
12334: douta=16'hb3a6;
12335: douta=16'hbbc6;
12336: douta=16'hbbe6;
12337: douta=16'hbbe5;
12338: douta=16'hc406;
12339: douta=16'hc406;
12340: douta=16'hc405;
12341: douta=16'hc426;
12342: douta=16'hc426;
12343: douta=16'hc446;
12344: douta=16'hc446;
12345: douta=16'hc446;
12346: douta=16'hcc47;
12347: douta=16'hcc47;
12348: douta=16'hcc47;
12349: douta=16'hcc47;
12350: douta=16'hcc67;
12351: douta=16'hcc67;
12352: douta=16'hcc46;
12353: douta=16'hcc67;
12354: douta=16'hcc67;
12355: douta=16'hd468;
12356: douta=16'hd468;
12357: douta=16'hd468;
12358: douta=16'hd467;
12359: douta=16'hd487;
12360: douta=16'hd467;
12361: douta=16'hd487;
12362: douta=16'hd487;
12363: douta=16'hd488;
12364: douta=16'hd488;
12365: douta=16'hd488;
12366: douta=16'hd488;
12367: douta=16'hd488;
12368: douta=16'hd488;
12369: douta=16'hacce;
12370: douta=16'hcc03;
12371: douta=16'hcc46;
12372: douta=16'hcc04;
12373: douta=16'hc426;
12374: douta=16'h8c30;
12375: douta=16'h7b8f;
12376: douta=16'h5a48;
12377: douta=16'h4a06;
12378: douta=16'h732a;
12379: douta=16'h6b0b;
12380: douta=16'h734b;
12381: douta=16'h8bed;
12382: douta=16'hb511;
12383: douta=16'ha48f;
12384: douta=16'hb510;
12385: douta=16'hbd10;
12386: douta=16'hd5d3;
12387: douta=16'h62aa;
12388: douta=16'hbd32;
12389: douta=16'hcd93;
12390: douta=16'hd5f4;
12391: douta=16'hde15;
12392: douta=16'hd5b3;
12393: douta=16'hacf3;
12394: douta=16'h9c94;
12395: douta=16'h9cb4;
12396: douta=16'h9cb4;
12397: douta=16'h8c53;
12398: douta=16'h8433;
12399: douta=16'h7390;
12400: douta=16'h6b2d;
12401: douta=16'h41c7;
12402: douta=16'h3144;
12403: douta=16'h2903;
12404: douta=16'h31ea;
12405: douta=16'h52ac;
12406: douta=16'h2126;
12407: douta=16'h2127;
12408: douta=16'h5a8a;
12409: douta=16'h59e6;
12410: douta=16'h59c6;
12411: douta=16'h59e6;
12412: douta=16'h6206;
12413: douta=16'h6206;
12414: douta=16'h6206;
12415: douta=16'h6206;
12416: douta=16'hb534;
12417: douta=16'had15;
12418: douta=16'hcdd6;
12419: douta=16'hbd55;
12420: douta=16'h9493;
12421: douta=16'ha4f5;
12422: douta=16'h94b5;
12423: douta=16'h8453;
12424: douta=16'h8c75;
12425: douta=16'h20c3;
12426: douta=16'h20e3;
12427: douta=16'h20c3;
12428: douta=16'h20c3;
12429: douta=16'h20c3;
12430: douta=16'h1881;
12431: douta=16'h20a2;
12432: douta=16'h20a2;
12433: douta=16'h20a2;
12434: douta=16'h20c2;
12435: douta=16'h28c2;
12436: douta=16'h28c2;
12437: douta=16'h30e2;
12438: douta=16'h3103;
12439: douta=16'h3903;
12440: douta=16'h10a4;
12441: douta=16'h4964;
12442: douta=16'h51a4;
12443: douta=16'h59a4;
12444: douta=16'h59c4;
12445: douta=16'h61c3;
12446: douta=16'h940c;
12447: douta=16'h7224;
12448: douta=16'h7224;
12449: douta=16'h7a44;
12450: douta=16'h82a4;
12451: douta=16'h7aa5;
12452: douta=16'h8265;
12453: douta=16'h8285;
12454: douta=16'h82a4;
12455: douta=16'h8ac5;
12456: douta=16'h9305;
12457: douta=16'h9b25;
12458: douta=16'ha346;
12459: douta=16'hab66;
12460: douta=16'hab85;
12461: douta=16'hb3c6;
12462: douta=16'hb3a6;
12463: douta=16'hbbe6;
12464: douta=16'hbbe5;
12465: douta=16'hc405;
12466: douta=16'hc406;
12467: douta=16'hc406;
12468: douta=16'hc426;
12469: douta=16'hc426;
12470: douta=16'hc446;
12471: douta=16'hcc26;
12472: douta=16'hcc27;
12473: douta=16'hcc47;
12474: douta=16'hcc47;
12475: douta=16'hcc47;
12476: douta=16'hcc47;
12477: douta=16'hcc68;
12478: douta=16'hcc66;
12479: douta=16'hcc67;
12480: douta=16'hcc67;
12481: douta=16'hcc87;
12482: douta=16'hd467;
12483: douta=16'hd468;
12484: douta=16'hd467;
12485: douta=16'hcc67;
12486: douta=16'hd488;
12487: douta=16'hd487;
12488: douta=16'hd467;
12489: douta=16'hcc45;
12490: douta=16'hcc25;
12491: douta=16'hcc25;
12492: douta=16'hcc89;
12493: douta=16'hd52e;
12494: douta=16'hddf2;
12495: douta=16'he6b6;
12496: douta=16'hf77b;
12497: douta=16'hf79b;
12498: douta=16'hfffd;
12499: douta=16'hf799;
12500: douta=16'heed6;
12501: douta=16'he612;
12502: douta=16'hcd0c;
12503: douta=16'h7b6c;
12504: douta=16'h734b;
12505: douta=16'h7b6c;
12506: douta=16'h7b4c;
12507: douta=16'h944f;
12508: douta=16'hacd0;
12509: douta=16'hacaf;
12510: douta=16'h9c2e;
12511: douta=16'hde35;
12512: douta=16'hd5f5;
12513: douta=16'hd5f4;
12514: douta=16'hc5b4;
12515: douta=16'hc5d4;
12516: douta=16'hacd1;
12517: douta=16'hd5b4;
12518: douta=16'hacb3;
12519: douta=16'h9453;
12520: douta=16'h8453;
12521: douta=16'h7bf1;
12522: douta=16'h7bf1;
12523: douta=16'h7bd1;
12524: douta=16'h6b0d;
12525: douta=16'h49e7;
12526: douta=16'h18a2;
12527: douta=16'h3144;
12528: douta=16'h5208;
12529: douta=16'h6aea;
12530: douta=16'h734e;
12531: douta=16'h52cd;
12532: douta=16'h5b31;
12533: douta=16'h6b4f;
12534: douta=16'h320b;
12535: douta=16'h2127;
12536: douta=16'h0022;
12537: douta=16'h6206;
12538: douta=16'h6207;
12539: douta=16'h61e6;
12540: douta=16'h61c5;
12541: douta=16'h59a5;
12542: douta=16'h6a47;
12543: douta=16'h7b4b;
12544: douta=16'hc554;
12545: douta=16'had34;
12546: douta=16'hc596;
12547: douta=16'had15;
12548: douta=16'h9494;
12549: douta=16'h94b4;
12550: douta=16'h94b5;
12551: douta=16'h8c95;
12552: douta=16'h73f2;
12553: douta=16'h20c3;
12554: douta=16'h20c3;
12555: douta=16'h20e3;
12556: douta=16'h20a3;
12557: douta=16'h20c3;
12558: douta=16'h20a2;
12559: douta=16'h1881;
12560: douta=16'h20a2;
12561: douta=16'h28e2;
12562: douta=16'h20c2;
12563: douta=16'h28c3;
12564: douta=16'h28e3;
12565: douta=16'h30e2;
12566: douta=16'h3103;
12567: douta=16'h4185;
12568: douta=16'h18e4;
12569: douta=16'h4984;
12570: douta=16'h51a4;
12571: douta=16'h59c4;
12572: douta=16'h59c4;
12573: douta=16'h6a25;
12574: douta=16'h7ae7;
12575: douta=16'h7245;
12576: douta=16'h7244;
12577: douta=16'h7a64;
12578: douta=16'h7224;
12579: douta=16'h82a5;
12580: douta=16'h8285;
12581: douta=16'h8aa5;
12582: douta=16'h8ac5;
12583: douta=16'h8ac5;
12584: douta=16'h9305;
12585: douta=16'h9b26;
12586: douta=16'ha325;
12587: douta=16'hab66;
12588: douta=16'hab85;
12589: douta=16'hb3c6;
12590: douta=16'hbbc6;
12591: douta=16'hbbe6;
12592: douta=16'hbbe5;
12593: douta=16'hbbe5;
12594: douta=16'hc406;
12595: douta=16'hc406;
12596: douta=16'hc406;
12597: douta=16'hc427;
12598: douta=16'hc426;
12599: douta=16'hc446;
12600: douta=16'hc446;
12601: douta=16'hcc67;
12602: douta=16'hcc47;
12603: douta=16'hcc67;
12604: douta=16'hcc47;
12605: douta=16'hcc67;
12606: douta=16'hcc67;
12607: douta=16'hcc46;
12608: douta=16'hcc25;
12609: douta=16'hcc04;
12610: douta=16'hcc25;
12611: douta=16'hccaa;
12612: douta=16'hd56f;
12613: douta=16'he655;
12614: douta=16'hef5a;
12615: douta=16'hf7dc;
12616: douta=16'hfffd;
12617: douta=16'hffdb;
12618: douta=16'hf738;
12619: douta=16'he673;
12620: douta=16'hddaf;
12621: douta=16'hd4ea;
12622: douta=16'hcc87;
12623: douta=16'hcc46;
12624: douta=16'hcc46;
12625: douta=16'hcc68;
12626: douta=16'hd489;
12627: douta=16'hd489;
12628: douta=16'hcc68;
12629: douta=16'hcc68;
12630: douta=16'hd466;
12631: douta=16'h942e;
12632: douta=16'h9c6f;
12633: douta=16'h9c6f;
12634: douta=16'h9c6f;
12635: douta=16'hb511;
12636: douta=16'hc552;
12637: douta=16'hc593;
12638: douta=16'hac90;
12639: douta=16'hacd2;
12640: douta=16'hb514;
12641: douta=16'h9452;
12642: douta=16'hb512;
12643: douta=16'h9453;
12644: douta=16'hddf5;
12645: douta=16'h9494;
12646: douta=16'h7c11;
12647: douta=16'h73d1;
12648: douta=16'h5acd;
12649: douta=16'h49e7;
12650: douta=16'h1881;
12651: douta=16'h2103;
12652: douta=16'h41e5;
12653: douta=16'h5247;
12654: douta=16'h5a48;
12655: douta=16'h730c;
12656: douta=16'h83cd;
12657: douta=16'h9c2e;
12658: douta=16'h5249;
12659: douta=16'h424b;
12660: douta=16'h3a2b;
12661: douta=16'h4a4b;
12662: douta=16'h3a0b;
12663: douta=16'h2126;
12664: douta=16'h0883;
12665: douta=16'h18e4;
12666: douta=16'ha4b2;
12667: douta=16'h8c0e;
12668: douta=16'h730a;
12669: douta=16'h6a68;
12670: douta=16'h6226;
12671: douta=16'h6a05;
12672: douta=16'hb555;
12673: douta=16'hcdb6;
12674: douta=16'hbd75;
12675: douta=16'h94b4;
12676: douta=16'h9cb4;
12677: douta=16'h94d5;
12678: douta=16'h8cb5;
12679: douta=16'h9d17;
12680: douta=16'h2061;
12681: douta=16'h20e3;
12682: douta=16'h20c3;
12683: douta=16'h20e3;
12684: douta=16'h20a3;
12685: douta=16'h20c3;
12686: douta=16'h2082;
12687: douta=16'h20a2;
12688: douta=16'h20a2;
12689: douta=16'h20a2;
12690: douta=16'h20c2;
12691: douta=16'h28e2;
12692: douta=16'h30e2;
12693: douta=16'h30e3;
12694: douta=16'h3903;
12695: douta=16'h4209;
12696: douta=16'h3903;
12697: douta=16'h51a4;
12698: douta=16'h51a3;
12699: douta=16'h59a4;
12700: douta=16'h61e4;
12701: douta=16'h6ac9;
12702: douta=16'h6a03;
12703: douta=16'h7244;
12704: douta=16'h7a44;
12705: douta=16'h7a64;
12706: douta=16'h51c4;
12707: douta=16'h8285;
12708: douta=16'h82a5;
12709: douta=16'h8ac5;
12710: douta=16'h8ac5;
12711: douta=16'h8ac5;
12712: douta=16'h9305;
12713: douta=16'ha326;
12714: douta=16'ha346;
12715: douta=16'haba6;
12716: douta=16'hb3a5;
12717: douta=16'hb3c6;
12718: douta=16'hbbc6;
12719: douta=16'hbbe6;
12720: douta=16'hbbe6;
12721: douta=16'hbc05;
12722: douta=16'hc406;
12723: douta=16'hc426;
12724: douta=16'hc427;
12725: douta=16'hc425;
12726: douta=16'hc405;
12727: douta=16'hc3e3;
12728: douta=16'hc404;
12729: douta=16'hc447;
12730: douta=16'hcccb;
12731: douta=16'hddb0;
12732: douta=16'he6d7;
12733: douta=16'hf77b;
12734: douta=16'hffdc;
12735: douta=16'hffdc;
12736: douta=16'hf759;
12737: douta=16'he694;
12738: douta=16'hddd0;
12739: douta=16'hd52b;
12740: douta=16'hd489;
12741: douta=16'hcc45;
12742: douta=16'hcc46;
12743: douta=16'hcc47;
12744: douta=16'hd467;
12745: douta=16'hd467;
12746: douta=16'hcc87;
12747: douta=16'hd488;
12748: douta=16'hd488;
12749: douta=16'hd488;
12750: douta=16'hcc88;
12751: douta=16'hcc88;
12752: douta=16'hd488;
12753: douta=16'hcc88;
12754: douta=16'hd488;
12755: douta=16'hcc88;
12756: douta=16'hcc67;
12757: douta=16'hcc68;
12758: douta=16'hd467;
12759: douta=16'h9c70;
12760: douta=16'h9c2f;
12761: douta=16'ha4b0;
12762: douta=16'hbd31;
12763: douta=16'hcd94;
12764: douta=16'hcdd4;
12765: douta=16'hd5f5;
12766: douta=16'hb4d2;
12767: douta=16'hacf4;
12768: douta=16'hbd74;
12769: douta=16'h8c74;
12770: douta=16'h73f2;
12771: douta=16'h8433;
12772: douta=16'h6370;
12773: douta=16'h4a6a;
12774: douta=16'h18a3;
12775: douta=16'h2923;
12776: douta=16'h3145;
12777: douta=16'h5227;
12778: douta=16'h732a;
12779: douta=16'h6ac9;
12780: douta=16'h734b;
12781: douta=16'h7b4b;
12782: douta=16'h7b6b;
12783: douta=16'ha46f;
12784: douta=16'hac8f;
12785: douta=16'ha46f;
12786: douta=16'h8bee;
12787: douta=16'h3a2b;
12788: douta=16'h18e5;
12789: douta=16'h0882;
12790: douta=16'h10a4;
12791: douta=16'h10e5;
12792: douta=16'h2167;
12793: douta=16'h1948;
12794: douta=16'h82a7;
12795: douta=16'h7286;
12796: douta=16'h7a67;
12797: douta=16'h7a87;
12798: douta=16'h7a87;
12799: douta=16'h7a87;
12800: douta=16'hacf5;
12801: douta=16'hcdf6;
12802: douta=16'hbd75;
12803: douta=16'h8412;
12804: douta=16'ha4f5;
12805: douta=16'h94d5;
12806: douta=16'h8454;
12807: douta=16'h8453;
12808: douta=16'h20e3;
12809: douta=16'h20c3;
12810: douta=16'h20c3;
12811: douta=16'h20e3;
12812: douta=16'h20c3;
12813: douta=16'h1882;
12814: douta=16'h20a2;
12815: douta=16'h20a2;
12816: douta=16'h20a2;
12817: douta=16'h20c2;
12818: douta=16'h28e3;
12819: douta=16'h28e2;
12820: douta=16'h3103;
12821: douta=16'h3103;
12822: douta=16'h3923;
12823: douta=16'h424b;
12824: douta=16'h5184;
12825: douta=16'h5184;
12826: douta=16'h51a4;
12827: douta=16'h61c4;
12828: douta=16'h61e4;
12829: douta=16'h8c2f;
12830: douta=16'h71e3;
12831: douta=16'h7244;
12832: douta=16'h7a64;
12833: douta=16'h7a64;
12834: douta=16'h7a85;
12835: douta=16'h8aa5;
12836: douta=16'h8284;
12837: douta=16'h8aa5;
12838: douta=16'h8ac5;
12839: douta=16'h8ac5;
12840: douta=16'h9306;
12841: douta=16'h9b26;
12842: douta=16'ha345;
12843: douta=16'hab85;
12844: douta=16'hab65;
12845: douta=16'hb384;
12846: douta=16'hb364;
12847: douta=16'hbbc6;
12848: douta=16'hc44a;
12849: douta=16'hcd2d;
12850: douta=16'hde54;
12851: douta=16'hef18;
12852: douta=16'hf79b;
12853: douta=16'hf7bb;
12854: douta=16'hef58;
12855: douta=16'he694;
12856: douta=16'hddcf;
12857: douta=16'hd50b;
12858: douta=16'hcc87;
12859: douta=16'hcc27;
12860: douta=16'hcc25;
12861: douta=16'hcc46;
12862: douta=16'hcc47;
12863: douta=16'hd468;
12864: douta=16'hcc68;
12865: douta=16'hcc68;
12866: douta=16'hd488;
12867: douta=16'hd488;
12868: douta=16'hd488;
12869: douta=16'hd488;
12870: douta=16'hd488;
12871: douta=16'hd488;
12872: douta=16'hd487;
12873: douta=16'hd488;
12874: douta=16'hcc67;
12875: douta=16'hcc88;
12876: douta=16'hd488;
12877: douta=16'hd488;
12878: douta=16'hd488;
12879: douta=16'hcc68;
12880: douta=16'hcc88;
12881: douta=16'hd488;
12882: douta=16'hd488;
12883: douta=16'hd488;
12884: douta=16'hd488;
12885: douta=16'hcc68;
12886: douta=16'hd467;
12887: douta=16'h9c4e;
12888: douta=16'hacd2;
12889: douta=16'hb4f2;
12890: douta=16'hbd52;
12891: douta=16'hc594;
12892: douta=16'hacf4;
12893: douta=16'h9473;
12894: douta=16'h8432;
12895: douta=16'h6bb1;
12896: douta=16'h6bb1;
12897: douta=16'h736f;
12898: douta=16'h39a6;
12899: douta=16'h3124;
12900: douta=16'h0860;
12901: douta=16'h62ca;
12902: douta=16'h7b6b;
12903: douta=16'h8bad;
12904: douta=16'h83ad;
12905: douta=16'h838c;
12906: douta=16'h7b6b;
12907: douta=16'h9c2e;
12908: douta=16'hac8f;
12909: douta=16'hb510;
12910: douta=16'hcd71;
12911: douta=16'hcd72;
12912: douta=16'hc551;
12913: douta=16'hac8f;
12914: douta=16'h9410;
12915: douta=16'h632d;
12916: douta=16'h31a8;
12917: douta=16'h2126;
12918: douta=16'h2987;
12919: douta=16'h10c4;
12920: douta=16'h10c4;
12921: douta=16'h2169;
12922: douta=16'h59e6;
12923: douta=16'h7aa6;
12924: douta=16'h82a7;
12925: douta=16'h82a7;
12926: douta=16'h82a7;
12927: douta=16'h82a7;
12928: douta=16'had35;
12929: douta=16'hc5b5;
12930: douta=16'hb555;
12931: douta=16'ha557;
12932: douta=16'h9cf5;
12933: douta=16'h94d5;
12934: douta=16'h8c95;
12935: douta=16'h1060;
12936: douta=16'h20e3;
12937: douta=16'h20e3;
12938: douta=16'h20c3;
12939: douta=16'h20c3;
12940: douta=16'h20c3;
12941: douta=16'h1882;
12942: douta=16'h20a2;
12943: douta=16'h20a2;
12944: douta=16'h20a2;
12945: douta=16'h20c2;
12946: douta=16'h28e2;
12947: douta=16'h28e2;
12948: douta=16'h3123;
12949: douta=16'h3103;
12950: douta=16'h3923;
12951: douta=16'h424a;
12952: douta=16'h51a4;
12953: douta=16'h51a4;
12954: douta=16'h59a4;
12955: douta=16'h59c4;
12956: douta=16'h61e4;
12957: douta=16'hb594;
12958: douta=16'h7224;
12959: douta=16'h7244;
12960: douta=16'h7a64;
12961: douta=16'h7a85;
12962: douta=16'h8aa4;
12963: douta=16'h8244;
12964: douta=16'h7a24;
12965: douta=16'h82c6;
12966: douta=16'h9369;
12967: douta=16'hb4af;
12968: douta=16'hc592;
12969: douta=16'hde96;
12970: douta=16'he718;
12971: douta=16'hf779;
12972: douta=16'hef17;
12973: douta=16'hde32;
12974: douta=16'hd54d;
12975: douta=16'hc4ca;
12976: douta=16'hbc27;
12977: douta=16'hbbe5;
12978: douta=16'hc3c5;
12979: douta=16'hc3e5;
12980: douta=16'hc426;
12981: douta=16'hc427;
12982: douta=16'hc446;
12983: douta=16'hcc47;
12984: douta=16'hcc67;
12985: douta=16'hcc47;
12986: douta=16'hcc68;
12987: douta=16'hcc47;
12988: douta=16'hcc67;
12989: douta=16'hcc48;
12990: douta=16'hcc67;
12991: douta=16'hcc68;
12992: douta=16'hcc68;
12993: douta=16'hcc68;
12994: douta=16'hcc88;
12995: douta=16'hcc68;
12996: douta=16'hcc68;
12997: douta=16'hd488;
12998: douta=16'hd488;
12999: douta=16'hd488;
13000: douta=16'hd487;
13001: douta=16'hd488;
13002: douta=16'hcc88;
13003: douta=16'hcc88;
13004: douta=16'hcc88;
13005: douta=16'hd488;
13006: douta=16'hd488;
13007: douta=16'hd488;
13008: douta=16'hd488;
13009: douta=16'hcc68;
13010: douta=16'hd489;
13011: douta=16'hd488;
13012: douta=16'hcc46;
13013: douta=16'hcc25;
13014: douta=16'hcc67;
13015: douta=16'hccec;
13016: douta=16'hacd2;
13017: douta=16'hacd2;
13018: douta=16'hacd3;
13019: douta=16'h9cb4;
13020: douta=16'h8412;
13021: douta=16'h7bf2;
13022: douta=16'h738f;
13023: douta=16'h3944;
13024: douta=16'h41c4;
13025: douta=16'h72e9;
13026: douta=16'h838b;
13027: douta=16'h8bcd;
13028: douta=16'h942e;
13029: douta=16'h9c6f;
13030: douta=16'hbd51;
13031: douta=16'h730b;
13032: douta=16'hacd1;
13033: douta=16'hbd52;
13034: douta=16'hbd31;
13035: douta=16'hd5b3;
13036: douta=16'hd5b3;
13037: douta=16'hd5b3;
13038: douta=16'hcd52;
13039: douta=16'hc532;
13040: douta=16'hb4d1;
13041: douta=16'hac91;
13042: douta=16'h8bf0;
13043: douta=16'h8c10;
13044: douta=16'h5b0d;
13045: douta=16'h3a2a;
13046: douta=16'h2126;
13047: douta=16'h1906;
13048: douta=16'h18c4;
13049: douta=16'h1128;
13050: douta=16'h936a;
13051: douta=16'h8ac7;
13052: douta=16'h8ac7;
13053: douta=16'h8ac7;
13054: douta=16'h8ac7;
13055: douta=16'h8ae7;
13056: douta=16'hcdb5;
13057: douta=16'hc596;
13058: douta=16'h9494;
13059: douta=16'had57;
13060: douta=16'h9cf6;
13061: douta=16'h8c75;
13062: douta=16'ha558;
13063: douta=16'h3165;
13064: douta=16'h1882;
13065: douta=16'h20e3;
13066: douta=16'h20e3;
13067: douta=16'h20e3;
13068: douta=16'h20c3;
13069: douta=16'h18a2;
13070: douta=16'h20a2;
13071: douta=16'h20c2;
13072: douta=16'h20a2;
13073: douta=16'h20a2;
13074: douta=16'h28e2;
13075: douta=16'h28e2;
13076: douta=16'h3103;
13077: douta=16'h3923;
13078: douta=16'h3923;
13079: douta=16'h31a8;
13080: douta=16'h5184;
13081: douta=16'h5163;
13082: douta=16'h5163;
13083: douta=16'h5984;
13084: douta=16'h61e4;
13085: douta=16'had51;
13086: douta=16'h9c4c;
13087: douta=16'hb4f1;
13088: douta=16'hce13;
13089: douta=16'hd674;
13090: douta=16'hd654;
13091: douta=16'h8ba9;
13092: douta=16'hb4cd;
13093: douta=16'ha42b;
13094: douta=16'h9b88;
13095: douta=16'h8ae5;
13096: douta=16'h92c5;
13097: douta=16'h9b05;
13098: douta=16'hab46;
13099: douta=16'hab87;
13100: douta=16'hb3c7;
13101: douta=16'hbbc7;
13102: douta=16'hbbc6;
13103: douta=16'hbbe7;
13104: douta=16'hc406;
13105: douta=16'hc406;
13106: douta=16'hc427;
13107: douta=16'hc447;
13108: douta=16'hc427;
13109: douta=16'hc427;
13110: douta=16'hcc47;
13111: douta=16'hcc47;
13112: douta=16'hcc67;
13113: douta=16'hcc67;
13114: douta=16'hcc67;
13115: douta=16'hcc68;
13116: douta=16'hcc67;
13117: douta=16'hcc67;
13118: douta=16'hcc68;
13119: douta=16'hcc68;
13120: douta=16'hcc88;
13121: douta=16'hcc68;
13122: douta=16'hd488;
13123: douta=16'hcc68;
13124: douta=16'hd488;
13125: douta=16'hcc88;
13126: douta=16'hd488;
13127: douta=16'hd488;
13128: douta=16'hd487;
13129: douta=16'hcc46;
13130: douta=16'hcc25;
13131: douta=16'hcc26;
13132: douta=16'hcc89;
13133: douta=16'hd50d;
13134: douta=16'hddb1;
13135: douta=16'he655;
13136: douta=16'hef19;
13137: douta=16'hf79c;
13138: douta=16'hfffe;
13139: douta=16'hf758;
13140: douta=16'hee94;
13141: douta=16'he5d0;
13142: douta=16'hd50a;
13143: douta=16'hd486;
13144: douta=16'ha4b2;
13145: douta=16'ha492;
13146: douta=16'h9432;
13147: douta=16'h83f0;
13148: douta=16'h49c6;
13149: douta=16'h49e6;
13150: douta=16'h62a9;
13151: douta=16'h7b2b;
13152: douta=16'h838b;
13153: douta=16'ha42e;
13154: douta=16'hac8f;
13155: douta=16'h8bed;
13156: douta=16'hd593;
13157: douta=16'hacd1;
13158: douta=16'h736d;
13159: douta=16'he615;
13160: douta=16'hc573;
13161: douta=16'hb513;
13162: douta=16'h9472;
13163: douta=16'h7bf1;
13164: douta=16'h7bd1;
13165: douta=16'h8c74;
13166: douta=16'h8c74;
13167: douta=16'h8c74;
13168: douta=16'h9473;
13169: douta=16'h9473;
13170: douta=16'h8412;
13171: douta=16'h9453;
13172: douta=16'h73d2;
13173: douta=16'h73f2;
13174: douta=16'h428e;
13175: douta=16'h320a;
13176: douta=16'h2946;
13177: douta=16'h1907;
13178: douta=16'h5acb;
13179: douta=16'h92e8;
13180: douta=16'h92e8;
13181: douta=16'h8ae7;
13182: douta=16'h8ae8;
13183: douta=16'h9307;
13184: douta=16'hcdd6;
13185: douta=16'hbd95;
13186: douta=16'h9453;
13187: douta=16'h9cf5;
13188: douta=16'h94d5;
13189: douta=16'h8433;
13190: douta=16'h2103;
13191: douta=16'h20c3;
13192: douta=16'h3987;
13193: douta=16'h426b;
13194: douta=16'h2104;
13195: douta=16'h20a2;
13196: douta=16'h20e3;
13197: douta=16'h20a2;
13198: douta=16'h2082;
13199: douta=16'h1861;
13200: douta=16'h2081;
13201: douta=16'h2082;
13202: douta=16'h28e3;
13203: douta=16'h3965;
13204: douta=16'h5227;
13205: douta=16'h62c9;
13206: douta=16'h7b6c;
13207: douta=16'h1906;
13208: douta=16'h9c90;
13209: douta=16'h944e;
13210: douta=16'h8bcb;
13211: douta=16'h7b29;
13212: douta=16'h72a6;
13213: douta=16'h7224;
13214: douta=16'h7224;
13215: douta=16'h7203;
13216: douta=16'h7a44;
13217: douta=16'h8285;
13218: douta=16'h82a6;
13219: douta=16'h51a4;
13220: douta=16'h8ac6;
13221: douta=16'h92e5;
13222: douta=16'h92e5;
13223: douta=16'h9306;
13224: douta=16'h9306;
13225: douta=16'ha366;
13226: douta=16'hab86;
13227: douta=16'hb3a6;
13228: douta=16'hb3c7;
13229: douta=16'hbbe7;
13230: douta=16'hbbc6;
13231: douta=16'hbbe6;
13232: douta=16'hc407;
13233: douta=16'hc407;
13234: douta=16'hc406;
13235: douta=16'hc426;
13236: douta=16'hc447;
13237: douta=16'hcc47;
13238: douta=16'hc446;
13239: douta=16'hcc47;
13240: douta=16'hcc47;
13241: douta=16'hcc67;
13242: douta=16'hcc68;
13243: douta=16'hcc48;
13244: douta=16'hcc67;
13245: douta=16'hcc67;
13246: douta=16'hcc25;
13247: douta=16'hcc25;
13248: douta=16'hc404;
13249: douta=16'hcc68;
13250: douta=16'hd50b;
13251: douta=16'hdd8f;
13252: douta=16'hde34;
13253: douta=16'heef8;
13254: douta=16'hf79c;
13255: douta=16'hffdc;
13256: douta=16'hffdb;
13257: douta=16'hf738;
13258: douta=16'heeb5;
13259: douta=16'hddcf;
13260: douta=16'hd54d;
13261: douta=16'hcca9;
13262: douta=16'hcc66;
13263: douta=16'hcc26;
13264: douta=16'hcc46;
13265: douta=16'had11;
13266: douta=16'hcc26;
13267: douta=16'hd4a9;
13268: douta=16'hd488;
13269: douta=16'hcc88;
13270: douta=16'hcc89;
13271: douta=16'hcc68;
13272: douta=16'h9493;
13273: douta=16'h62aa;
13274: douta=16'h3985;
13275: douta=16'h730a;
13276: douta=16'h7b4b;
13277: douta=16'h8c0e;
13278: douta=16'h940d;
13279: douta=16'hacaf;
13280: douta=16'hbd11;
13281: douta=16'hcd73;
13282: douta=16'hc572;
13283: douta=16'h8bad;
13284: douta=16'hd5b3;
13285: douta=16'hacb3;
13286: douta=16'h9473;
13287: douta=16'h7390;
13288: douta=16'hacb3;
13289: douta=16'h8c32;
13290: douta=16'h83f1;
13291: douta=16'h7390;
13292: douta=16'h630e;
13293: douta=16'h738f;
13294: douta=16'h73b0;
13295: douta=16'h6b4f;
13296: douta=16'h7390;
13297: douta=16'h73b1;
13298: douta=16'h73d1;
13299: douta=16'h6b70;
13300: douta=16'h7bf3;
13301: douta=16'h6370;
13302: douta=16'h7c75;
13303: douta=16'h3a2a;
13304: douta=16'h29c9;
13305: douta=16'hffff;
13306: douta=16'hffff;
13307: douta=16'h9b49;
13308: douta=16'h9308;
13309: douta=16'h9328;
13310: douta=16'h9307;
13311: douta=16'h9328;
13312: douta=16'hcdd6;
13313: douta=16'hb555;
13314: douta=16'had57;
13315: douta=16'ha516;
13316: douta=16'h9cf6;
13317: douta=16'ha558;
13318: douta=16'h28e3;
13319: douta=16'h28e3;
13320: douta=16'h20c3;
13321: douta=16'h28c3;
13322: douta=16'h20e3;
13323: douta=16'h31c8;
13324: douta=16'h39e9;
13325: douta=16'h31c7;
13326: douta=16'h31c7;
13327: douta=16'h3165;
13328: douta=16'h3144;
13329: douta=16'h3124;
13330: douta=16'h3103;
13331: douta=16'h30e2;
13332: douta=16'h30e2;
13333: douta=16'h3902;
13334: douta=16'h41a6;
13335: douta=16'h10a5;
13336: douta=16'h51a4;
13337: douta=16'h59c4;
13338: douta=16'h61e4;
13339: douta=16'h69e4;
13340: douta=16'h7224;
13341: douta=16'h7244;
13342: douta=16'h7a65;
13343: douta=16'h7a64;
13344: douta=16'h8285;
13345: douta=16'h82a5;
13346: douta=16'h82c6;
13347: douta=16'h6a24;
13348: douta=16'h8ac6;
13349: douta=16'h9306;
13350: douta=16'h9306;
13351: douta=16'h9306;
13352: douta=16'h9b47;
13353: douta=16'hab87;
13354: douta=16'haba7;
13355: douta=16'hb3a7;
13356: douta=16'hb3c7;
13357: douta=16'hbbe7;
13358: douta=16'hbbe6;
13359: douta=16'hc3e7;
13360: douta=16'hc407;
13361: douta=16'hc427;
13362: douta=16'hc406;
13363: douta=16'hc406;
13364: douta=16'hc3e3;
13365: douta=16'hc404;
13366: douta=16'hcc28;
13367: douta=16'hcccb;
13368: douta=16'hd56f;
13369: douta=16'hde33;
13370: douta=16'heed8;
13371: douta=16'hf77a;
13372: douta=16'hf7dc;
13373: douta=16'hf79b;
13374: douta=16'hef37;
13375: douta=16'heeb4;
13376: douta=16'hddd1;
13377: douta=16'hd52c;
13378: douta=16'hcca8;
13379: douta=16'hcc66;
13380: douta=16'hcc26;
13381: douta=16'hcc45;
13382: douta=16'hd467;
13383: douta=16'hd488;
13384: douta=16'hcc88;
13385: douta=16'hd488;
13386: douta=16'hd488;
13387: douta=16'hd488;
13388: douta=16'hd488;
13389: douta=16'hcc88;
13390: douta=16'hd488;
13391: douta=16'hd4a9;
13392: douta=16'hcc69;
13393: douta=16'had31;
13394: douta=16'hcc25;
13395: douta=16'hcc68;
13396: douta=16'hcc88;
13397: douta=16'hcc68;
13398: douta=16'hcc68;
13399: douta=16'hcc69;
13400: douta=16'h9beb;
13401: douta=16'h7b4a;
13402: douta=16'h83ad;
13403: douta=16'hac90;
13404: douta=16'hac8f;
13405: douta=16'hb4f0;
13406: douta=16'hc552;
13407: douta=16'hd5b3;
13408: douta=16'hcd93;
13409: douta=16'hcd53;
13410: douta=16'hb511;
13411: douta=16'hacb2;
13412: douta=16'h83d1;
13413: douta=16'h9474;
13414: douta=16'h8c74;
13415: douta=16'h6b70;
13416: douta=16'h7b90;
13417: douta=16'h736f;
13418: douta=16'h6b4f;
13419: douta=16'h6b6f;
13420: douta=16'h634e;
13421: douta=16'h632f;
13422: douta=16'h62cd;
13423: douta=16'h62cd;
13424: douta=16'h62cc;
13425: douta=16'h62cc;
13426: douta=16'h6b0d;
13427: douta=16'h6b4f;
13428: douta=16'h4aad;
13429: douta=16'h6bb1;
13430: douta=16'h8c73;
13431: douta=16'h4acf;
13432: douta=16'h39cc;
13433: douta=16'hffff;
13434: douta=16'hffff;
13435: douta=16'h7aa6;
13436: douta=16'h9b28;
13437: douta=16'h9b48;
13438: douta=16'h9b28;
13439: douta=16'h9b48;
13440: douta=16'hc595;
13441: douta=16'h9494;
13442: douta=16'had36;
13443: douta=16'ha4f5;
13444: douta=16'h8c94;
13445: douta=16'h31c7;
13446: douta=16'h28e4;
13447: douta=16'h28e3;
13448: douta=16'h28e3;
13449: douta=16'h20e3;
13450: douta=16'h20e3;
13451: douta=16'h20e3;
13452: douta=16'h18a2;
13453: douta=16'h20a2;
13454: douta=16'h20c2;
13455: douta=16'h20a2;
13456: douta=16'h20c2;
13457: douta=16'h28e3;
13458: douta=16'h28e3;
13459: douta=16'h3123;
13460: douta=16'h3943;
13461: douta=16'h4144;
13462: douta=16'h4a49;
13463: douta=16'h18a5;
13464: douta=16'h51a4;
13465: douta=16'h61e4;
13466: douta=16'h61e4;
13467: douta=16'h6a04;
13468: douta=16'h7224;
13469: douta=16'h7a64;
13470: douta=16'h7a65;
13471: douta=16'h8286;
13472: douta=16'h7a85;
13473: douta=16'h82a5;
13474: douta=16'h82c5;
13475: douta=16'h9326;
13476: douta=16'h9b26;
13477: douta=16'h9306;
13478: douta=16'h9305;
13479: douta=16'h9326;
13480: douta=16'h9306;
13481: douta=16'ha326;
13482: douta=16'ha325;
13483: douta=16'hab64;
13484: douta=16'hb3c6;
13485: douta=16'hc4ac;
13486: douta=16'hcd70;
13487: douta=16'hde53;
13488: douta=16'he718;
13489: douta=16'hf77a;
13490: douta=16'hf79a;
13491: douta=16'hef38;
13492: douta=16'he6b4;
13493: douta=16'hddf1;
13494: douta=16'hcd4d;
13495: douta=16'hcca8;
13496: douta=16'hcc46;
13497: douta=16'hcc25;
13498: douta=16'hcc25;
13499: douta=16'hcc46;
13500: douta=16'hcc67;
13501: douta=16'hcc67;
13502: douta=16'hcc68;
13503: douta=16'hcc67;
13504: douta=16'hcc68;
13505: douta=16'hd488;
13506: douta=16'hcc68;
13507: douta=16'hcc88;
13508: douta=16'hcc88;
13509: douta=16'hcc88;
13510: douta=16'hd488;
13511: douta=16'hcc88;
13512: douta=16'hcc88;
13513: douta=16'hcc88;
13514: douta=16'hd488;
13515: douta=16'hd4a9;
13516: douta=16'hd489;
13517: douta=16'hd4a9;
13518: douta=16'hd488;
13519: douta=16'hd488;
13520: douta=16'hd488;
13521: douta=16'had31;
13522: douta=16'hcc26;
13523: douta=16'hcc68;
13524: douta=16'hcc68;
13525: douta=16'hcc88;
13526: douta=16'hcc68;
13527: douta=16'hcc68;
13528: douta=16'ha40a;
13529: douta=16'h8bcd;
13530: douta=16'h9c2f;
13531: douta=16'hbd12;
13532: douta=16'hc553;
13533: douta=16'hbd73;
13534: douta=16'hcdb4;
13535: douta=16'hcd92;
13536: douta=16'hacd2;
13537: douta=16'h8c32;
13538: douta=16'h9432;
13539: douta=16'h8c32;
13540: douta=16'h83f2;
13541: douta=16'h7bb0;
13542: douta=16'h630d;
13543: douta=16'h630e;
13544: douta=16'h62ed;
13545: douta=16'h736f;
13546: douta=16'h5acc;
13547: douta=16'h5acc;
13548: douta=16'h5aab;
13549: douta=16'h526a;
13550: douta=16'h62ac;
13551: douta=16'h8c32;
13552: douta=16'h8413;
13553: douta=16'h8432;
13554: douta=16'h632f;
13555: douta=16'h634e;
13556: douta=16'hb5d7;
13557: douta=16'h6c94;
13558: douta=16'hce7b;
13559: douta=16'hddb2;
13560: douta=16'hb2c5;
13561: douta=16'ha368;
13562: douta=16'ha368;
13563: douta=16'ha369;
13564: douta=16'ha369;
13565: douta=16'h9b48;
13566: douta=16'ha349;
13567: douta=16'h9b48;
13568: douta=16'hbd95;
13569: douta=16'h8c53;
13570: douta=16'ha515;
13571: douta=16'ha4d5;
13572: douta=16'h9d38;
13573: douta=16'h2041;
13574: douta=16'h28e3;
13575: douta=16'h28e3;
13576: douta=16'h28e3;
13577: douta=16'h28e3;
13578: douta=16'h20e3;
13579: douta=16'h20e3;
13580: douta=16'h1882;
13581: douta=16'h20a2;
13582: douta=16'h20a2;
13583: douta=16'h20a2;
13584: douta=16'h28e3;
13585: douta=16'h28e3;
13586: douta=16'h3103;
13587: douta=16'h3123;
13588: douta=16'h3944;
13589: douta=16'h4143;
13590: douta=16'h424a;
13591: douta=16'h3104;
13592: douta=16'h59a4;
13593: douta=16'h61c4;
13594: douta=16'h6204;
13595: douta=16'h6a24;
13596: douta=16'h7224;
13597: douta=16'h7a64;
13598: douta=16'h7a44;
13599: douta=16'h7a24;
13600: douta=16'h7a44;
13601: douta=16'h8285;
13602: douta=16'h8b28;
13603: douta=16'ha42b;
13604: douta=16'h9bcb;
13605: douta=16'hcdf2;
13606: douta=16'hd674;
13607: douta=16'hde73;
13608: douta=16'hd653;
13609: douta=16'hd5d1;
13610: douta=16'hc52e;
13611: douta=16'hbcab;
13612: douta=16'hbc28;
13613: douta=16'hbbe6;
13614: douta=16'hbba5;
13615: douta=16'hbba4;
13616: douta=16'hbbe5;
13617: douta=16'hc406;
13618: douta=16'hc426;
13619: douta=16'hc447;
13620: douta=16'hc447;
13621: douta=16'hcc47;
13622: douta=16'hcc47;
13623: douta=16'hcc47;
13624: douta=16'hcc67;
13625: douta=16'hcc67;
13626: douta=16'hcc47;
13627: douta=16'hcc67;
13628: douta=16'hcc68;
13629: douta=16'hcc68;
13630: douta=16'hcc67;
13631: douta=16'hcc68;
13632: douta=16'hcc88;
13633: douta=16'hcc68;
13634: douta=16'hcc68;
13635: douta=16'hcc68;
13636: douta=16'hcc68;
13637: douta=16'hcc88;
13638: douta=16'hd488;
13639: douta=16'hd488;
13640: douta=16'hcc88;
13641: douta=16'hd488;
13642: douta=16'hcc88;
13643: douta=16'hd489;
13644: douta=16'hd488;
13645: douta=16'hd4a9;
13646: douta=16'hd4a9;
13647: douta=16'hd489;
13648: douta=16'hcc88;
13649: douta=16'had31;
13650: douta=16'hcc25;
13651: douta=16'hcc88;
13652: douta=16'hcc88;
13653: douta=16'hcc88;
13654: douta=16'hcc88;
13655: douta=16'hcc68;
13656: douta=16'hcc69;
13657: douta=16'h9c4f;
13658: douta=16'ha4b1;
13659: douta=16'hb533;
13660: douta=16'hc574;
13661: douta=16'hb534;
13662: douta=16'ha4b3;
13663: douta=16'h8c73;
13664: douta=16'h9453;
13665: douta=16'h8c53;
13666: douta=16'h6b2f;
13667: douta=16'h6b4f;
13668: douta=16'h6b2e;
13669: douta=16'h5acd;
13670: douta=16'h630d;
13671: douta=16'h736f;
13672: douta=16'h5a8c;
13673: douta=16'h522a;
13674: douta=16'h7b8f;
13675: douta=16'ha4b3;
13676: douta=16'h83d1;
13677: douta=16'h7390;
13678: douta=16'h736f;
13679: douta=16'h5aee;
13680: douta=16'h7c73;
13681: douta=16'hffff;
13682: douta=16'hffff;
13683: douta=16'hdcd0;
13684: douta=16'h9aa3;
13685: douta=16'h9b67;
13686: douta=16'ha368;
13687: douta=16'ha367;
13688: douta=16'ha368;
13689: douta=16'ha368;
13690: douta=16'ha388;
13691: douta=16'ha368;
13692: douta=16'ha368;
13693: douta=16'ha368;
13694: douta=16'ha348;
13695: douta=16'ha349;
13696: douta=16'had56;
13697: douta=16'ha515;
13698: douta=16'had16;
13699: douta=16'ha4f5;
13700: douta=16'h634e;
13701: douta=16'h3125;
13702: douta=16'h426c;
13703: douta=16'h424b;
13704: douta=16'h28e3;
13705: douta=16'h28c3;
13706: douta=16'h20e3;
13707: douta=16'h20e3;
13708: douta=16'h20a2;
13709: douta=16'h20a2;
13710: douta=16'h20c2;
13711: douta=16'h20a2;
13712: douta=16'h28e3;
13713: douta=16'h28e2;
13714: douta=16'h28e2;
13715: douta=16'h3103;
13716: douta=16'h30c2;
13717: douta=16'h3902;
13718: douta=16'h39e9;
13719: douta=16'h51c5;
13720: douta=16'h6ac8;
13721: douta=16'h838b;
13722: douta=16'h9c6e;
13723: douta=16'had30;
13724: douta=16'hbd92;
13725: douta=16'hbd71;
13726: douta=16'hb50f;
13727: douta=16'ha44c;
13728: douta=16'h9389;
13729: douta=16'h8b07;
13730: douta=16'h8aa5;
13731: douta=16'h8285;
13732: douta=16'h51c5;
13733: douta=16'h92c5;
13734: douta=16'h9305;
13735: douta=16'h9306;
13736: douta=16'h9326;
13737: douta=16'hab86;
13738: douta=16'haba6;
13739: douta=16'hb3c7;
13740: douta=16'hbbe7;
13741: douta=16'hbbe7;
13742: douta=16'hbbe7;
13743: douta=16'hbc06;
13744: douta=16'hc407;
13745: douta=16'hc447;
13746: douta=16'hc447;
13747: douta=16'hc448;
13748: douta=16'hcc47;
13749: douta=16'hcc47;
13750: douta=16'hcc47;
13751: douta=16'hcc67;
13752: douta=16'hcc47;
13753: douta=16'hcc48;
13754: douta=16'hcc68;
13755: douta=16'hcc48;
13756: douta=16'hcc68;
13757: douta=16'hcc68;
13758: douta=16'hcc68;
13759: douta=16'hcc68;
13760: douta=16'hcc68;
13761: douta=16'hcc68;
13762: douta=16'hcc68;
13763: douta=16'hcc68;
13764: douta=16'hcc88;
13765: douta=16'hd488;
13766: douta=16'hcc68;
13767: douta=16'hcc88;
13768: douta=16'hd4a9;
13769: douta=16'hd4a9;
13770: douta=16'hcc89;
13771: douta=16'hd489;
13772: douta=16'hd488;
13773: douta=16'hd488;
13774: douta=16'hcc88;
13775: douta=16'hd4a9;
13776: douta=16'hd4a9;
13777: douta=16'had32;
13778: douta=16'hcc25;
13779: douta=16'hd488;
13780: douta=16'hcc88;
13781: douta=16'hcc89;
13782: douta=16'hcc89;
13783: douta=16'hcc69;
13784: douta=16'hd488;
13785: douta=16'h8bef;
13786: douta=16'ha492;
13787: douta=16'ha4d4;
13788: douta=16'h9cb3;
13789: douta=16'h9452;
13790: douta=16'h8412;
13791: douta=16'h6b90;
13792: douta=16'h6b4f;
13793: douta=16'h630e;
13794: douta=16'h632e;
13795: douta=16'h630e;
13796: douta=16'h5aac;
13797: douta=16'h62ed;
13798: douta=16'h83f0;
13799: douta=16'h8bf1;
13800: douta=16'h8410;
13801: douta=16'h7bb0;
13802: douta=16'h6acd;
13803: douta=16'h6b0d;
13804: douta=16'hadd7;
13805: douta=16'hffff;
13806: douta=16'hffbd;
13807: douta=16'hbb87;
13808: douta=16'ha304;
13809: douta=16'haba8;
13810: douta=16'haba7;
13811: douta=16'haba8;
13812: douta=16'hab88;
13813: douta=16'ha388;
13814: douta=16'hab88;
13815: douta=16'hab88;
13816: douta=16'hab88;
13817: douta=16'ha388;
13818: douta=16'hab88;
13819: douta=16'ha368;
13820: douta=16'ha368;
13821: douta=16'ha368;
13822: douta=16'hab68;
13823: douta=16'ha368;
13824: douta=16'h9494;
13825: douta=16'had36;
13826: douta=16'had15;
13827: douta=16'h94b5;
13828: douta=16'h1040;
13829: douta=16'h28e3;
13830: douta=16'h28e3;
13831: douta=16'h28e3;
13832: douta=16'h20c2;
13833: douta=16'h428c;
13834: douta=16'h428c;
13835: douta=16'h2925;
13836: douta=16'h2945;
13837: douta=16'h3186;
13838: douta=16'h39a6;
13839: douta=16'h41e8;
13840: douta=16'h528a;
13841: douta=16'h5aaa;
13842: douta=16'h5aca;
13843: douta=16'h62c9;
13844: douta=16'h5a47;
13845: douta=16'h5226;
13846: douta=16'h2167;
13847: douta=16'h59a4;
13848: douta=16'h5184;
13849: douta=16'h59a4;
13850: douta=16'h61c4;
13851: douta=16'h6a04;
13852: douta=16'h838c;
13853: douta=16'h7a85;
13854: douta=16'h82a5;
13855: douta=16'h82a5;
13856: douta=16'h82c5;
13857: douta=16'h8aa5;
13858: douta=16'h8ac6;
13859: douta=16'h8ac6;
13860: douta=16'h59e5;
13861: douta=16'h9326;
13862: douta=16'h9326;
13863: douta=16'h9326;
13864: douta=16'h9b26;
13865: douta=16'hab86;
13866: douta=16'hb3a7;
13867: douta=16'hb3c7;
13868: douta=16'hb3e6;
13869: douta=16'hbbe6;
13870: douta=16'hbbe7;
13871: douta=16'hc407;
13872: douta=16'hc407;
13873: douta=16'hc426;
13874: douta=16'hc426;
13875: douta=16'hc448;
13876: douta=16'hc448;
13877: douta=16'hc447;
13878: douta=16'hcc47;
13879: douta=16'hcc47;
13880: douta=16'hcc47;
13881: douta=16'hcc48;
13882: douta=16'hcc68;
13883: douta=16'hcc68;
13884: douta=16'hcc68;
13885: douta=16'hcc48;
13886: douta=16'hcc68;
13887: douta=16'hcc68;
13888: douta=16'hcc68;
13889: douta=16'hcc68;
13890: douta=16'hcc88;
13891: douta=16'hcc88;
13892: douta=16'hcc68;
13893: douta=16'hcc88;
13894: douta=16'hd4a9;
13895: douta=16'hd4a9;
13896: douta=16'hcc88;
13897: douta=16'hd488;
13898: douta=16'hd489;
13899: douta=16'hcc89;
13900: douta=16'hd489;
13901: douta=16'hd488;
13902: douta=16'hcc88;
13903: douta=16'hcc88;
13904: douta=16'hcc89;
13905: douta=16'had33;
13906: douta=16'hcc26;
13907: douta=16'hcc89;
13908: douta=16'hcc88;
13909: douta=16'hcc69;
13910: douta=16'hcc69;
13911: douta=16'hcc69;
13912: douta=16'hcc69;
13913: douta=16'h9c50;
13914: douta=16'h9451;
13915: douta=16'h8c12;
13916: douta=16'h7bd1;
13917: douta=16'h8432;
13918: douta=16'h632e;
13919: douta=16'h6b0e;
13920: douta=16'h5aab;
13921: douta=16'h5aed;
13922: douta=16'h83f1;
13923: douta=16'h9472;
13924: douta=16'h9432;
13925: douta=16'h730e;
13926: douta=16'h7b8f;
13927: douta=16'h9d14;
13928: douta=16'hf7ff;
13929: douta=16'hffff;
13930: douta=16'hfe15;
13931: douta=16'hbb46;
13932: douta=16'hab66;
13933: douta=16'hb3c8;
13934: douta=16'hb3a8;
13935: douta=16'hb3c8;
13936: douta=16'hb3a8;
13937: douta=16'hb3a8;
13938: douta=16'haba8;
13939: douta=16'hb3c8;
13940: douta=16'hab88;
13941: douta=16'hb3c8;
13942: douta=16'hb3a8;
13943: douta=16'haba8;
13944: douta=16'hab88;
13945: douta=16'hab89;
13946: douta=16'haba9;
13947: douta=16'hab88;
13948: douta=16'hab88;
13949: douta=16'hab68;
13950: douta=16'ha368;
13951: douta=16'ha368;
13952: douta=16'h9c94;
13953: douta=16'h9cb4;
13954: douta=16'had15;
13955: douta=16'h8c96;
13956: douta=16'h28e3;
13957: douta=16'h28e3;
13958: douta=16'h28e3;
13959: douta=16'h28e3;
13960: douta=16'h28e3;
13961: douta=16'h20a3;
13962: douta=16'h2082;
13963: douta=16'h20c3;
13964: douta=16'h20a2;
13965: douta=16'h2082;
13966: douta=16'h20a2;
13967: douta=16'h20c2;
13968: douta=16'h28e2;
13969: douta=16'h30e2;
13970: douta=16'h3123;
13971: douta=16'h4143;
13972: douta=16'h4143;
13973: douta=16'h49a6;
13974: douta=16'h10e4;
13975: douta=16'h59c4;
13976: douta=16'h59c4;
13977: douta=16'h61e4;
13978: douta=16'h6a04;
13979: douta=16'h6a04;
13980: douta=16'h94b1;
13981: douta=16'h7a84;
13982: douta=16'h7a85;
13983: douta=16'h82a5;
13984: douta=16'h82a5;
13985: douta=16'h8ac6;
13986: douta=16'h8ac6;
13987: douta=16'h8ac6;
13988: douta=16'h7265;
13989: douta=16'h9306;
13990: douta=16'h9326;
13991: douta=16'h9326;
13992: douta=16'h9b26;
13993: douta=16'ha386;
13994: douta=16'hb3a7;
13995: douta=16'hb3c7;
13996: douta=16'hbbe7;
13997: douta=16'hbbe7;
13998: douta=16'hbc07;
13999: douta=16'hc407;
14000: douta=16'hc427;
14001: douta=16'hc427;
14002: douta=16'hc428;
14003: douta=16'hc428;
14004: douta=16'hc428;
14005: douta=16'hcc47;
14006: douta=16'hcc47;
14007: douta=16'hcc47;
14008: douta=16'hcc67;
14009: douta=16'hcc68;
14010: douta=16'hcc68;
14011: douta=16'hcc48;
14012: douta=16'hcc68;
14013: douta=16'hcc68;
14014: douta=16'hcc68;
14015: douta=16'hcc68;
14016: douta=16'hcc68;
14017: douta=16'hcc69;
14018: douta=16'hcc88;
14019: douta=16'hcc88;
14020: douta=16'hcc88;
14021: douta=16'hcc89;
14022: douta=16'hcc88;
14023: douta=16'hcc88;
14024: douta=16'hd488;
14025: douta=16'hd488;
14026: douta=16'hcc89;
14027: douta=16'hcc89;
14028: douta=16'hd489;
14029: douta=16'hcc88;
14030: douta=16'hd489;
14031: douta=16'hcc89;
14032: douta=16'hcc89;
14033: douta=16'had33;
14034: douta=16'hcc26;
14035: douta=16'hcc89;
14036: douta=16'hcc89;
14037: douta=16'hcc89;
14038: douta=16'hcc89;
14039: douta=16'hcc68;
14040: douta=16'hcc69;
14041: douta=16'hdc86;
14042: douta=16'h9431;
14043: douta=16'h7390;
14044: douta=16'h6b6f;
14045: douta=16'h6b4f;
14046: douta=16'h4a6b;
14047: douta=16'h62ee;
14048: douta=16'hacd4;
14049: douta=16'h7b90;
14050: douta=16'h62cd;
14051: douta=16'h8431;
14052: douta=16'hd71d;
14053: douta=16'hffff;
14054: douta=16'he5d3;
14055: douta=16'hcbc7;
14056: douta=16'hbba5;
14057: douta=16'hbc08;
14058: douta=16'hbbe8;
14059: douta=16'hb3c9;
14060: douta=16'hb3e9;
14061: douta=16'hbbc9;
14062: douta=16'hb3e9;
14063: douta=16'hb3c8;
14064: douta=16'hb3c8;
14065: douta=16'hb3a8;
14066: douta=16'hb3a8;
14067: douta=16'hb3a8;
14068: douta=16'hb3c8;
14069: douta=16'hb3c8;
14070: douta=16'hb3c8;
14071: douta=16'haba8;
14072: douta=16'hb3a8;
14073: douta=16'hab88;
14074: douta=16'hab88;
14075: douta=16'hab88;
14076: douta=16'hab89;
14077: douta=16'hab88;
14078: douta=16'hab88;
14079: douta=16'ha368;
14080: douta=16'h9cb4;
14081: douta=16'hb534;
14082: douta=16'h9cd6;
14083: douta=16'h8cd7;
14084: douta=16'h28e3;
14085: douta=16'h28e3;
14086: douta=16'h28e3;
14087: douta=16'h28e3;
14088: douta=16'h20c3;
14089: douta=16'h28e3;
14090: douta=16'h20a3;
14091: douta=16'h18a1;
14092: douta=16'h20a2;
14093: douta=16'h20c2;
14094: douta=16'h28c3;
14095: douta=16'h28e3;
14096: douta=16'h30e3;
14097: douta=16'h3103;
14098: douta=16'h3923;
14099: douta=16'h3943;
14100: douta=16'h4163;
14101: douta=16'h4a08;
14102: douta=16'h0884;
14103: douta=16'h51a4;
14104: douta=16'h61c4;
14105: douta=16'h6204;
14106: douta=16'h6a04;
14107: douta=16'h6a24;
14108: douta=16'had53;
14109: douta=16'h7a64;
14110: douta=16'h7a85;
14111: douta=16'h82a5;
14112: douta=16'h82a5;
14113: douta=16'h8ac6;
14114: douta=16'h8ac6;
14115: douta=16'h9307;
14116: douta=16'h7244;
14117: douta=16'h9326;
14118: douta=16'h9b47;
14119: douta=16'h9326;
14120: douta=16'h9b67;
14121: douta=16'hab87;
14122: douta=16'hb3c6;
14123: douta=16'hb3c7;
14124: douta=16'hbbe7;
14125: douta=16'hbbe7;
14126: douta=16'hbc07;
14127: douta=16'hbc07;
14128: douta=16'hc427;
14129: douta=16'hc428;
14130: douta=16'hc427;
14131: douta=16'hc448;
14132: douta=16'hc448;
14133: douta=16'hc448;
14134: douta=16'hc448;
14135: douta=16'hcc47;
14136: douta=16'hcc68;
14137: douta=16'hcc68;
14138: douta=16'hcc68;
14139: douta=16'hcc67;
14140: douta=16'hcc68;
14141: douta=16'hcc68;
14142: douta=16'hcc68;
14143: douta=16'hcc68;
14144: douta=16'hcc69;
14145: douta=16'hcc69;
14146: douta=16'hcc88;
14147: douta=16'hcc88;
14148: douta=16'hd4a9;
14149: douta=16'hcc89;
14150: douta=16'hcc89;
14151: douta=16'hcc89;
14152: douta=16'hd489;
14153: douta=16'hd489;
14154: douta=16'hcc89;
14155: douta=16'hcc89;
14156: douta=16'hcc89;
14157: douta=16'hd489;
14158: douta=16'hcc89;
14159: douta=16'hcc89;
14160: douta=16'hcc89;
14161: douta=16'had53;
14162: douta=16'hcc27;
14163: douta=16'hcc89;
14164: douta=16'hcc69;
14165: douta=16'hcc89;
14166: douta=16'hcc89;
14167: douta=16'hcc69;
14168: douta=16'hcc69;
14169: douta=16'hcc6a;
14170: douta=16'h8bef;
14171: douta=16'h528c;
14172: douta=16'h7bf1;
14173: douta=16'h9493;
14174: douta=16'h5acd;
14175: douta=16'h9d17;
14176: douta=16'hb6bf;
14177: douta=16'he7bf;
14178: douta=16'hd593;
14179: douta=16'hc3e7;
14180: douta=16'hc3e6;
14181: douta=16'hc428;
14182: douta=16'hc429;
14183: douta=16'hc429;
14184: douta=16'hbc09;
14185: douta=16'hbc09;
14186: douta=16'hbc08;
14187: douta=16'hbc09;
14188: douta=16'hbbe9;
14189: douta=16'hbbe9;
14190: douta=16'hbbe9;
14191: douta=16'hb3e8;
14192: douta=16'hb3e9;
14193: douta=16'hb3c9;
14194: douta=16'hb3c9;
14195: douta=16'hb3a8;
14196: douta=16'hb3a9;
14197: douta=16'hb3c8;
14198: douta=16'hb3c8;
14199: douta=16'hb3c8;
14200: douta=16'hb3a8;
14201: douta=16'haba9;
14202: douta=16'hab88;
14203: douta=16'ha388;
14204: douta=16'hab89;
14205: douta=16'hab89;
14206: douta=16'ha368;
14207: douta=16'ha388;
14208: douta=16'ha4f5;
14209: douta=16'hbd75;
14210: douta=16'h8c95;
14211: douta=16'h7c53;
14212: douta=16'h28e3;
14213: douta=16'h28e3;
14214: douta=16'h28e3;
14215: douta=16'h28e3;
14216: douta=16'h20c3;
14217: douta=16'h20c3;
14218: douta=16'h20c3;
14219: douta=16'h20a2;
14220: douta=16'h20a2;
14221: douta=16'h20c2;
14222: douta=16'h28c3;
14223: douta=16'h28e3;
14224: douta=16'h28e2;
14225: douta=16'h3103;
14226: douta=16'h3923;
14227: douta=16'h4144;
14228: douta=16'h4984;
14229: douta=16'h528b;
14230: douta=16'h18c4;
14231: douta=16'h59c4;
14232: douta=16'h61e4;
14233: douta=16'h6204;
14234: douta=16'h6a25;
14235: douta=16'h7203;
14236: douta=16'haccf;
14237: douta=16'h7a84;
14238: douta=16'h8285;
14239: douta=16'h8aa6;
14240: douta=16'h8aa5;
14241: douta=16'h8ac6;
14242: douta=16'h8ac6;
14243: douta=16'h9307;
14244: douta=16'h82a6;
14245: douta=16'h9b47;
14246: douta=16'h9b47;
14247: douta=16'h9326;
14248: douta=16'ha367;
14249: douta=16'hab86;
14250: douta=16'hb3c7;
14251: douta=16'hb3c7;
14252: douta=16'hbbe7;
14253: douta=16'hbbe7;
14254: douta=16'hbc07;
14255: douta=16'hbc07;
14256: douta=16'hc428;
14257: douta=16'hc427;
14258: douta=16'hc428;
14259: douta=16'hc448;
14260: douta=16'hcc48;
14261: douta=16'hc447;
14262: douta=16'hcc48;
14263: douta=16'hcc67;
14264: douta=16'hcc68;
14265: douta=16'hcc68;
14266: douta=16'hcc68;
14267: douta=16'hcc68;
14268: douta=16'hcc68;
14269: douta=16'hcc68;
14270: douta=16'hcc68;
14271: douta=16'hcc68;
14272: douta=16'hcc68;
14273: douta=16'hcc68;
14274: douta=16'hcc89;
14275: douta=16'hd489;
14276: douta=16'hcc89;
14277: douta=16'hd489;
14278: douta=16'hcc89;
14279: douta=16'hd48a;
14280: douta=16'hd489;
14281: douta=16'hd489;
14282: douta=16'hcc89;
14283: douta=16'hcc69;
14284: douta=16'hd48a;
14285: douta=16'hcc89;
14286: douta=16'hcc89;
14287: douta=16'hcc89;
14288: douta=16'hcc69;
14289: douta=16'had33;
14290: douta=16'hcc47;
14291: douta=16'hcc89;
14292: douta=16'hcc69;
14293: douta=16'hcc69;
14294: douta=16'hcc89;
14295: douta=16'hcc69;
14296: douta=16'hcc69;
14297: douta=16'hcc69;
14298: douta=16'hcc69;
14299: douta=16'hc449;
14300: douta=16'hcc49;
14301: douta=16'hd485;
14302: douta=16'hd618;
14303: douta=16'hc428;
14304: douta=16'hc448;
14305: douta=16'hcc4a;
14306: douta=16'hcc49;
14307: douta=16'hc448;
14308: douta=16'hc428;
14309: douta=16'hc449;
14310: douta=16'hc429;
14311: douta=16'hbc08;
14312: douta=16'hc429;
14313: douta=16'hbc09;
14314: douta=16'hbc09;
14315: douta=16'hbc09;
14316: douta=16'hbc09;
14317: douta=16'hbbe9;
14318: douta=16'hb3c8;
14319: douta=16'hb3e9;
14320: douta=16'hb3c9;
14321: douta=16'hb3c8;
14322: douta=16'hb3c8;
14323: douta=16'hb3c8;
14324: douta=16'hb3c8;
14325: douta=16'hb3c8;
14326: douta=16'hb3c8;
14327: douta=16'hb3a8;
14328: douta=16'hab89;
14329: douta=16'haba9;
14330: douta=16'haba9;
14331: douta=16'haba8;
14332: douta=16'haba8;
14333: douta=16'ha388;
14334: douta=16'ha389;
14335: douta=16'ha389;
14336: douta=16'ha4d5;
14337: douta=16'ha515;
14338: douta=16'h94b6;
14339: douta=16'h3186;
14340: douta=16'h28e3;
14341: douta=16'h28e3;
14342: douta=16'h28e3;
14343: douta=16'h28e3;
14344: douta=16'h28e3;
14345: douta=16'h20a3;
14346: douta=16'h20e3;
14347: douta=16'h20a2;
14348: douta=16'h20c2;
14349: douta=16'h20a2;
14350: douta=16'h28e3;
14351: douta=16'h30e3;
14352: douta=16'h30e3;
14353: douta=16'h3103;
14354: douta=16'h3923;
14355: douta=16'h4144;
14356: douta=16'h4963;
14357: douta=16'h4a49;
14358: douta=16'h3924;
14359: douta=16'h59c4;
14360: douta=16'h61e4;
14361: douta=16'h6a24;
14362: douta=16'h6a24;
14363: douta=16'h7245;
14364: douta=16'h93aa;
14365: douta=16'h7a85;
14366: douta=16'h7a85;
14367: douta=16'h8aa6;
14368: douta=16'h8ac6;
14369: douta=16'h8ac6;
14370: douta=16'h8ac6;
14371: douta=16'h9306;
14372: douta=16'h9b47;
14373: douta=16'ha347;
14374: douta=16'h9b47;
14375: douta=16'h9b47;
14376: douta=16'ha367;
14377: douta=16'haba7;
14378: douta=16'hb3c7;
14379: douta=16'hbbe7;
14380: douta=16'hbbe7;
14381: douta=16'hbbe7;
14382: douta=16'hbc07;
14383: douta=16'hc407;
14384: douta=16'hc428;
14385: douta=16'hc428;
14386: douta=16'hc428;
14387: douta=16'hc448;
14388: douta=16'hcc67;
14389: douta=16'hcc47;
14390: douta=16'hcc48;
14391: douta=16'hcc68;
14392: douta=16'hcc68;
14393: douta=16'hcc68;
14394: douta=16'hcc68;
14395: douta=16'hcc68;
14396: douta=16'hcc68;
14397: douta=16'hcc88;
14398: douta=16'hcc88;
14399: douta=16'hcc68;
14400: douta=16'hcc88;
14401: douta=16'hcc68;
14402: douta=16'hcc69;
14403: douta=16'hcc69;
14404: douta=16'hcc89;
14405: douta=16'hcc89;
14406: douta=16'hcc69;
14407: douta=16'hcc69;
14408: douta=16'hcc89;
14409: douta=16'hcc89;
14410: douta=16'hd489;
14411: douta=16'hcc69;
14412: douta=16'hd48a;
14413: douta=16'hcc89;
14414: douta=16'hcc89;
14415: douta=16'hcc69;
14416: douta=16'hcc89;
14417: douta=16'had53;
14418: douta=16'hcc27;
14419: douta=16'hcc69;
14420: douta=16'hcc89;
14421: douta=16'hcc69;
14422: douta=16'hcc69;
14423: douta=16'hcc69;
14424: douta=16'hcc69;
14425: douta=16'hcc49;
14426: douta=16'hcc69;
14427: douta=16'hcc49;
14428: douta=16'hcc69;
14429: douta=16'hcc69;
14430: douta=16'hcc69;
14431: douta=16'hcc49;
14432: douta=16'hc449;
14433: douta=16'hcc49;
14434: douta=16'hcc49;
14435: douta=16'hc428;
14436: douta=16'hc449;
14437: douta=16'hc429;
14438: douta=16'hc429;
14439: douta=16'hc429;
14440: douta=16'hc429;
14441: douta=16'hc429;
14442: douta=16'hbc09;
14443: douta=16'hbc09;
14444: douta=16'hbc09;
14445: douta=16'hb3e8;
14446: douta=16'hbbe9;
14447: douta=16'hbbe9;
14448: douta=16'hb3e9;
14449: douta=16'hb3c8;
14450: douta=16'hb3c8;
14451: douta=16'hb3c8;
14452: douta=16'hb3c8;
14453: douta=16'hb3c9;
14454: douta=16'hb3c8;
14455: douta=16'hb3a9;
14456: douta=16'haba9;
14457: douta=16'haba9;
14458: douta=16'habc9;
14459: douta=16'hab88;
14460: douta=16'hab89;
14461: douta=16'ha368;
14462: douta=16'ha389;
14463: douta=16'ha388;
14464: douta=16'ha4f5;
14465: douta=16'h8c95;
14466: douta=16'h8c96;
14467: douta=16'h2082;
14468: douta=16'h28e3;
14469: douta=16'h28e3;
14470: douta=16'h28e3;
14471: douta=16'h28e3;
14472: douta=16'h28e3;
14473: douta=16'h20c3;
14474: douta=16'h20e3;
14475: douta=16'h20c2;
14476: douta=16'h20a2;
14477: douta=16'h28c3;
14478: douta=16'h28e3;
14479: douta=16'h28e2;
14480: douta=16'h30e3;
14481: douta=16'h3103;
14482: douta=16'h4123;
14483: douta=16'h4143;
14484: douta=16'h4963;
14485: douta=16'h31a7;
14486: douta=16'h5184;
14487: douta=16'h59c4;
14488: douta=16'h6204;
14489: douta=16'h6204;
14490: douta=16'h6a24;
14491: douta=16'h6a46;
14492: douta=16'h7245;
14493: douta=16'h7a85;
14494: douta=16'h8285;
14495: douta=16'h8aa6;
14496: douta=16'h8ac6;
14497: douta=16'h8ac6;
14498: douta=16'h92e7;
14499: douta=16'h9306;
14500: douta=16'h9b47;
14501: douta=16'h7265;
14502: douta=16'h8a82;
14503: douta=16'h7a23;
14504: douta=16'h8aa2;
14505: douta=16'haba6;
14506: douta=16'hb3c7;
14507: douta=16'hb3e7;
14508: douta=16'hbbe7;
14509: douta=16'hbc07;
14510: douta=16'hbc08;
14511: douta=16'hc428;
14512: douta=16'hc428;
14513: douta=16'hc427;
14514: douta=16'hc428;
14515: douta=16'hc448;
14516: douta=16'hc448;
14517: douta=16'hc448;
14518: douta=16'hcc48;
14519: douta=16'hcc68;
14520: douta=16'hcc68;
14521: douta=16'hcc68;
14522: douta=16'hcc68;
14523: douta=16'hcc68;
14524: douta=16'hcc68;
14525: douta=16'hcc68;
14526: douta=16'hcc68;
14527: douta=16'hcc68;
14528: douta=16'hcc69;
14529: douta=16'hcc89;
14530: douta=16'hcc89;
14531: douta=16'hcc89;
14532: douta=16'hcc89;
14533: douta=16'hcc89;
14534: douta=16'hcc69;
14535: douta=16'hcc89;
14536: douta=16'hcc69;
14537: douta=16'hcc69;
14538: douta=16'hd489;
14539: douta=16'hcc89;
14540: douta=16'hd48a;
14541: douta=16'hcc69;
14542: douta=16'hcc89;
14543: douta=16'hcc89;
14544: douta=16'hcc89;
14545: douta=16'had73;
14546: douta=16'hcc47;
14547: douta=16'hcc69;
14548: douta=16'hcc69;
14549: douta=16'hcc69;
14550: douta=16'hcc69;
14551: douta=16'hcc69;
14552: douta=16'hcc69;
14553: douta=16'hcc69;
14554: douta=16'hcc69;
14555: douta=16'hcc69;
14556: douta=16'hcc69;
14557: douta=16'hcc69;
14558: douta=16'hcc69;
14559: douta=16'hcc69;
14560: douta=16'hc449;
14561: douta=16'hcc49;
14562: douta=16'hc449;
14563: douta=16'hc449;
14564: douta=16'hc449;
14565: douta=16'hc429;
14566: douta=16'hc429;
14567: douta=16'hc429;
14568: douta=16'hbc08;
14569: douta=16'hbc09;
14570: douta=16'hbc09;
14571: douta=16'hbc09;
14572: douta=16'hbc09;
14573: douta=16'hbbe9;
14574: douta=16'hbbe9;
14575: douta=16'hbbe9;
14576: douta=16'hbbe9;
14577: douta=16'hb3e9;
14578: douta=16'hb3c9;
14579: douta=16'hb3c8;
14580: douta=16'hb3c9;
14581: douta=16'hb3c8;
14582: douta=16'hb3c8;
14583: douta=16'haba9;
14584: douta=16'haba8;
14585: douta=16'haba9;
14586: douta=16'haba9;
14587: douta=16'hab88;
14588: douta=16'hab88;
14589: douta=16'ha389;
14590: douta=16'hab89;
14591: douta=16'ha368;
14592: douta=16'h94b4;
14593: douta=16'h94d6;
14594: douta=16'h8475;
14595: douta=16'h2904;
14596: douta=16'h2904;
14597: douta=16'h28e3;
14598: douta=16'h28e3;
14599: douta=16'h28e3;
14600: douta=16'h20e3;
14601: douta=16'h20e3;
14602: douta=16'h20a2;
14603: douta=16'h20a2;
14604: douta=16'h20c2;
14605: douta=16'h20c2;
14606: douta=16'h28e3;
14607: douta=16'h28e2;
14608: douta=16'h30e2;
14609: douta=16'h3103;
14610: douta=16'h4124;
14611: douta=16'h4163;
14612: douta=16'h4984;
14613: douta=16'h1905;
14614: douta=16'h61c3;
14615: douta=16'h59c4;
14616: douta=16'h6204;
14617: douta=16'h6a04;
14618: douta=16'h7224;
14619: douta=16'h7b6c;
14620: douta=16'h7223;
14621: douta=16'h7a85;
14622: douta=16'h82a5;
14623: douta=16'h82a6;
14624: douta=16'h8ac6;
14625: douta=16'h8ae7;
14626: douta=16'h8ac6;
14627: douta=16'h9306;
14628: douta=16'h9326;
14629: douta=16'h6a24;
14630: douta=16'hde97;
14631: douta=16'hd635;
14632: douta=16'hde97;
14633: douta=16'hb3e7;
14634: douta=16'hb3c7;
14635: douta=16'hb3e7;
14636: douta=16'hbbe7;
14637: douta=16'hbc07;
14638: douta=16'hbc07;
14639: douta=16'hbc07;
14640: douta=16'hc428;
14641: douta=16'hc428;
14642: douta=16'hc448;
14643: douta=16'hc448;
14644: douta=16'hc448;
14645: douta=16'hc448;
14646: douta=16'hcc49;
14647: douta=16'hc448;
14648: douta=16'hcc68;
14649: douta=16'hcc68;
14650: douta=16'hcc68;
14651: douta=16'hcc68;
14652: douta=16'hcc68;
14653: douta=16'hcc68;
14654: douta=16'hcc68;
14655: douta=16'hcc89;
14656: douta=16'hcc89;
14657: douta=16'hcc69;
14658: douta=16'hcc69;
14659: douta=16'hcc89;
14660: douta=16'hcc89;
14661: douta=16'hcc89;
14662: douta=16'hcc89;
14663: douta=16'hcc89;
14664: douta=16'hcc89;
14665: douta=16'hcc8a;
14666: douta=16'hcc89;
14667: douta=16'hd48a;
14668: douta=16'hcc8a;
14669: douta=16'hcc89;
14670: douta=16'hcc89;
14671: douta=16'hcc89;
14672: douta=16'hcc89;
14673: douta=16'had73;
14674: douta=16'hcc47;
14675: douta=16'hcc69;
14676: douta=16'hcc89;
14677: douta=16'hcc69;
14678: douta=16'hcc69;
14679: douta=16'hcc69;
14680: douta=16'hcc69;
14681: douta=16'hcc69;
14682: douta=16'hcc69;
14683: douta=16'hcc69;
14684: douta=16'hcc69;
14685: douta=16'hcc69;
14686: douta=16'hcc69;
14687: douta=16'hc448;
14688: douta=16'hcc69;
14689: douta=16'hc449;
14690: douta=16'hc449;
14691: douta=16'hc449;
14692: douta=16'hc429;
14693: douta=16'hc429;
14694: douta=16'hbc09;
14695: douta=16'hc429;
14696: douta=16'hc429;
14697: douta=16'hbc29;
14698: douta=16'hbc29;
14699: douta=16'hbc09;
14700: douta=16'hbc09;
14701: douta=16'hbc09;
14702: douta=16'hbbe9;
14703: douta=16'hbbe9;
14704: douta=16'hbbe9;
14705: douta=16'hb3e9;
14706: douta=16'hb3c8;
14707: douta=16'hb3e9;
14708: douta=16'hb3c9;
14709: douta=16'hb3c9;
14710: douta=16'hb3c9;
14711: douta=16'habc9;
14712: douta=16'haba9;
14713: douta=16'haba8;
14714: douta=16'haba9;
14715: douta=16'haba9;
14716: douta=16'hab89;
14717: douta=16'hab89;
14718: douta=16'ha388;
14719: douta=16'ha368;
14720: douta=16'h8c95;
14721: douta=16'h94f7;
14722: douta=16'h2924;
14723: douta=16'h28e3;
14724: douta=16'h3124;
14725: douta=16'h28e3;
14726: douta=16'h28e3;
14727: douta=16'h28e3;
14728: douta=16'h20c3;
14729: douta=16'h20e3;
14730: douta=16'h20a2;
14731: douta=16'h20c2;
14732: douta=16'h20c2;
14733: douta=16'h28e3;
14734: douta=16'h28e3;
14735: douta=16'h28e3;
14736: douta=16'h3103;
14737: douta=16'h3123;
14738: douta=16'h4124;
14739: douta=16'h4963;
14740: douta=16'h49c7;
14741: douta=16'h0884;
14742: douta=16'h59c4;
14743: douta=16'h59c4;
14744: douta=16'h6204;
14745: douta=16'h6a24;
14746: douta=16'h7224;
14747: douta=16'h9cd1;
14748: douta=16'h7a64;
14749: douta=16'h7a85;
14750: douta=16'h82a5;
14751: douta=16'h82c6;
14752: douta=16'h8ac6;
14753: douta=16'h8ae6;
14754: douta=16'h9307;
14755: douta=16'h9306;
14756: douta=16'h9b27;
14757: douta=16'h8aa5;
14758: douta=16'h2985;
14759: douta=16'h0000;
14760: douta=16'had52;
14761: douta=16'hb3c7;
14762: douta=16'haba7;
14763: douta=16'hb3e7;
14764: douta=16'hbbe7;
14765: douta=16'hbc07;
14766: douta=16'hbc07;
14767: douta=16'hc428;
14768: douta=16'hc428;
14769: douta=16'hc428;
14770: douta=16'hc448;
14771: douta=16'hc448;
14772: douta=16'hcc68;
14773: douta=16'hcc49;
14774: douta=16'hcc49;
14775: douta=16'hcc68;
14776: douta=16'hcc68;
14777: douta=16'hcc68;
14778: douta=16'hcc68;
14779: douta=16'hcc68;
14780: douta=16'hcc68;
14781: douta=16'hcc68;
14782: douta=16'hcc69;
14783: douta=16'hcc69;
14784: douta=16'hcc68;
14785: douta=16'hcc89;
14786: douta=16'hcc89;
14787: douta=16'hcc8a;
14788: douta=16'hcc89;
14789: douta=16'hcc89;
14790: douta=16'hcc89;
14791: douta=16'hcc89;
14792: douta=16'hcc89;
14793: douta=16'hcc8a;
14794: douta=16'hcc69;
14795: douta=16'hcc89;
14796: douta=16'hcc89;
14797: douta=16'hcc89;
14798: douta=16'hcc89;
14799: douta=16'hcc89;
14800: douta=16'hcc89;
14801: douta=16'hb594;
14802: douta=16'hcc47;
14803: douta=16'hcc69;
14804: douta=16'hcc69;
14805: douta=16'hcc69;
14806: douta=16'hcc69;
14807: douta=16'hcc89;
14808: douta=16'hcc89;
14809: douta=16'hcc69;
14810: douta=16'hcc69;
14811: douta=16'hcc69;
14812: douta=16'hcc49;
14813: douta=16'hcc69;
14814: douta=16'hcc69;
14815: douta=16'hcc49;
14816: douta=16'hc449;
14817: douta=16'hc449;
14818: douta=16'hc449;
14819: douta=16'hc429;
14820: douta=16'hc429;
14821: douta=16'hc449;
14822: douta=16'hc449;
14823: douta=16'hc429;
14824: douta=16'hc429;
14825: douta=16'hbc29;
14826: douta=16'hc429;
14827: douta=16'hbc09;
14828: douta=16'hbbe9;
14829: douta=16'hbc09;
14830: douta=16'hbbe9;
14831: douta=16'hb3e9;
14832: douta=16'hb3e9;
14833: douta=16'hbc09;
14834: douta=16'hb3c9;
14835: douta=16'hb3e9;
14836: douta=16'hb3c9;
14837: douta=16'hb3c9;
14838: douta=16'hb3c9;
14839: douta=16'haba9;
14840: douta=16'haba9;
14841: douta=16'haba9;
14842: douta=16'haba9;
14843: douta=16'haba8;
14844: douta=16'haba9;
14845: douta=16'haba9;
14846: douta=16'ha389;
14847: douta=16'ha389;
14848: douta=16'h94b6;
14849: douta=16'h8496;
14850: douta=16'h2082;
14851: douta=16'h28e3;
14852: douta=16'h28e3;
14853: douta=16'h28e3;
14854: douta=16'h28e3;
14855: douta=16'h20e3;
14856: douta=16'h20e3;
14857: douta=16'h20e3;
14858: douta=16'h20a2;
14859: douta=16'h20c2;
14860: douta=16'h28c3;
14861: douta=16'h28e3;
14862: douta=16'h3103;
14863: douta=16'h30e3;
14864: douta=16'h3103;
14865: douta=16'h3923;
14866: douta=16'h4143;
14867: douta=16'h4964;
14868: douta=16'h524a;
14869: douta=16'h1084;
14870: douta=16'h61c4;
14871: douta=16'h59c4;
14872: douta=16'h6204;
14873: douta=16'h6a24;
14874: douta=16'h7224;
14875: douta=16'hb593;
14876: douta=16'h7a64;
14877: douta=16'h7a85;
14878: douta=16'h82a5;
14879: douta=16'h82c6;
14880: douta=16'h8ae7;
14881: douta=16'h8ae7;
14882: douta=16'h9307;
14883: douta=16'h9326;
14884: douta=16'h9b47;
14885: douta=16'h9b46;
14886: douta=16'h8caf;
14887: douta=16'h7b8a;
14888: douta=16'h7bad;
14889: douta=16'hb3c7;
14890: douta=16'hb3c8;
14891: douta=16'hbc08;
14892: douta=16'hbc07;
14893: douta=16'hbc07;
14894: douta=16'hbc07;
14895: douta=16'hc428;
14896: douta=16'hc428;
14897: douta=16'hc428;
14898: douta=16'hc448;
14899: douta=16'hc428;
14900: douta=16'hc448;
14901: douta=16'hc448;
14902: douta=16'hcc68;
14903: douta=16'hc448;
14904: douta=16'hcc68;
14905: douta=16'hcc68;
14906: douta=16'hcc68;
14907: douta=16'hcc69;
14908: douta=16'hcc68;
14909: douta=16'hcc89;
14910: douta=16'hcc69;
14911: douta=16'hcc69;
14912: douta=16'hcc69;
14913: douta=16'hcc69;
14914: douta=16'hcc69;
14915: douta=16'hcc89;
14916: douta=16'hcc89;
14917: douta=16'hcc89;
14918: douta=16'hcc89;
14919: douta=16'hcc89;
14920: douta=16'hcc89;
14921: douta=16'hcc89;
14922: douta=16'hcc89;
14923: douta=16'hcc89;
14924: douta=16'hcc89;
14925: douta=16'hcc89;
14926: douta=16'hcc69;
14927: douta=16'hcc69;
14928: douta=16'hcc69;
14929: douta=16'hb594;
14930: douta=16'hcc48;
14931: douta=16'hcc69;
14932: douta=16'hcc69;
14933: douta=16'hcc69;
14934: douta=16'hcc69;
14935: douta=16'hcc69;
14936: douta=16'hcc69;
14937: douta=16'hcc69;
14938: douta=16'hcc49;
14939: douta=16'hcc69;
14940: douta=16'hcc49;
14941: douta=16'hcc49;
14942: douta=16'hcc49;
14943: douta=16'hcc69;
14944: douta=16'hcc69;
14945: douta=16'hc449;
14946: douta=16'hc449;
14947: douta=16'hc429;
14948: douta=16'hc429;
14949: douta=16'hc429;
14950: douta=16'hbc29;
14951: douta=16'hc429;
14952: douta=16'hc429;
14953: douta=16'hbc29;
14954: douta=16'hbc09;
14955: douta=16'hbc29;
14956: douta=16'hbc09;
14957: douta=16'hbc09;
14958: douta=16'hbc09;
14959: douta=16'hbbe9;
14960: douta=16'hbbe9;
14961: douta=16'hb3e9;
14962: douta=16'hb3c9;
14963: douta=16'hb3c9;
14964: douta=16'hb3e9;
14965: douta=16'hb3c9;
14966: douta=16'hb3c9;
14967: douta=16'hb3c9;
14968: douta=16'haba9;
14969: douta=16'haba9;
14970: douta=16'haba9;
14971: douta=16'haba9;
14972: douta=16'haba9;
14973: douta=16'ha389;
14974: douta=16'ha389;
14975: douta=16'ha389;
14976: douta=16'h94b5;
14977: douta=16'h9518;
14978: douta=16'h2903;
14979: douta=16'h28e3;
14980: douta=16'h28e3;
14981: douta=16'h28e3;
14982: douta=16'h20e3;
14983: douta=16'h20e3;
14984: douta=16'h20e3;
14985: douta=16'h28e3;
14986: douta=16'h20c3;
14987: douta=16'h20c3;
14988: douta=16'h28c3;
14989: douta=16'h28e3;
14990: douta=16'h3103;
14991: douta=16'h3103;
14992: douta=16'h3103;
14993: douta=16'h3923;
14994: douta=16'h4143;
14995: douta=16'h4964;
14996: douta=16'h528b;
14997: douta=16'h3104;
14998: douta=16'h59c4;
14999: douta=16'h61e4;
15000: douta=16'h6a24;
15001: douta=16'h7245;
15002: douta=16'h7223;
15003: douta=16'hacf0;
15004: douta=16'h7a85;
15005: douta=16'h7a85;
15006: douta=16'h82a6;
15007: douta=16'h82c6;
15008: douta=16'h8ac6;
15009: douta=16'h8ae6;
15010: douta=16'h9307;
15011: douta=16'h9b27;
15012: douta=16'h9b47;
15013: douta=16'hac4b;
15014: douta=16'hacb0;
15015: douta=16'hb44e;
15016: douta=16'h5a47;
15017: douta=16'haba7;
15018: douta=16'hb3c7;
15019: douta=16'hbbe8;
15020: douta=16'hbbe7;
15021: douta=16'hbc08;
15022: douta=16'hc407;
15023: douta=16'hc407;
15024: douta=16'hc448;
15025: douta=16'hc448;
15026: douta=16'hc448;
15027: douta=16'hcc49;
15028: douta=16'hc428;
15029: douta=16'hc449;
15030: douta=16'hcc49;
15031: douta=16'hc448;
15032: douta=16'hcc68;
15033: douta=16'hcc68;
15034: douta=16'hcc68;
15035: douta=16'hcc68;
15036: douta=16'hcc68;
15037: douta=16'hcc69;
15038: douta=16'hcc69;
15039: douta=16'hcc69;
15040: douta=16'hcc69;
15041: douta=16'hcc69;
15042: douta=16'hcc89;
15043: douta=16'hcc89;
15044: douta=16'hcc89;
15045: douta=16'hcc89;
15046: douta=16'hcc89;
15047: douta=16'hcc89;
15048: douta=16'hcc89;
15049: douta=16'hcc69;
15050: douta=16'hcc89;
15051: douta=16'hcc89;
15052: douta=16'hcc89;
15053: douta=16'hcc69;
15054: douta=16'hcc89;
15055: douta=16'hcc69;
15056: douta=16'hcc69;
15057: douta=16'hb594;
15058: douta=16'hcc48;
15059: douta=16'hcc69;
15060: douta=16'hcc69;
15061: douta=16'hcc69;
15062: douta=16'hcc69;
15063: douta=16'hcc69;
15064: douta=16'hcc69;
15065: douta=16'hcc69;
15066: douta=16'hcc8a;
15067: douta=16'hcc69;
15068: douta=16'hc449;
15069: douta=16'hcc69;
15070: douta=16'hc449;
15071: douta=16'hc449;
15072: douta=16'hc449;
15073: douta=16'hc449;
15074: douta=16'hc429;
15075: douta=16'hc429;
15076: douta=16'hc429;
15077: douta=16'hc429;
15078: douta=16'hc429;
15079: douta=16'hc429;
15080: douta=16'hc429;
15081: douta=16'hbc29;
15082: douta=16'hbc29;
15083: douta=16'hbc09;
15084: douta=16'hbc2a;
15085: douta=16'hbc09;
15086: douta=16'hbc09;
15087: douta=16'hbc09;
15088: douta=16'hbc09;
15089: douta=16'hbbe9;
15090: douta=16'hb3e9;
15091: douta=16'hb3e9;
15092: douta=16'hb3e9;
15093: douta=16'hb3c9;
15094: douta=16'habc9;
15095: douta=16'haba9;
15096: douta=16'habc9;
15097: douta=16'haba9;
15098: douta=16'haba9;
15099: douta=16'haba9;
15100: douta=16'haba9;
15101: douta=16'haba9;
15102: douta=16'ha389;
15103: douta=16'ha389;
15104: douta=16'h8cb6;
15105: douta=16'h528c;
15106: douta=16'h2904;
15107: douta=16'h2904;
15108: douta=16'h20e3;
15109: douta=16'h2904;
15110: douta=16'h28e3;
15111: douta=16'h2904;
15112: douta=16'h20e3;
15113: douta=16'h20e3;
15114: douta=16'h20a3;
15115: douta=16'h28e3;
15116: douta=16'h28e3;
15117: douta=16'h28e3;
15118: douta=16'h30e3;
15119: douta=16'h3103;
15120: douta=16'h3123;
15121: douta=16'h3943;
15122: douta=16'h4144;
15123: douta=16'h4964;
15124: douta=16'h4249;
15125: douta=16'h4984;
15126: douta=16'h59c4;
15127: douta=16'h61e4;
15128: douta=16'h6a24;
15129: douta=16'h7245;
15130: douta=16'h7224;
15131: douta=16'h93eb;
15132: douta=16'h7a85;
15133: douta=16'h8285;
15134: douta=16'h82c6;
15135: douta=16'h82c6;
15136: douta=16'h8ae7;
15137: douta=16'h8ae7;
15138: douta=16'h9307;
15139: douta=16'h9b27;
15140: douta=16'h9b27;
15141: douta=16'hcd52;
15142: douta=16'h0000;
15143: douta=16'hcdb3;
15144: douta=16'h59a4;
15145: douta=16'haba7;
15146: douta=16'hb3c7;
15147: douta=16'hb3c7;
15148: douta=16'hbc08;
15149: douta=16'hbc08;
15150: douta=16'hbc08;
15151: douta=16'hc428;
15152: douta=16'hc428;
15153: douta=16'hc448;
15154: douta=16'hcc49;
15155: douta=16'hc428;
15156: douta=16'hc448;
15157: douta=16'hc449;
15158: douta=16'hc448;
15159: douta=16'hc448;
15160: douta=16'hcc69;
15161: douta=16'hcc49;
15162: douta=16'hcc68;
15163: douta=16'hcc69;
15164: douta=16'hcc69;
15165: douta=16'hcc69;
15166: douta=16'hcc69;
15167: douta=16'hcc89;
15168: douta=16'hcc89;
15169: douta=16'hcc69;
15170: douta=16'hcc89;
15171: douta=16'hcc89;
15172: douta=16'hcc89;
15173: douta=16'hcc89;
15174: douta=16'hcc89;
15175: douta=16'hcc69;
15176: douta=16'hcc89;
15177: douta=16'hcc89;
15178: douta=16'hcc89;
15179: douta=16'hcc89;
15180: douta=16'hcc89;
15181: douta=16'hcc69;
15182: douta=16'hcc69;
15183: douta=16'hcc89;
15184: douta=16'hcc69;
15185: douta=16'hb5b5;
15186: douta=16'hcc48;
15187: douta=16'hcc69;
15188: douta=16'hcc6a;
15189: douta=16'hcc69;
15190: douta=16'hcc69;
15191: douta=16'hcc69;
15192: douta=16'hcc6a;
15193: douta=16'hcc69;
15194: douta=16'hcc69;
15195: douta=16'hcc49;
15196: douta=16'hc449;
15197: douta=16'hcc49;
15198: douta=16'hcc49;
15199: douta=16'hc449;
15200: douta=16'hc429;
15201: douta=16'hc449;
15202: douta=16'hc429;
15203: douta=16'hc429;
15204: douta=16'hc429;
15205: douta=16'hbc29;
15206: douta=16'hc429;
15207: douta=16'hc429;
15208: douta=16'hc429;
15209: douta=16'hbc29;
15210: douta=16'hbc09;
15211: douta=16'hbc2a;
15212: douta=16'hbc09;
15213: douta=16'hbc09;
15214: douta=16'hbc09;
15215: douta=16'hbc09;
15216: douta=16'hbbe9;
15217: douta=16'hbc09;
15218: douta=16'hb3c9;
15219: douta=16'hbbe9;
15220: douta=16'hb3e9;
15221: douta=16'hb3e9;
15222: douta=16'habc9;
15223: douta=16'hb3c9;
15224: douta=16'haba9;
15225: douta=16'habc9;
15226: douta=16'haba9;
15227: douta=16'haba8;
15228: douta=16'hab89;
15229: douta=16'ha388;
15230: douta=16'ha389;
15231: douta=16'ha389;
15232: douta=16'h84b7;
15233: douta=16'h1861;
15234: douta=16'h2904;
15235: douta=16'h20e3;
15236: douta=16'h28e3;
15237: douta=16'h2904;
15238: douta=16'h2904;
15239: douta=16'h20e3;
15240: douta=16'h20e3;
15241: douta=16'h20a3;
15242: douta=16'h20c2;
15243: douta=16'h20c2;
15244: douta=16'h28e3;
15245: douta=16'h28e3;
15246: douta=16'h30e3;
15247: douta=16'h3103;
15248: douta=16'h3923;
15249: douta=16'h3944;
15250: douta=16'h4164;
15251: douta=16'h4964;
15252: douta=16'h2947;
15253: douta=16'h6204;
15254: douta=16'h59c4;
15255: douta=16'h6204;
15256: douta=16'h6a25;
15257: douta=16'h6a44;
15258: douta=16'h7288;
15259: douta=16'h7a85;
15260: douta=16'h7a85;
15261: douta=16'h82a5;
15262: douta=16'h82c6;
15263: douta=16'h82c6;
15264: douta=16'h8ae7;
15265: douta=16'h8b07;
15266: douta=16'h8b07;
15267: douta=16'h9b47;
15268: douta=16'h9b27;
15269: douta=16'hde77;
15270: douta=16'he6b7;
15271: douta=16'hde76;
15272: douta=16'h7a23;
15273: douta=16'habc8;
15274: douta=16'hb3c7;
15275: douta=16'hb3e8;
15276: douta=16'hbc08;
15277: douta=16'hbc08;
15278: douta=16'hc408;
15279: douta=16'hc428;
15280: douta=16'hc448;
15281: douta=16'hc448;
15282: douta=16'hc428;
15283: douta=16'hc448;
15284: douta=16'hc448;
15285: douta=16'hc448;
15286: douta=16'hc449;
15287: douta=16'hc448;
15288: douta=16'hcc49;
15289: douta=16'hcc69;
15290: douta=16'hcc69;
15291: douta=16'hcc68;
15292: douta=16'hcc69;
15293: douta=16'hcc89;
15294: douta=16'hcc69;
15295: douta=16'hcc69;
15296: douta=16'hcc69;
15297: douta=16'hcc69;
15298: douta=16'hcc89;
15299: douta=16'hcc69;
15300: douta=16'hcc89;
15301: douta=16'hcc69;
15302: douta=16'hcc89;
15303: douta=16'hcc89;
15304: douta=16'hcc89;
15305: douta=16'hcc89;
15306: douta=16'hcc69;
15307: douta=16'hcc89;
15308: douta=16'hcc89;
15309: douta=16'hcc69;
15310: douta=16'hcc69;
15311: douta=16'hcc89;
15312: douta=16'hcc89;
15313: douta=16'hb595;
15314: douta=16'hcc49;
15315: douta=16'hcc6a;
15316: douta=16'hcc69;
15317: douta=16'hcc6a;
15318: douta=16'hcc6a;
15319: douta=16'hcc69;
15320: douta=16'hcc69;
15321: douta=16'hcc49;
15322: douta=16'hcc69;
15323: douta=16'hc449;
15324: douta=16'hcc69;
15325: douta=16'hcc49;
15326: douta=16'hc449;
15327: douta=16'hc449;
15328: douta=16'hc469;
15329: douta=16'hc449;
15330: douta=16'hc449;
15331: douta=16'hc449;
15332: douta=16'hc44a;
15333: douta=16'hc429;
15334: douta=16'hbc29;
15335: douta=16'hc429;
15336: douta=16'hc429;
15337: douta=16'hc40a;
15338: douta=16'hbc2a;
15339: douta=16'hbc2a;
15340: douta=16'hbc09;
15341: douta=16'hbc09;
15342: douta=16'hbc09;
15343: douta=16'hbc09;
15344: douta=16'hbbe9;
15345: douta=16'hb3e9;
15346: douta=16'hb3e9;
15347: douta=16'hb3e9;
15348: douta=16'hb3e9;
15349: douta=16'hb3c9;
15350: douta=16'hb3c9;
15351: douta=16'habc9;
15352: douta=16'habc9;
15353: douta=16'habc9;
15354: douta=16'haba9;
15355: douta=16'habc9;
15356: douta=16'haba9;
15357: douta=16'haba9;
15358: douta=16'ha389;
15359: douta=16'ha389;
15360: douta=16'h955a;
15361: douta=16'h2924;
15362: douta=16'h2904;
15363: douta=16'h2904;
15364: douta=16'h2904;
15365: douta=16'h2904;
15366: douta=16'h28e3;
15367: douta=16'h20e3;
15368: douta=16'h20e3;
15369: douta=16'h20a3;
15370: douta=16'h20c2;
15371: douta=16'h28c3;
15372: douta=16'h28e3;
15373: douta=16'h28e3;
15374: douta=16'h3103;
15375: douta=16'h3103;
15376: douta=16'h3923;
15377: douta=16'h3944;
15378: douta=16'h4164;
15379: douta=16'h4985;
15380: douta=16'h10e5;
15381: douta=16'h61e4;
15382: douta=16'h59c4;
15383: douta=16'h6204;
15384: douta=16'h6a44;
15385: douta=16'h7245;
15386: douta=16'h736b;
15387: douta=16'h7203;
15388: douta=16'h7a85;
15389: douta=16'h82c6;
15390: douta=16'h82c6;
15391: douta=16'h82c6;
15392: douta=16'h8ae7;
15393: douta=16'h8ae7;
15394: douta=16'h9307;
15395: douta=16'h9b47;
15396: douta=16'h9b47;
15397: douta=16'ha38b;
15398: douta=16'h9b48;
15399: douta=16'h9b05;
15400: douta=16'habc8;
15401: douta=16'hb3c7;
15402: douta=16'hb3e8;
15403: douta=16'hb3e8;
15404: douta=16'hbc08;
15405: douta=16'hbc28;
15406: douta=16'hbc29;
15407: douta=16'hbc28;
15408: douta=16'hc428;
15409: douta=16'hc449;
15410: douta=16'hc449;
15411: douta=16'hc428;
15412: douta=16'hc448;
15413: douta=16'hc448;
15414: douta=16'hcc69;
15415: douta=16'hcc69;
15416: douta=16'hcc69;
15417: douta=16'hcc69;
15418: douta=16'hcc69;
15419: douta=16'hcc69;
15420: douta=16'hcc69;
15421: douta=16'hcc69;
15422: douta=16'hcc69;
15423: douta=16'hcc89;
15424: douta=16'hcc89;
15425: douta=16'hcc69;
15426: douta=16'hcc69;
15427: douta=16'hcc89;
15428: douta=16'hcc89;
15429: douta=16'hcc89;
15430: douta=16'hcc89;
15431: douta=16'hcc89;
15432: douta=16'hcc69;
15433: douta=16'hcc69;
15434: douta=16'hcc69;
15435: douta=16'hcc69;
15436: douta=16'hcc69;
15437: douta=16'hcc89;
15438: douta=16'hcc89;
15439: douta=16'hc489;
15440: douta=16'hcc89;
15441: douta=16'hb5b5;
15442: douta=16'hcc69;
15443: douta=16'hcc6a;
15444: douta=16'hcc89;
15445: douta=16'hcc69;
15446: douta=16'hcc69;
15447: douta=16'hcc69;
15448: douta=16'hcc69;
15449: douta=16'hcc49;
15450: douta=16'hcc69;
15451: douta=16'hc449;
15452: douta=16'hcc6a;
15453: douta=16'hcc49;
15454: douta=16'hc449;
15455: douta=16'hc44a;
15456: douta=16'hc449;
15457: douta=16'hc449;
15458: douta=16'hc449;
15459: douta=16'hc449;
15460: douta=16'hc429;
15461: douta=16'hc44a;
15462: douta=16'hc429;
15463: douta=16'hc429;
15464: douta=16'hc429;
15465: douta=16'hbc09;
15466: douta=16'hbc09;
15467: douta=16'hbc29;
15468: douta=16'hbc09;
15469: douta=16'hbc09;
15470: douta=16'hbc09;
15471: douta=16'hbc09;
15472: douta=16'hbc09;
15473: douta=16'hb3e9;
15474: douta=16'hbc09;
15475: douta=16'hb3e9;
15476: douta=16'hb3e9;
15477: douta=16'hb3e9;
15478: douta=16'hb3ca;
15479: douta=16'hb3c9;
15480: douta=16'habc9;
15481: douta=16'habc9;
15482: douta=16'habc9;
15483: douta=16'habc9;
15484: douta=16'haba9;
15485: douta=16'ha389;
15486: douta=16'habaa;
15487: douta=16'ha389;
15488: douta=16'h4a8b;
15489: douta=16'h2904;
15490: douta=16'h2904;
15491: douta=16'h2904;
15492: douta=16'h2904;
15493: douta=16'h2904;
15494: douta=16'h2904;
15495: douta=16'h20e3;
15496: douta=16'h20e3;
15497: douta=16'h20c2;
15498: douta=16'h20c3;
15499: douta=16'h28e3;
15500: douta=16'h28e3;
15501: douta=16'h2903;
15502: douta=16'h3103;
15503: douta=16'h3903;
15504: douta=16'h3923;
15505: douta=16'h4144;
15506: douta=16'h4964;
15507: douta=16'h4a28;
15508: douta=16'h1085;
15509: douta=16'h59c4;
15510: douta=16'h59e4;
15511: douta=16'h6204;
15512: douta=16'h6a25;
15513: douta=16'h7245;
15514: douta=16'h9491;
15515: douta=16'h7244;
15516: douta=16'h82a5;
15517: douta=16'h82a6;
15518: douta=16'h82c6;
15519: douta=16'h8ae6;
15520: douta=16'h8ac6;
15521: douta=16'h9307;
15522: douta=16'h9327;
15523: douta=16'h9b47;
15524: douta=16'h9b47;
15525: douta=16'ha368;
15526: douta=16'ha368;
15527: douta=16'ha388;
15528: douta=16'haba8;
15529: douta=16'hb3c8;
15530: douta=16'hb3e8;
15531: douta=16'hb3e8;
15532: douta=16'hbbe8;
15533: douta=16'hbc08;
15534: douta=16'hbc08;
15535: douta=16'hbc28;
15536: douta=16'hc429;
15537: douta=16'hc449;
15538: douta=16'hc449;
15539: douta=16'hc449;
15540: douta=16'hc449;
15541: douta=16'hc468;
15542: douta=16'hcc49;
15543: douta=16'hcc69;
15544: douta=16'hcc69;
15545: douta=16'hcc69;
15546: douta=16'hcc69;
15547: douta=16'hcc69;
15548: douta=16'hcc69;
15549: douta=16'hcc89;
15550: douta=16'hcc69;
15551: douta=16'hcc69;
15552: douta=16'hcc89;
15553: douta=16'hcc89;
15554: douta=16'hcc89;
15555: douta=16'hcc69;
15556: douta=16'hcc69;
15557: douta=16'hcc89;
15558: douta=16'hcc89;
15559: douta=16'hcc69;
15560: douta=16'hcc69;
15561: douta=16'hcc89;
15562: douta=16'hcc69;
15563: douta=16'hcc69;
15564: douta=16'hcc69;
15565: douta=16'hcc69;
15566: douta=16'hcc89;
15567: douta=16'hc489;
15568: douta=16'hcc69;
15569: douta=16'hb5d5;
15570: douta=16'hc448;
15571: douta=16'hcc69;
15572: douta=16'hcc6a;
15573: douta=16'hcc69;
15574: douta=16'hcc8a;
15575: douta=16'hcc69;
15576: douta=16'hcc6a;
15577: douta=16'hcc6a;
15578: douta=16'hcc49;
15579: douta=16'hcc6a;
15580: douta=16'hc449;
15581: douta=16'hc449;
15582: douta=16'hc449;
15583: douta=16'hc449;
15584: douta=16'hc449;
15585: douta=16'hc449;
15586: douta=16'hc44a;
15587: douta=16'hc44a;
15588: douta=16'hc429;
15589: douta=16'hc42a;
15590: douta=16'hc40a;
15591: douta=16'hbc29;
15592: douta=16'hbc09;
15593: douta=16'hbc0a;
15594: douta=16'hbc09;
15595: douta=16'hbc2a;
15596: douta=16'hbc09;
15597: douta=16'hbc09;
15598: douta=16'hbc09;
15599: douta=16'hbc09;
15600: douta=16'hbc09;
15601: douta=16'hbc09;
15602: douta=16'hbbe9;
15603: douta=16'hb3e9;
15604: douta=16'hb3c9;
15605: douta=16'hb3c9;
15606: douta=16'habc9;
15607: douta=16'haba9;
15608: douta=16'hb3ca;
15609: douta=16'habc9;
15610: douta=16'habc9;
15611: douta=16'haba9;
15612: douta=16'haba9;
15613: douta=16'ha389;
15614: douta=16'ha389;
15615: douta=16'ha389;
15616: douta=16'h1881;
15617: douta=16'h2924;
15618: douta=16'h3124;
15619: douta=16'h3124;
15620: douta=16'h2904;
15621: douta=16'h2904;
15622: douta=16'h2103;
15623: douta=16'h2103;
15624: douta=16'h2904;
15625: douta=16'h20c3;
15626: douta=16'h28e3;
15627: douta=16'h28e3;
15628: douta=16'h28e3;
15629: douta=16'h28e3;
15630: douta=16'h3123;
15631: douta=16'h3923;
15632: douta=16'h3943;
15633: douta=16'h4144;
15634: douta=16'h4984;
15635: douta=16'h528b;
15636: douta=16'h18a4;
15637: douta=16'h59e4;
15638: douta=16'h61e4;
15639: douta=16'h6204;
15640: douta=16'h6a25;
15641: douta=16'h7245;
15642: douta=16'hb594;
15643: douta=16'h7a85;
15644: douta=16'h82a5;
15645: douta=16'h82c6;
15646: douta=16'h82c6;
15647: douta=16'h8b07;
15648: douta=16'h8b07;
15649: douta=16'h8b07;
15650: douta=16'h9328;
15651: douta=16'h9b47;
15652: douta=16'h9b68;
15653: douta=16'h9b67;
15654: douta=16'h9b67;
15655: douta=16'ha367;
15656: douta=16'hab87;
15657: douta=16'hb3c8;
15658: douta=16'hb3e8;
15659: douta=16'hb3e8;
15660: douta=16'hbbe8;
15661: douta=16'hbc28;
15662: douta=16'hc429;
15663: douta=16'hc449;
15664: douta=16'hc429;
15665: douta=16'hc429;
15666: douta=16'hc429;
15667: douta=16'hc449;
15668: douta=16'hc449;
15669: douta=16'hcc49;
15670: douta=16'hcc69;
15671: douta=16'hcc49;
15672: douta=16'hcc49;
15673: douta=16'hcc69;
15674: douta=16'hcc69;
15675: douta=16'hcc69;
15676: douta=16'hcc6a;
15677: douta=16'hcc6a;
15678: douta=16'hcc6a;
15679: douta=16'hcc6a;
15680: douta=16'hcc6a;
15681: douta=16'hcc69;
15682: douta=16'hcc69;
15683: douta=16'hcc89;
15684: douta=16'hcc89;
15685: douta=16'hcc69;
15686: douta=16'hcc69;
15687: douta=16'hcc6a;
15688: douta=16'hcc69;
15689: douta=16'hcc69;
15690: douta=16'hcc69;
15691: douta=16'hcc6a;
15692: douta=16'hcc6a;
15693: douta=16'hcc89;
15694: douta=16'hcc69;
15695: douta=16'hcc6a;
15696: douta=16'hcc69;
15697: douta=16'hb5b5;
15698: douta=16'hc468;
15699: douta=16'hcc6a;
15700: douta=16'hcc6a;
15701: douta=16'hcc69;
15702: douta=16'hcc8a;
15703: douta=16'hcc49;
15704: douta=16'hcc6a;
15705: douta=16'hcc6a;
15706: douta=16'hcc69;
15707: douta=16'hc449;
15708: douta=16'hc469;
15709: douta=16'hc449;
15710: douta=16'hc44a;
15711: douta=16'hc449;
15712: douta=16'hc469;
15713: douta=16'hc44a;
15714: douta=16'hc44a;
15715: douta=16'hc429;
15716: douta=16'hc429;
15717: douta=16'hc42a;
15718: douta=16'hbc2a;
15719: douta=16'hbc29;
15720: douta=16'hbc09;
15721: douta=16'hbc29;
15722: douta=16'hbc2a;
15723: douta=16'hbc09;
15724: douta=16'hbc09;
15725: douta=16'hbc09;
15726: douta=16'hbc09;
15727: douta=16'hbbe9;
15728: douta=16'hbbe9;
15729: douta=16'hbbe9;
15730: douta=16'hbbe9;
15731: douta=16'hb3e9;
15732: douta=16'hb3e9;
15733: douta=16'hb3ca;
15734: douta=16'hb3c9;
15735: douta=16'hb3c9;
15736: douta=16'haba9;
15737: douta=16'haba9;
15738: douta=16'haba9;
15739: douta=16'haba9;
15740: douta=16'haba9;
15741: douta=16'ha389;
15742: douta=16'ha389;
15743: douta=16'ha369;
15744: douta=16'h2924;
15745: douta=16'h3125;
15746: douta=16'h3124;
15747: douta=16'h2924;
15748: douta=16'h2904;
15749: douta=16'h2904;
15750: douta=16'h28e3;
15751: douta=16'h2103;
15752: douta=16'h2924;
15753: douta=16'h20e3;
15754: douta=16'h28e3;
15755: douta=16'h2903;
15756: douta=16'h2903;
15757: douta=16'h28e3;
15758: douta=16'h3923;
15759: douta=16'h3923;
15760: douta=16'h3944;
15761: douta=16'h4143;
15762: douta=16'h4984;
15763: douta=16'h4a4a;
15764: douta=16'h3924;
15765: douta=16'h59e4;
15766: douta=16'h6205;
15767: douta=16'h6a25;
15768: douta=16'h6a45;
15769: douta=16'h7224;
15770: douta=16'hb572;
15771: douta=16'h7a85;
15772: douta=16'h82a5;
15773: douta=16'h82c6;
15774: douta=16'h8ac7;
15775: douta=16'h8ae7;
15776: douta=16'h8ae7;
15777: douta=16'h9327;
15778: douta=16'h9328;
15779: douta=16'h9b47;
15780: douta=16'h9b68;
15781: douta=16'h9b68;
15782: douta=16'h9b67;
15783: douta=16'ha387;
15784: douta=16'hab87;
15785: douta=16'hb3c8;
15786: douta=16'hb408;
15787: douta=16'hb408;
15788: douta=16'hbc09;
15789: douta=16'hbc09;
15790: douta=16'hbc09;
15791: douta=16'hbc29;
15792: douta=16'hbc49;
15793: douta=16'hc449;
15794: douta=16'hc449;
15795: douta=16'hc449;
15796: douta=16'hc469;
15797: douta=16'hc469;
15798: douta=16'hc46a;
15799: douta=16'hcc8a;
15800: douta=16'hcc6a;
15801: douta=16'hcc6a;
15802: douta=16'hc469;
15803: douta=16'hcc69;
15804: douta=16'hcc8a;
15805: douta=16'hcc69;
15806: douta=16'hcc6a;
15807: douta=16'hcc6a;
15808: douta=16'hcc8a;
15809: douta=16'hcc69;
15810: douta=16'hcc89;
15811: douta=16'hcc89;
15812: douta=16'hcc69;
15813: douta=16'hcc69;
15814: douta=16'hcc69;
15815: douta=16'hcc69;
15816: douta=16'hcc69;
15817: douta=16'hcc69;
15818: douta=16'hcc69;
15819: douta=16'hcc6a;
15820: douta=16'hcc69;
15821: douta=16'hcc69;
15822: douta=16'hcc6a;
15823: douta=16'hcc6a;
15824: douta=16'hcc6a;
15825: douta=16'hb5d5;
15826: douta=16'hcc49;
15827: douta=16'hcc6a;
15828: douta=16'hcc69;
15829: douta=16'hcc69;
15830: douta=16'hcc6a;
15831: douta=16'hcc69;
15832: douta=16'hcc6a;
15833: douta=16'hc46a;
15834: douta=16'hcc69;
15835: douta=16'hc469;
15836: douta=16'hc449;
15837: douta=16'hc449;
15838: douta=16'hc469;
15839: douta=16'hc469;
15840: douta=16'hc44a;
15841: douta=16'hc44a;
15842: douta=16'hc44a;
15843: douta=16'hc44a;
15844: douta=16'hc44a;
15845: douta=16'hc44a;
15846: douta=16'hc42a;
15847: douta=16'hbc2a;
15848: douta=16'hbc2a;
15849: douta=16'hbc2a;
15850: douta=16'hbc09;
15851: douta=16'hbc0a;
15852: douta=16'hbc09;
15853: douta=16'hbc09;
15854: douta=16'hbc09;
15855: douta=16'hbbe9;
15856: douta=16'hbc09;
15857: douta=16'hbbe9;
15858: douta=16'hb3e9;
15859: douta=16'hb3e9;
15860: douta=16'hb3ca;
15861: douta=16'hb3c9;
15862: douta=16'hb3c9;
15863: douta=16'habc9;
15864: douta=16'haba9;
15865: douta=16'haba9;
15866: douta=16'haba9;
15867: douta=16'haba9;
15868: douta=16'haba9;
15869: douta=16'ha389;
15870: douta=16'ha389;
15871: douta=16'ha389;
15872: douta=16'h2945;
15873: douta=16'h2924;
15874: douta=16'h2924;
15875: douta=16'h2924;
15876: douta=16'h2924;
15877: douta=16'h2924;
15878: douta=16'h2904;
15879: douta=16'h2104;
15880: douta=16'h28e3;
15881: douta=16'h20e3;
15882: douta=16'h28e3;
15883: douta=16'h2903;
15884: douta=16'h2904;
15885: douta=16'h3104;
15886: douta=16'h3123;
15887: douta=16'h3923;
15888: douta=16'h3923;
15889: douta=16'h4123;
15890: douta=16'h4984;
15891: douta=16'h39a8;
15892: douta=16'h51a5;
15893: douta=16'h59e5;
15894: douta=16'h6205;
15895: douta=16'h6a25;
15896: douta=16'h6a45;
15897: douta=16'h7245;
15898: douta=16'h9c2d;
15899: douta=16'h7a85;
15900: douta=16'h82a6;
15901: douta=16'h82c6;
15902: douta=16'h82c6;
15903: douta=16'h8ae7;
15904: douta=16'h8ae6;
15905: douta=16'h8b07;
15906: douta=16'h9328;
15907: douta=16'h9b48;
15908: douta=16'h9b68;
15909: douta=16'h9b68;
15910: douta=16'ha368;
15911: douta=16'ha388;
15912: douta=16'haba8;
15913: douta=16'hb3e8;
15914: douta=16'hb3e9;
15915: douta=16'hbc08;
15916: douta=16'hbc29;
15917: douta=16'hbc29;
15918: douta=16'hbc29;
15919: douta=16'hbc29;
15920: douta=16'hbc29;
15921: douta=16'hc449;
15922: douta=16'hc449;
15923: douta=16'hc449;
15924: douta=16'hc469;
15925: douta=16'hc46a;
15926: douta=16'hc46a;
15927: douta=16'hc469;
15928: douta=16'hcc6a;
15929: douta=16'hc469;
15930: douta=16'hcc6a;
15931: douta=16'hcc6a;
15932: douta=16'hcc6a;
15933: douta=16'hcc8a;
15934: douta=16'hc469;
15935: douta=16'hcc6a;
15936: douta=16'hcc8a;
15937: douta=16'hcc6a;
15938: douta=16'hcc6a;
15939: douta=16'hcc6a;
15940: douta=16'hcc6a;
15941: douta=16'hcc69;
15942: douta=16'hcc69;
15943: douta=16'hcc6a;
15944: douta=16'hcc69;
15945: douta=16'hcc69;
15946: douta=16'hcc8a;
15947: douta=16'hcc6a;
15948: douta=16'hcc6a;
15949: douta=16'hcc69;
15950: douta=16'hc469;
15951: douta=16'hcc8a;
15952: douta=16'hcc69;
15953: douta=16'hbdd5;
15954: douta=16'hc449;
15955: douta=16'hcc6a;
15956: douta=16'hcc6a;
15957: douta=16'hc46a;
15958: douta=16'hcc69;
15959: douta=16'hcc69;
15960: douta=16'hcc69;
15961: douta=16'hcc6a;
15962: douta=16'hc46a;
15963: douta=16'hc469;
15964: douta=16'hc46a;
15965: douta=16'hc44a;
15966: douta=16'hc44a;
15967: douta=16'hc44a;
15968: douta=16'hc44a;
15969: douta=16'hc429;
15970: douta=16'hc429;
15971: douta=16'hc44a;
15972: douta=16'hc44a;
15973: douta=16'hc42a;
15974: douta=16'hbc2a;
15975: douta=16'hbc2a;
15976: douta=16'hbc29;
15977: douta=16'hbc2a;
15978: douta=16'hbc0a;
15979: douta=16'hbc0a;
15980: douta=16'hbc0a;
15981: douta=16'hbc09;
15982: douta=16'hbc09;
15983: douta=16'hbc09;
15984: douta=16'hb3e9;
15985: douta=16'hb3e9;
15986: douta=16'hb3e9;
15987: douta=16'hb3e9;
15988: douta=16'hb3ca;
15989: douta=16'hb3ca;
15990: douta=16'haba9;
15991: douta=16'haba9;
15992: douta=16'haba9;
15993: douta=16'haba9;
15994: douta=16'haba9;
15995: douta=16'hab89;
15996: douta=16'hab89;
15997: douta=16'ha389;
15998: douta=16'hab89;
15999: douta=16'ha389;
16000: douta=16'h3145;
16001: douta=16'h2924;
16002: douta=16'h2904;
16003: douta=16'h2904;
16004: douta=16'h2924;
16005: douta=16'h2904;
16006: douta=16'h2924;
16007: douta=16'h2104;
16008: douta=16'h20c3;
16009: douta=16'h20e3;
16010: douta=16'h28e3;
16011: douta=16'h28e3;
16012: douta=16'h2903;
16013: douta=16'h3103;
16014: douta=16'h3123;
16015: douta=16'h3923;
16016: douta=16'h3923;
16017: douta=16'h4164;
16018: douta=16'h4163;
16019: douta=16'h1906;
16020: douta=16'h59c4;
16021: douta=16'h59e5;
16022: douta=16'h6205;
16023: douta=16'h6a25;
16024: douta=16'h7265;
16025: douta=16'h7ae9;
16026: douta=16'h82e7;
16027: douta=16'h82a6;
16028: douta=16'h82c6;
16029: douta=16'h82c6;
16030: douta=16'h8ac7;
16031: douta=16'h8ae7;
16032: douta=16'h8b07;
16033: douta=16'h8b07;
16034: douta=16'h9328;
16035: douta=16'h9b28;
16036: douta=16'h9b48;
16037: douta=16'ha388;
16038: douta=16'ha368;
16039: douta=16'ha387;
16040: douta=16'haba8;
16041: douta=16'hb3e8;
16042: douta=16'hb409;
16043: douta=16'hb409;
16044: douta=16'hbc2a;
16045: douta=16'hbc2a;
16046: douta=16'hc42a;
16047: douta=16'hbc29;
16048: douta=16'hbc29;
16049: douta=16'hc449;
16050: douta=16'hc449;
16051: douta=16'hc469;
16052: douta=16'hc44a;
16053: douta=16'hc46a;
16054: douta=16'hcc8b;
16055: douta=16'hc46a;
16056: douta=16'hc46a;
16057: douta=16'hc48a;
16058: douta=16'hcc8a;
16059: douta=16'hcc89;
16060: douta=16'hcc6a;
16061: douta=16'hcc6a;
16062: douta=16'hcc6a;
16063: douta=16'hc469;
16064: douta=16'hcc6a;
16065: douta=16'hcc89;
16066: douta=16'hcc8a;
16067: douta=16'hcc6a;
16068: douta=16'hcc6a;
16069: douta=16'hcc6a;
16070: douta=16'hcc69;
16071: douta=16'hcc6a;
16072: douta=16'hcc6a;
16073: douta=16'hcc6a;
16074: douta=16'hcc6a;
16075: douta=16'hcc6a;
16076: douta=16'hcc69;
16077: douta=16'hcc6a;
16078: douta=16'hcc8a;
16079: douta=16'hcc8a;
16080: douta=16'hcc69;
16081: douta=16'hbdd6;
16082: douta=16'hcc49;
16083: douta=16'hcc6a;
16084: douta=16'hc46a;
16085: douta=16'hc46a;
16086: douta=16'hc469;
16087: douta=16'hc449;
16088: douta=16'hc46a;
16089: douta=16'hc44a;
16090: douta=16'hc449;
16091: douta=16'hc469;
16092: douta=16'hc44a;
16093: douta=16'hc44a;
16094: douta=16'hc44a;
16095: douta=16'hc44a;
16096: douta=16'hc44a;
16097: douta=16'hc44a;
16098: douta=16'hc44a;
16099: douta=16'hc44a;
16100: douta=16'hbc2a;
16101: douta=16'hbc2a;
16102: douta=16'hbc2a;
16103: douta=16'hbc2a;
16104: douta=16'hbc29;
16105: douta=16'hbc2a;
16106: douta=16'hbc0a;
16107: douta=16'hbc09;
16108: douta=16'hbc09;
16109: douta=16'hbc09;
16110: douta=16'hbc09;
16111: douta=16'hb3ea;
16112: douta=16'hb3e9;
16113: douta=16'hb3e9;
16114: douta=16'hb3e9;
16115: douta=16'hb3ca;
16116: douta=16'hb3ca;
16117: douta=16'hb3e9;
16118: douta=16'habca;
16119: douta=16'haba9;
16120: douta=16'haba9;
16121: douta=16'haba9;
16122: douta=16'habaa;
16123: douta=16'ha389;
16124: douta=16'hab89;
16125: douta=16'ha369;
16126: douta=16'ha389;
16127: douta=16'ha389;
16128: douta=16'h3145;
16129: douta=16'h2944;
16130: douta=16'h2924;
16131: douta=16'h28e3;
16132: douta=16'h2904;
16133: douta=16'h2904;
16134: douta=16'h2104;
16135: douta=16'h20e4;
16136: douta=16'h20c3;
16137: douta=16'h20e3;
16138: douta=16'h28e3;
16139: douta=16'h2903;
16140: douta=16'h3104;
16141: douta=16'h3124;
16142: douta=16'h3944;
16143: douta=16'h3944;
16144: douta=16'h4164;
16145: douta=16'h4964;
16146: douta=16'h4965;
16147: douta=16'h10a3;
16148: douta=16'h59c4;
16149: douta=16'h59e5;
16150: douta=16'h6205;
16151: douta=16'h6a45;
16152: douta=16'h7266;
16153: douta=16'h7bcf;
16154: douta=16'h7245;
16155: douta=16'h82a6;
16156: douta=16'h82c7;
16157: douta=16'h8ae7;
16158: douta=16'h8ae6;
16159: douta=16'h8b07;
16160: douta=16'h8b07;
16161: douta=16'h9308;
16162: douta=16'h9348;
16163: douta=16'h9b48;
16164: douta=16'h9b69;
16165: douta=16'h9b48;
16166: douta=16'ha388;
16167: douta=16'ha3a8;
16168: douta=16'haba8;
16169: douta=16'hb3e9;
16170: douta=16'hb3e9;
16171: douta=16'hbc09;
16172: douta=16'hbc2a;
16173: douta=16'hbc2a;
16174: douta=16'hbc2a;
16175: douta=16'hbc49;
16176: douta=16'hbc29;
16177: douta=16'hc44a;
16178: douta=16'hc44a;
16179: douta=16'hc44a;
16180: douta=16'hc44a;
16181: douta=16'hc48a;
16182: douta=16'hc46a;
16183: douta=16'hc48a;
16184: douta=16'hc46a;
16185: douta=16'hcc6a;
16186: douta=16'hc48a;
16187: douta=16'hcc8a;
16188: douta=16'hcc6a;
16189: douta=16'hcc6a;
16190: douta=16'hcc6a;
16191: douta=16'hcc8a;
16192: douta=16'hcc6a;
16193: douta=16'hc489;
16194: douta=16'hc469;
16195: douta=16'hcc6a;
16196: douta=16'hcc6a;
16197: douta=16'hcc6a;
16198: douta=16'hcc69;
16199: douta=16'hcc6a;
16200: douta=16'hcc6a;
16201: douta=16'hcc6a;
16202: douta=16'hcc6a;
16203: douta=16'hcc6a;
16204: douta=16'hcc6a;
16205: douta=16'hcc6a;
16206: douta=16'hcc6a;
16207: douta=16'hcc6a;
16208: douta=16'hcc69;
16209: douta=16'hbdf6;
16210: douta=16'hcc69;
16211: douta=16'hcc6a;
16212: douta=16'hcc8a;
16213: douta=16'hc469;
16214: douta=16'hc469;
16215: douta=16'hc469;
16216: douta=16'hc469;
16217: douta=16'hc469;
16218: douta=16'hc469;
16219: douta=16'hc44a;
16220: douta=16'hc44a;
16221: douta=16'hc44a;
16222: douta=16'hc429;
16223: douta=16'hc44a;
16224: douta=16'hc44a;
16225: douta=16'hc44a;
16226: douta=16'hc42a;
16227: douta=16'hc42a;
16228: douta=16'hc42a;
16229: douta=16'hbc2a;
16230: douta=16'hbc2a;
16231: douta=16'hbc2a;
16232: douta=16'hbc0a;
16233: douta=16'hbc09;
16234: douta=16'hbc0a;
16235: douta=16'hbc09;
16236: douta=16'hb3e9;
16237: douta=16'hbc0a;
16238: douta=16'hb40a;
16239: douta=16'hb40a;
16240: douta=16'hb3ea;
16241: douta=16'hb3e9;
16242: douta=16'hb3ca;
16243: douta=16'hb3ca;
16244: douta=16'hb3e9;
16245: douta=16'habc9;
16246: douta=16'habc9;
16247: douta=16'habc9;
16248: douta=16'hb3ca;
16249: douta=16'habaa;
16250: douta=16'habaa;
16251: douta=16'ha389;
16252: douta=16'habaa;
16253: douta=16'ha38a;
16254: douta=16'ha369;
16255: douta=16'ha38a;
16256: douta=16'h2925;
16257: douta=16'h2924;
16258: douta=16'h2924;
16259: douta=16'h2104;
16260: douta=16'h2104;
16261: douta=16'h2104;
16262: douta=16'h2104;
16263: douta=16'h2924;
16264: douta=16'h20e3;
16265: douta=16'h20e3;
16266: douta=16'h28e3;
16267: douta=16'h28e3;
16268: douta=16'h3124;
16269: douta=16'h3124;
16270: douta=16'h3924;
16271: douta=16'h4144;
16272: douta=16'h4164;
16273: douta=16'h4185;
16274: douta=16'h49c6;
16275: douta=16'h1084;
16276: douta=16'h59c5;
16277: douta=16'h59e4;
16278: douta=16'h6205;
16279: douta=16'h6a25;
16280: douta=16'h7266;
16281: douta=16'h94f4;
16282: douta=16'h7a66;
16283: douta=16'h82a7;
16284: douta=16'h82c7;
16285: douta=16'h82c6;
16286: douta=16'h8ae6;
16287: douta=16'h8b07;
16288: douta=16'h9308;
16289: douta=16'h9328;
16290: douta=16'h9348;
16291: douta=16'h9b48;
16292: douta=16'h9b69;
16293: douta=16'h9b48;
16294: douta=16'ha369;
16295: douta=16'ha388;
16296: douta=16'habc8;
16297: douta=16'hb3e9;
16298: douta=16'hb3e9;
16299: douta=16'hb409;
16300: douta=16'hb42a;
16301: douta=16'hbc2a;
16302: douta=16'hbc2a;
16303: douta=16'hbc2a;
16304: douta=16'hbc2a;
16305: douta=16'hc44a;
16306: douta=16'hc44a;
16307: douta=16'hc44a;
16308: douta=16'hc46b;
16309: douta=16'hc46a;
16310: douta=16'hc46a;
16311: douta=16'hc48a;
16312: douta=16'hc46a;
16313: douta=16'hc46a;
16314: douta=16'hc46a;
16315: douta=16'hcc8a;
16316: douta=16'hc48a;
16317: douta=16'hc46a;
16318: douta=16'hc489;
16319: douta=16'hcc6a;
16320: douta=16'hcc6a;
16321: douta=16'hcc6a;
16322: douta=16'hcc6a;
16323: douta=16'hcc6a;
16324: douta=16'hcc6a;
16325: douta=16'hc469;
16326: douta=16'hc469;
16327: douta=16'hcc6a;
16328: douta=16'hcc6a;
16329: douta=16'hc46a;
16330: douta=16'hc46a;
16331: douta=16'hcc6a;
16332: douta=16'hcc6a;
16333: douta=16'hcc6a;
16334: douta=16'hcc6a;
16335: douta=16'hc46a;
16336: douta=16'hcc69;
16337: douta=16'hbe16;
16338: douta=16'hc44a;
16339: douta=16'hc469;
16340: douta=16'hc46a;
16341: douta=16'hc469;
16342: douta=16'hc46a;
16343: douta=16'hc469;
16344: douta=16'hc469;
16345: douta=16'hc46a;
16346: douta=16'hc44a;
16347: douta=16'hc44a;
16348: douta=16'hc44a;
16349: douta=16'hc44a;
16350: douta=16'hc44a;
16351: douta=16'hc44a;
16352: douta=16'hc42a;
16353: douta=16'hc44a;
16354: douta=16'hc44a;
16355: douta=16'hc42a;
16356: douta=16'hbc2a;
16357: douta=16'hbc2a;
16358: douta=16'hbc2a;
16359: douta=16'hbc2a;
16360: douta=16'hbc0a;
16361: douta=16'hbc0a;
16362: douta=16'hbc0a;
16363: douta=16'hbc09;
16364: douta=16'hb40a;
16365: douta=16'hb40a;
16366: douta=16'hb3ea;
16367: douta=16'hb3ea;
16368: douta=16'hb3e9;
16369: douta=16'hb3ea;
16370: douta=16'habc9;
16371: douta=16'habca;
16372: douta=16'hb3ca;
16373: douta=16'habca;
16374: douta=16'habca;
16375: douta=16'haba9;
16376: douta=16'habaa;
16377: douta=16'habaa;
16378: douta=16'habaa;
16379: douta=16'hab89;
16380: douta=16'ha389;
16381: douta=16'ha389;
16382: douta=16'ha369;
16383: douta=16'ha369;

default :douta  =	16'h	0000;
endcase
end


endmodule 
