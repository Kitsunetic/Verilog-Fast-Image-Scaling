module bufferram (
  input [16:0] addra,      
  output reg [15:0] douta 
);

always@(*) begin
  case(addra)
0	:douta	=	16'h	74d9;
1	:douta	=	16'h	5c16;
2	:douta	=	16'h	6cba;
3	:douta	=	16'h	32b0;
4	:douta	=	16'h	4311;
5	:douta	=	16'h	5394;
6	:douta	=	16'h	6436;
7	:douta	=	16'h	6c77;
8	:douta	=	16'h	6c14;
9	:douta	=	16'h	7c98;
10	:douta	=	16'h	7414;
11	:douta	=	16'h	7c76;
12	:douta	=	16'h	6435;
13	:douta	=	16'h	4b32;
14	:douta	=	16'h	31ea;
15	:douta	=	16'h	6c15;
16	:douta	=	16'h	31c8;
17	:douta	=	16'h	10a3;
18	:douta	=	16'h	b536;
19	:douta	=	16'h	a536;
20	:douta	=	16'h	b597;
21	:douta	=	16'h	84d6;
22	:douta	=	16'h	6bd3;
23	:douta	=	16'h	9516;
24	:douta	=	16'h	322d;
25	:douta	=	16'h	63b2;
26	:douta	=	16'h	326f;
27	:douta	=	16'h	9d37;
28	:douta	=	16'h	9d36;
29	:douta	=	16'h	a578;
30	:douta	=	16'h	ce19;
31	:douta	=	16'h	84b6;
32	:douta	=	16'h	8c95;
33	:douta	=	16'h	b5d8;
34	:douta	=	16'h	5bb2;
35	:douta	=	16'h	8494;
36	:douta	=	16'h	94f6;
37	:douta	=	16'h	bdf8;
38	:douta	=	16'h	c659;
39	:douta	=	16'h	d618;
40	:douta	=	16'h	ffbc;
41	:douta	=	16'h	b5d9;
42	:douta	=	16'h	8454;
43	:douta	=	16'h	6b50;
44	:douta	=	16'h	6bd2;
45	:douta	=	16'h	9d15;
46	:douta	=	16'h	5bd4;
47	:douta	=	16'h	94f5;
48	:douta	=	16'h	e6fb;
49	:douta	=	16'h	ce18;
50	:douta	=	16'h	d6da;
51	:douta	=	16'h	5b52;
52	:douta	=	16'h	8cb4;
53	:douta	=	16'h	53d4;
54	:douta	=	16'h	63b2;
55	:douta	=	16'h	ad36;
56	:douta	=	16'h	d678;
57	:douta	=	16'h	de99;
58	:douta	=	16'h	94d6;
59	:douta	=	16'h	f77b;
60	:douta	=	16'h	7c75;
61	:douta	=	16'h	9cd6;
62	:douta	=	16'h	ad97;
63	:douta	=	16'h	3ad1;
64	:douta	=	16'h	7454;
65	:douta	=	16'h	7c54;
66	:douta	=	16'h	ad77;
67	:douta	=	16'h	b5b8;
68	:douta	=	16'h	e6b9;
69	:douta	=	16'h	be18;
70	:douta	=	16'h	94d6;
71	:douta	=	16'h	ad98;
72	:douta	=	16'h	9cd4;
73	:douta	=	16'h	73d3;
74	:douta	=	16'h	5392;
75	:douta	=	16'h	3b11;
76	:douta	=	16'h	b5d8;
77	:douta	=	16'h	b556;
78	:douta	=	16'h	a576;
79	:douta	=	16'h	7415;
80	:douta	=	16'h	b5b8;
81	:douta	=	16'h	adda;
82	:douta	=	16'h	6c58;
83	:douta	=	16'h	d6ba;
84	:douta	=	16'h	2a90;
85	:douta	=	16'h	7455;
86	:douta	=	16'h	8cd3;
87	:douta	=	16'h	7cb6;
88	:douta	=	16'h	d6fa;
89	:douta	=	16'h	be7b;
90	:douta	=	16'h	cebb;
91	:douta	=	16'h	ae1b;
92	:douta	=	16'h	6437;
93	:douta	=	16'h	a599;
94	:douta	=	16'h	4b73;
95	:douta	=	16'h	6435;
96	:douta	=	16'h	7454;
97	:douta	=	16'h	7cd7;
98	:douta	=	16'h	c67a;
99	:douta	=	16'h	a598;
100	:douta	=	16'h	ad98;
101	:douta	=	16'h	a5ba;
102	:douta	=	16'h	5bd5;
103	:douta	=	16'h	94d6;
104	:douta	=	16'h	3b11;
105	:douta	=	16'h	8c95;
106	:douta	=	16'h	b639;
107	:douta	=	16'h	bdd8;
108	:douta	=	16'h	ce9b;
109	:douta	=	16'h	959b;
110	:douta	=	16'h	7c34;
111	:douta	=	16'h	6c76;
112	:douta	=	16'h	6c35;
113	:douta	=	16'h	2ab0;
114	:douta	=	16'h	7474;
115	:douta	=	16'h	9598;
116	:douta	=	16'h	a578;
117	:douta	=	16'h	cedc;
118	:douta	=	16'h	7455;
119	:douta	=	16'h	a536;
120	:douta	=	16'h	add8;
121	:douta	=	16'h	5b0f;
122	:douta	=	16'h	9d15;
123	:douta	=	16'h	21ab;
124	:douta	=	16'h	5b71;
125	:douta	=	16'h	8c93;
126	:douta	=	16'h	2a2c;
127	:douta	=	16'h	7474;
128	:douta	=	16'h	bdd8;
129	:douta	=	16'h	94f6;
130	:douta	=	16'h	f77c;
131	:douta	=	16'h	ce18;
132	:douta	=	16'h	bdd7;
133	:douta	=	16'h	5b50;
134	:douta	=	16'h	6b90;
135	:douta	=	16'h	8c92;
136	:douta	=	16'h	638f;
137	:douta	=	16'h	8432;
138	:douta	=	16'h	e6f9;
139	:douta	=	16'h	8472;
140	:douta	=	16'h	d636;
141	:douta	=	16'h	734f;
142	:douta	=	16'h	9c30;
143	:douta	=	16'h	5b4f;
144	:douta	=	16'h	2169;
145	:douta	=	16'h	29a8;
146	:douta	=	16'h	94d2;
147	:douta	=	16'h	ce99;
148	:douta	=	16'h	6b90;
149	:douta	=	16'h	630d;
150	:douta	=	16'h	d677;
151	:douta	=	16'h	5a6b;
152	:douta	=	16'h	736f;
153	:douta	=	16'h	1107;
154	:douta	=	16'h	08a5;
155	:douta	=	16'h	52ee;
156	:douta	=	16'h	5b4f;
157	:douta	=	16'h	534e;
158	:douta	=	16'h	8c72;
159	:douta	=	16'h	9d14;
160	:douta	=	16'h	a4f2;
161	:douta	=	16'h	b575;
162	:douta	=	16'h	5b0e;
163	:douta	=	16'h	8c10;
164	:douta	=	16'h	8430;
165	:douta	=	16'h	6b6f;
166	:douta	=	16'h	0908;
167	:douta	=	16'h	1149;
168	:douta	=	16'h	6b6f;
169	:douta	=	16'h	b575;
170	:douta	=	16'h	5acc;
171	:douta	=	16'h	e695;
172	:douta	=	16'h	5b30;
173	:douta	=	16'h	b533;
174	:douta	=	16'h	c5d6;
175	:douta	=	16'h	1109;
176	:douta	=	16'h	52ac;
177	:douta	=	16'h	324c;
178	:douta	=	16'h	324c;
179	:douta	=	16'h	326d;
180	:douta	=	16'h	29c9;
181	:douta	=	16'h	8431;
182	:douta	=	16'h	7411;
183	:douta	=	16'h	a4d3;
184	:douta	=	16'h	94b2;
185	:douta	=	16'h	ad34;
186	:douta	=	16'h	94b4;
187	:douta	=	16'h	2966;
188	:douta	=	16'h	10e5;
189	:douta	=	16'h	10c4;
190	:douta	=	16'h	0043;
191	:douta	=	16'h	7bcf;
192	:douta	=	16'h	8452;
193	:douta	=	16'h	a4f3;
194	:douta	=	16'h	5ace;
195	:douta	=	16'h	7c74;
196	:douta	=	16'h	42f0;
197	:douta	=	16'h	636f;
198	:douta	=	16'h	532f;
199	:douta	=	16'h	73f2;
200	:douta	=	16'h	94f5;
201	:douta	=	16'h	63f4;
202	:douta	=	16'h	8453;
203	:douta	=	16'h	7c54;
204	:douta	=	16'h	4b31;
205	:douta	=	16'h	7c55;
206	:douta	=	16'h	3ad0;
207	:douta	=	16'h	5b71;
208	:douta	=	16'h	3ace;
209	:douta	=	16'h	8493;
210	:douta	=	16'h	b5d7;
211	:douta	=	16'h	6bf4;
212	:douta	=	16'h	a515;
213	:douta	=	16'h	5372;
214	:douta	=	16'h	73f4;
215	:douta	=	16'h	19ee;
216	:douta	=	16'h	63f4;
217	:douta	=	16'h	bdd8;
218	:douta	=	16'h	9518;
219	:douta	=	16'h	a599;
220	:douta	=	16'h	74b8;
221	:douta	=	16'h	7c96;
222	:douta	=	16'h	a558;
223	:douta	=	16'h	4373;
224	:douta	=	16'h	5bd4;
225	:douta	=	16'h	2a90;
226	:douta	=	16'h	4b11;
227	:douta	=	16'h	5371;
228	:douta	=	16'h	84d5;
229	:douta	=	16'h	c67a;
230	:douta	=	16'h	6c99;
231	:douta	=	16'h	7cb8;
232	:douta	=	16'h	7d19;
233	:douta	=	16'h	3b12;
234	:douta	=	16'h	2a6f;
235	:douta	=	16'h	5352;
236	:douta	=	16'h	5b92;
237	:douta	=	16'h	7cb7;
238	:douta	=	16'h	a5bb;
239	:douta	=	16'h	74d9;
240	:douta	=	16'h	118a;
241	:douta	=	16'h	3ab0;
242	:douta	=	16'h	19ed;
243	:douta	=	16'h	6c55;
244	:douta	=	16'h	7476;
245	:douta	=	16'h	9d9b;
246	:douta	=	16'h	8d7c;
247	:douta	=	16'h	7cd9;
248	:douta	=	16'h	2b35;
249	:douta	=	16'h	2ab2;
250	:douta	=	16'h	4b53;
251	:douta	=	16'h	6c57;
252	:douta	=	16'h	8519;
253	:douta	=	16'h	7cf9;
254	:douta	=	16'h	3b54;
255	:douta	=	16'h	5c37;
256	:douta	=	16'h	3ad2;
257	:douta	=	16'h	328f;
258	:douta	=	16'h	2a4f;
259	:douta	=	16'h	5373;
260	:douta	=	16'h	7497;
261	:douta	=	16'h	5bb4;
262	:douta	=	16'h	7498;
263	:douta	=	16'h	53f6;
264	:douta	=	16'h	42f1;
265	:douta	=	16'h	4af0;
266	:douta	=	16'h	5b72;
267	:douta	=	16'h	8cd7;
268	:douta	=	16'h	84b6;
269	:douta	=	16'h	9d79;
270	:douta	=	16'h	ad78;
271	:douta	=	16'h	8d18;
272	:douta	=	16'h	528d;
273	:douta	=	16'h	2127;
274	:douta	=	16'h	6392;
275	:douta	=	16'h	8494;
276	:douta	=	16'h	8c94;
277	:douta	=	16'h	adb8;
278	:douta	=	16'h	8495;
279	:douta	=	16'h	ded9;
280	:douta	=	16'h	ce39;
281	:douta	=	16'h	deba;
282	:douta	=	16'h	adb9;
283	:douta	=	16'h	a537;
284	:douta	=	16'h	8c96;
285	:douta	=	16'h	5b52;
286	:douta	=	16'h	6bf2;
287	:douta	=	16'h	8cb6;
288	:douta	=	16'h	a577;
289	:douta	=	16'h	deba;
290	:douta	=	16'h	d65a;
291	:douta	=	16'h	d6ba;
292	:douta	=	16'h	9d17;
293	:douta	=	16'h	a557;
294	:douta	=	16'h	9599;
295	:douta	=	16'h	3a4c;
296	:douta	=	16'h	a4d3;
297	:douta	=	16'h	7bf3;
298	:douta	=	16'h	d679;
299	:douta	=	16'h	e6da;
300	:douta	=	16'h	ce7a;
301	:douta	=	16'h	e6da;
302	:douta	=	16'h	7cb7;
303	:douta	=	16'h	8434;
304	:douta	=	16'h	c67a;
305	:douta	=	16'h	7c95;
306	:douta	=	16'h	84b5;
307	:douta	=	16'h	a536;
308	:douta	=	16'h	f73c;
309	:douta	=	16'h	b5f9;
310	:douta	=	16'h	be5a;
311	:douta	=	16'h	7436;
312	:douta	=	16'h	8c73;
313	:douta	=	16'h	b597;
314	:douta	=	16'h	226e;
315	:douta	=	16'h	bdf8;
316	:douta	=	16'h	a556;
317	:douta	=	16'h	e6da;
318	:douta	=	16'h	ef3b;
319	:douta	=	16'h	c5f8;
320	:douta	=	16'h	7455;
321	:douta	=	16'h	63b4;
322	:douta	=	16'h	d69a;
323	:douta	=	16'h	9559;
324	:douta	=	16'h	42cf;
325	:douta	=	16'h	9535;
326	:douta	=	16'h	7c54;
327	:douta	=	16'h	ad75;
328	:douta	=	16'h	c658;
329	:douta	=	16'h	e6ba;
330	:douta	=	16'h	adda;
331	:douta	=	16'h	8c97;
332	:douta	=	16'h	add8;
333	:douta	=	16'h	53b3;
334	:douta	=	16'h	bdb6;
335	:douta	=	16'h	6c15;
336	:douta	=	16'h	63f3;
337	:douta	=	16'h	6bf2;
338	:douta	=	16'h	7c96;
339	:douta	=	16'h	84b5;
340	:douta	=	16'h	bdf8;
341	:douta	=	16'h	d67a;
342	:douta	=	16'h	9dd9;
343	:douta	=	16'h	5373;
344	:douta	=	16'h	9558;
345	:douta	=	16'h	3b12;
346	:douta	=	16'h	be1a;
347	:douta	=	16'h	6c55;
348	:douta	=	16'h	7cb6;
349	:douta	=	16'h	be7b;
350	:douta	=	16'h	84f8;
351	:douta	=	16'h	d69b;
352	:douta	=	16'h	95db;
353	:douta	=	16'h	4b52;
354	:douta	=	16'h	3ab0;
355	:douta	=	16'h	19ee;
356	:douta	=	16'h	74d7;
357	:douta	=	16'h	74b8;
358	:douta	=	16'h	7415;
359	:douta	=	16'h	a5ba;
360	:douta	=	16'h	8cf9;
361	:douta	=	16'h	ceba;
362	:douta	=	16'h	42d0;
363	:douta	=	16'h	ad98;
364	:douta	=	16'h	9d98;
365	:douta	=	16'h	9558;
366	:douta	=	16'h	8cf6;
367	:douta	=	16'h	7c55;
368	:douta	=	16'h	c619;
369	:douta	=	16'h	7c98;
370	:douta	=	16'h	8cb7;
371	:douta	=	16'h	b67c;
372	:douta	=	16'h	7c55;
373	:douta	=	16'h	4b53;
374	:douta	=	16'h	4b0f;
375	:douta	=	16'h	7c12;
376	:douta	=	16'h	6412;
377	:douta	=	16'h	94d4;
378	:douta	=	16'h	7c75;
379	:douta	=	16'h	9d16;
380	:douta	=	16'h	a576;
381	:douta	=	16'h	d6bb;
382	:douta	=	16'h	a558;
383	:douta	=	16'h	8cd6;
384	:douta	=	16'h	4b10;
385	:douta	=	16'h	7454;
386	:douta	=	16'h	6bf3;
387	:douta	=	16'h	8c93;
388	:douta	=	16'h	8493;
389	:douta	=	16'h	a514;
390	:douta	=	16'h	8c12;
391	:douta	=	16'h	ce16;
392	:douta	=	16'h	4a6b;
393	:douta	=	16'h	bd96;
394	:douta	=	16'h	426d;
395	:douta	=	16'h	524a;
396	:douta	=	16'h	3a4b;
397	:douta	=	16'h	9d13;
398	:douta	=	16'h	d6d9;
399	:douta	=	16'h	8c72;
400	:douta	=	16'h	6b70;
401	:douta	=	16'h	8473;
402	:douta	=	16'h	530f;
403	:douta	=	16'h	1989;
404	:douta	=	16'h	634e;
405	:douta	=	16'h	8430;
406	:douta	=	16'h	9c91;
407	:douta	=	16'h	ce56;
408	:douta	=	16'h	b573;
409	:douta	=	16'h	83cf;
410	:douta	=	16'h	bd33;
411	:douta	=	16'h	52ac;
412	:douta	=	16'h	83f1;
413	:douta	=	16'h	6bd1;
414	:douta	=	16'h	31c9;
415	:douta	=	16'h	52ed;
416	:douta	=	16'h	2167;
417	:douta	=	16'h	322a;
418	:douta	=	16'h	6b6f;
419	:douta	=	16'h	ef3a;
420	:douta	=	16'h	d657;
421	:douta	=	16'h	a4d4;
422	:douta	=	16'h	63b1;
423	:douta	=	16'h	5b2f;
424	:douta	=	16'h	31e9;
425	:douta	=	16'h	3a0a;
426	:douta	=	16'h	7bf0;
427	:douta	=	16'h	6b8f;
428	:douta	=	16'h	424b;
429	:douta	=	16'h	8c92;
430	:douta	=	16'h	ad75;
431	:douta	=	16'h	9c92;
432	:douta	=	16'h	ff38;
433	:douta	=	16'h	4b0f;
434	:douta	=	16'h	d659;
435	:douta	=	16'h	5371;
436	:douta	=	16'h	9d16;
437	:douta	=	16'h	4aef;
438	:douta	=	16'h	29ea;
439	:douta	=	16'h	4aae;
440	:douta	=	16'h	4acd;
441	:douta	=	16'h	d677;
442	:douta	=	16'h	bdb6;
443	:douta	=	16'h	2145;
444	:douta	=	16'h	18e5;
445	:douta	=	16'h	10e5;
446	:douta	=	16'h	1905;
447	:douta	=	16'h	320b;
448	:douta	=	16'h	73b0;
449	:douta	=	16'h	00a6;
450	:douta	=	16'h	638e;
451	:douta	=	16'h	6370;
452	:douta	=	16'h	b555;
453	:douta	=	16'h	738f;
454	:douta	=	16'h	5b30;
455	:douta	=	16'h	5b31;
456	:douta	=	16'h	52cc;
457	:douta	=	16'h	94d4;
458	:douta	=	16'h	3a6b;
459	:douta	=	16'h	73f2;
460	:douta	=	16'h	adb6;
461	:douta	=	16'h	63f3;
462	:douta	=	16'h	428f;
463	:douta	=	16'h	ad57;
464	:douta	=	16'h	5bf5;
465	:douta	=	16'h	5393;
466	:douta	=	16'h	7c73;
467	:douta	=	16'h	6bd1;
468	:douta	=	16'h	4331;
469	:douta	=	16'h	ce79;
470	:douta	=	16'h	a577;
471	:douta	=	16'h	7455;
472	:douta	=	16'h	6b91;
473	:douta	=	16'h	6415;
474	:douta	=	16'h	5bd4;
475	:douta	=	16'h	3af0;
476	:douta	=	16'h	7456;
477	:douta	=	16'h	2a6f;
478	:douta	=	16'h	84b6;
479	:douta	=	16'h	ad98;
480	:douta	=	16'h	7477;
481	:douta	=	16'h	8cb5;
482	:douta	=	16'h	8518;
483	:douta	=	16'h	220e;
484	:douta	=	16'h	4b53;
485	:douta	=	16'h	32b0;
486	:douta	=	16'h	198a;
487	:douta	=	16'h	5393;
488	:douta	=	16'h	a578;
489	:douta	=	16'h	7476;
490	:douta	=	16'h	7c76;
491	:douta	=	16'h	6436;
492	:douta	=	16'h	3334;
493	:douta	=	16'h	3b12;
494	:douta	=	16'h	19ee;
495	:douta	=	16'h	3b12;
496	:douta	=	16'h	a5bb;
497	:douta	=	16'h	84b8;
498	:douta	=	16'h	8d7c;
499	:douta	=	16'h	326f;
500	:douta	=	16'h	5331;
501	:douta	=	16'h	5416;
502	:douta	=	16'h	53d5;
503	:douta	=	16'h	6478;
504	:douta	=	16'h	4bf6;
505	:douta	=	16'h	6435;
506	:douta	=	16'h	74d9;
507	:douta	=	16'h	4395;
508	:douta	=	16'h	116d;
509	:douta	=	16'h	32d1;
510	:douta	=	16'h	3b12;
511	:douta	=	16'h	6c77;
512	:douta	=	16'h	5c57;
513	:douta	=	16'h	2a4e;
514	:douta	=	16'h	4b52;
515	:douta	=	16'h	3b11;
516	:douta	=	16'h	4b31;
517	:douta	=	16'h	5b93;
518	:douta	=	16'h	8519;
519	:douta	=	16'h	74b8;
520	:douta	=	16'h	6c35;
521	:douta	=	16'h	5372;
522	:douta	=	16'h	5351;
523	:douta	=	16'h	63b3;
524	:douta	=	16'h	63d4;
525	:douta	=	16'h	6bf3;
526	:douta	=	16'h	c61a;
527	:douta	=	16'h	9537;
528	:douta	=	16'h	b5f9;
529	:douta	=	16'h	9d59;
530	:douta	=	16'h	73f3;
531	:douta	=	16'h	6c13;
532	:douta	=	16'h	52f0;
533	:douta	=	16'h	adb8;
534	:douta	=	16'h	9517;
535	:douta	=	16'h	8495;
536	:douta	=	16'h	ce39;
537	:douta	=	16'h	ce79;
538	:douta	=	16'h	9d37;
539	:douta	=	16'h	d6ba;
540	:douta	=	16'h	de99;
541	:douta	=	16'h	8cd7;
542	:douta	=	16'h	ad57;
543	:douta	=	16'h	3312;
544	:douta	=	16'h	7414;
545	:douta	=	16'h	8494;
546	:douta	=	16'h	adb8;
547	:douta	=	16'h	bdf7;
548	:douta	=	16'h	d679;
549	:douta	=	16'h	dedb;
550	:douta	=	16'h	9d99;
551	:douta	=	16'h	8c53;
552	:douta	=	16'h	cdf8;
553	:douta	=	16'h	7c55;
554	:douta	=	16'h	c618;
555	:douta	=	16'h	8c52;
556	:douta	=	16'h	bdf7;
557	:douta	=	16'h	d638;
558	:douta	=	16'h	ce59;
559	:douta	=	16'h	b5b8;
560	:douta	=	16'h	d6bb;
561	:douta	=	16'h	7c34;
562	:douta	=	16'h	7434;
563	:douta	=	16'h	3a6f;
564	:douta	=	16'h	8c94;
565	:douta	=	16'h	ad97;
566	:douta	=	16'h	c619;
567	:douta	=	16'h	c5f8;
568	:douta	=	16'h	c5f8;
569	:douta	=	16'h	de99;
570	:douta	=	16'h	326f;
571	:douta	=	16'h	6c54;
572	:douta	=	16'h	5b91;
573	:douta	=	16'h	adb7;
574	:douta	=	16'h	b5d8;
575	:douta	=	16'h	e719;
576	:douta	=	16'h	9d37;
577	:douta	=	16'h	a516;
578	:douta	=	16'h	ef3b;
579	:douta	=	16'h	ce7b;
580	:douta	=	16'h	bd97;
581	:douta	=	16'h	5393;
582	:douta	=	16'h	3ab0;
583	:douta	=	16'h	94d4;
584	:douta	=	16'h	84b5;
585	:douta	=	16'h	a555;
586	:douta	=	16'h	9d35;
587	:douta	=	16'h	a517;
588	:douta	=	16'h	defb;
589	:douta	=	16'h	9d36;
590	:douta	=	16'h	d679;
591	:douta	=	16'h	8475;
592	:douta	=	16'h	7455;
593	:douta	=	16'h	b5d8;
594	:douta	=	16'h	74d8;
595	:douta	=	16'h	8cb6;
596	:douta	=	16'h	9516;
597	:douta	=	16'h	ef3c;
598	:douta	=	16'h	9d99;
599	:douta	=	16'h	a516;
600	:douta	=	16'h	c6bd;
601	:douta	=	16'h	6c56;
602	:douta	=	16'h	c618;
603	:douta	=	16'h	4b52;
604	:douta	=	16'h	3a90;
605	:douta	=	16'h	6414;
606	:douta	=	16'h	7434;
607	:douta	=	16'h	be39;
608	:douta	=	16'h	ae1b;
609	:douta	=	16'h	9559;
610	:douta	=	16'h	9559;
611	:douta	=	16'h	5bb5;
612	:douta	=	16'h	63b4;
613	:douta	=	16'h	4332;
614	:douta	=	16'h	2a4e;
615	:douta	=	16'h	5bd3;
616	:douta	=	16'h	9558;
617	:douta	=	16'h	b619;
618	:douta	=	16'h	ad57;
619	:douta	=	16'h	eefa;
620	:douta	=	16'h	6cb8;
621	:douta	=	16'h	6415;
622	:douta	=	16'h	7435;
623	:douta	=	16'h	8cf7;
624	:douta	=	16'h	9579;
625	:douta	=	16'h	7476;
626	:douta	=	16'h	b619;
627	:douta	=	16'h	adda;
628	:douta	=	16'h	c69b;
629	:douta	=	16'h	7497;
630	:douta	=	16'h	6351;
631	:douta	=	16'h	d67a;
632	:douta	=	16'h	4b32;
633	:douta	=	16'h	2a2c;
634	:douta	=	16'h	326d;
635	:douta	=	16'h	84d4;
636	:douta	=	16'h	7412;
637	:douta	=	16'h	8d57;
638	:douta	=	16'h	ceba;
639	:douta	=	16'h	a577;
640	:douta	=	16'h	63d2;
641	:douta	=	16'h	8c74;
642	:douta	=	16'h	6392;
643	:douta	=	16'h	4a8c;
644	:douta	=	16'h	1948;
645	:douta	=	16'h	b575;
646	:douta	=	16'h	a535;
647	:douta	=	16'h	ce78;
648	:douta	=	16'h	a492;
649	:douta	=	16'h	ce16;
650	:douta	=	16'h	7390;
651	:douta	=	16'h	a491;
652	:douta	=	16'h	320a;
653	:douta	=	16'h	2188;
654	:douta	=	16'h	7411;
655	:douta	=	16'h	b595;
656	:douta	=	16'h	c5f7;
657	:douta	=	16'h	9493;
658	:douta	=	16'h	94d4;
659	:douta	=	16'h	42ef;
660	:douta	=	16'h	4a2a;
661	:douta	=	16'h	6b2d;
662	:douta	=	16'h	322a;
663	:douta	=	16'h	5b2c;
664	:douta	=	16'h	632d;
665	:douta	=	16'h	9cd2;
666	:douta	=	16'h	deb7;
667	:douta	=	16'h	9c91;
668	:douta	=	16'h	ce17;
669	:douta	=	16'h	7412;
670	:douta	=	16'h	83af;
671	:douta	=	16'h	94b4;
672	:douta	=	16'h	4a4a;
673	:douta	=	16'h	1927;
674	:douta	=	16'h	3a4b;
675	:douta	=	16'h	9d53;
676	:douta	=	16'h	9d34;
677	:douta	=	16'h	b596;
678	:douta	=	16'h	9d14;
679	:douta	=	16'h	8432;
680	:douta	=	16'h	8c51;
681	:douta	=	16'h	73b0;
682	:douta	=	16'h	634f;
683	:douta	=	16'h	8411;
684	:douta	=	16'h	7bf0;
685	:douta	=	16'h	3a4c;
686	:douta	=	16'h	322b;
687	:douta	=	16'h	636f;
688	:douta	=	16'h	ce57;
689	:douta	=	16'h	7bf1;
690	:douta	=	16'h	ce57;
691	:douta	=	16'h	4aaf;
692	:douta	=	16'h	bdb5;
693	:douta	=	16'h	6b72;
694	:douta	=	16'h	08e8;
695	:douta	=	16'h	42ad;
696	:douta	=	16'h	322c;
697	:douta	=	16'h	4b0c;
698	:douta	=	16'h	63b0;
699	:douta	=	16'h	3187;
700	:douta	=	16'h	10c5;
701	:douta	=	16'h	10c4;
702	:douta	=	16'h	18e6;
703	:douta	=	16'h	4aef;
704	:douta	=	16'h	94d3;
705	:douta	=	16'h	31eb;
706	:douta	=	16'h	21a9;
707	:douta	=	16'h	1968;
708	:douta	=	16'h	5b6e;
709	:douta	=	16'h	ad55;
710	:douta	=	16'h	8433;
711	:douta	=	16'h	7c13;
712	:douta	=	16'h	42af;
713	:douta	=	16'h	21aa;
714	:douta	=	16'h	29eb;
715	:douta	=	16'h	530f;
716	:douta	=	16'h	7433;
717	:douta	=	16'h	4ace;
718	:douta	=	16'h	b534;
719	:douta	=	16'h	c617;
720	:douta	=	16'h	6c15;
721	:douta	=	16'h	63f4;
722	:douta	=	16'h	3aae;
723	:douta	=	16'h	7412;
724	:douta	=	16'h	2ad1;
725	:douta	=	16'h	4311;
726	:douta	=	16'h	7454;
727	:douta	=	16'h	9516;
728	:douta	=	16'h	de9a;
729	:douta	=	16'h	7c56;
730	:douta	=	16'h	7477;
731	:douta	=	16'h	4333;
732	:douta	=	16'h	4331;
733	:douta	=	16'h	328f;
734	:douta	=	16'h	4b53;
735	:douta	=	16'h	84d5;
736	:douta	=	16'h	6c55;
737	:douta	=	16'h	f71b;
738	:douta	=	16'h	a5db;
739	:douta	=	16'h	6b71;
740	:douta	=	16'h	6436;
741	:douta	=	16'h	6c77;
742	:douta	=	16'h	5330;
743	:douta	=	16'h	6416;
744	:douta	=	16'h	3b52;
745	:douta	=	16'h	3ad1;
746	:douta	=	16'h	9517;
747	:douta	=	16'h	6c36;
748	:douta	=	16'h	4b53;
749	:douta	=	16'h	9559;
750	:douta	=	16'h	2a4f;
751	:douta	=	16'h	19cc;
752	:douta	=	16'h	4311;
753	:douta	=	16'h	a537;
754	:douta	=	16'h	5c57;
755	:douta	=	16'h	7c35;
756	:douta	=	16'h	84f8;
757	:douta	=	16'h	3b76;
758	:douta	=	16'h	3b54;
759	:douta	=	16'h	6499;
760	:douta	=	16'h	2270;
761	:douta	=	16'h	6415;
762	:douta	=	16'h	7cd9;
763	:douta	=	16'h	84f9;
764	:douta	=	16'h	4b75;
765	:douta	=	16'h	32f2;
766	:douta	=	16'h	1a2f;
767	:douta	=	16'h	5c15;
768	:douta	=	16'h	6c97;
769	:douta	=	16'h	2a8f;
770	:douta	=	16'h	53b4;
771	:douta	=	16'h	6457;
772	:douta	=	16'h	4b32;
773	:douta	=	16'h	4b73;
774	:douta	=	16'h	53b4;
775	:douta	=	16'h	53f5;
776	:douta	=	16'h	5352;
777	:douta	=	16'h	7c55;
778	:douta	=	16'h	7c75;
779	:douta	=	16'h	9517;
780	:douta	=	16'h	8497;
781	:douta	=	16'h	8cb5;
782	:douta	=	16'h	4333;
783	:douta	=	16'h	5311;
784	:douta	=	16'h	5b51;
785	:douta	=	16'h	5351;
786	:douta	=	16'h	9cd5;
787	:douta	=	16'h	ad98;
788	:douta	=	16'h	de99;
789	:douta	=	16'h	9d78;
790	:douta	=	16'h	add9;
791	:douta	=	16'h	8455;
792	:douta	=	16'h	6bd2;
793	:douta	=	16'h	ad78;
794	:douta	=	16'h	63b4;
795	:douta	=	16'h	8c95;
796	:douta	=	16'h	7454;
797	:douta	=	16'h	9cd6;
798	:douta	=	16'h	bdf7;
799	:douta	=	16'h	84d7;
800	:douta	=	16'h	a578;
801	:douta	=	16'h	e6da;
802	:douta	=	16'h	ad37;
803	:douta	=	16'h	bdd8;
804	:douta	=	16'h	5bb4;
805	:douta	=	16'h	8c94;
806	:douta	=	16'h	ce7a;
807	:douta	=	16'h	a598;
808	:douta	=	16'h	e71a;
809	:douta	=	16'h	b597;
810	:douta	=	16'h	d69a;
811	:douta	=	16'h	bdb6;
812	:douta	=	16'h	ce38;
813	:douta	=	16'h	ad76;
814	:douta	=	16'h	63d3;
815	:douta	=	16'h	73f2;
816	:douta	=	16'h	c638;
817	:douta	=	16'h	ce58;
818	:douta	=	16'h	cebb;
819	:douta	=	16'h	73b2;
820	:douta	=	16'h	f75b;
821	:douta	=	16'h	7c76;
822	:douta	=	16'h	9d77;
823	:douta	=	16'h	4333;
824	:douta	=	16'h	b596;
825	:douta	=	16'h	d678;
826	:douta	=	16'h	ad36;
827	:douta	=	16'h	be7a;
828	:douta	=	16'h	9516;
829	:douta	=	16'h	c5d7;
830	:douta	=	16'h	c699;
831	:douta	=	16'h	9d36;
832	:douta	=	16'h	3b11;
833	:douta	=	16'h	5331;
834	:douta	=	16'h	8412;
835	:douta	=	16'h	d658;
836	:douta	=	16'h	ef3a;
837	:douta	=	16'h	9d37;
838	:douta	=	16'h	b5b6;
839	:douta	=	16'h	d6b9;
840	:douta	=	16'h	9d78;
841	:douta	=	16'h	ce5a;
842	:douta	=	16'h	7496;
843	:douta	=	16'h	3b11;
844	:douta	=	16'h	6371;
845	:douta	=	16'h	8cd5;
846	:douta	=	16'h	84b6;
847	:douta	=	16'h	c5f8;
848	:douta	=	16'h	defb;
849	:douta	=	16'h	f79c;
850	:douta	=	16'h	be19;
851	:douta	=	16'h	c67a;
852	:douta	=	16'h	7435;
853	:douta	=	16'h	7c33;
854	:douta	=	16'h	84d5;
855	:douta	=	16'h	2af0;
856	:douta	=	16'h	4332;
857	:douta	=	16'h	9d36;
858	:douta	=	16'h	deba;
859	:douta	=	16'h	9d58;
860	:douta	=	16'h	d679;
861	:douta	=	16'h	7476;
862	:douta	=	16'h	8496;
863	:douta	=	16'h	8c95;
864	:douta	=	16'h	2250;
865	:douta	=	16'h	42d0;
866	:douta	=	16'h	4332;
867	:douta	=	16'h	84d6;
868	:douta	=	16'h	e75d;
869	:douta	=	16'h	7d3a;
870	:douta	=	16'h	7c77;
871	:douta	=	16'h	8538;
872	:douta	=	16'h	5bd5;
873	:douta	=	16'h	5bf4;
874	:douta	=	16'h	9d58;
875	:douta	=	16'h	9599;
876	:douta	=	16'h	7c96;
877	:douta	=	16'h	a5b9;
878	:douta	=	16'h	c69b;
879	:douta	=	16'h	be39;
880	:douta	=	16'h	9dba;
881	:douta	=	16'h	9cd7;
882	:douta	=	16'h	d69b;
883	:douta	=	16'h	3b32;
884	:douta	=	16'h	63d3;
885	:douta	=	16'h	6bd3;
886	:douta	=	16'h	ad55;
887	:douta	=	16'h	ce59;
888	:douta	=	16'h	9cb6;
889	:douta	=	16'h	ad97;
890	:douta	=	16'h	6c13;
891	:douta	=	16'h	a536;
892	:douta	=	16'h	ce59;
893	:douta	=	16'h	5bb3;
894	:douta	=	16'h	19cd;
895	:douta	=	16'h	21cd;
896	:douta	=	16'h	adb8;
897	:douta	=	16'h	be59;
898	:douta	=	16'h	8433;
899	:douta	=	16'h	ad55;
900	:douta	=	16'h	7c32;
901	:douta	=	16'h	5b0e;
902	:douta	=	16'h	8c52;
903	:douta	=	16'h	2188;
904	:douta	=	16'h	530f;
905	:douta	=	16'h	73f1;
906	:douta	=	16'h	ad54;
907	:douta	=	16'h	a555;
908	:douta	=	16'h	7c51;
909	:douta	=	16'h	d5f6;
910	:douta	=	16'h	9514;
911	:douta	=	16'h	5aee;
912	:douta	=	16'h	5b0f;
913	:douta	=	16'h	6b2e;
914	:douta	=	16'h	8493;
915	:douta	=	16'h	9cd3;
916	:douta	=	16'h	a4b2;
917	:douta	=	16'h	eed8;
918	:douta	=	16'h	52ac;
919	:douta	=	16'h	8c51;
920	:douta	=	16'h	4a8c;
921	:douta	=	16'h	2967;
922	:douta	=	16'h	424c;
923	:douta	=	16'h	634e;
924	:douta	=	16'h	3a6b;
925	:douta	=	16'h	4aad;
926	:douta	=	16'h	eef9;
927	:douta	=	16'h	bdb5;
928	:douta	=	16'h	d657;
929	:douta	=	16'h	630d;
930	:douta	=	16'h	41c9;
931	:douta	=	16'h	8c71;
932	:douta	=	16'h	5b2f;
933	:douta	=	16'h	21a9;
934	:douta	=	16'h	7c12;
935	:douta	=	16'h	636f;
936	:douta	=	16'h	9cd3;
937	:douta	=	16'h	b554;
938	:douta	=	16'h	8431;
939	:douta	=	16'h	73d0;
940	:douta	=	16'h	c5d6;
941	:douta	=	16'h	42f0;
942	:douta	=	16'h	6b4f;
943	:douta	=	16'h	6391;
944	:douta	=	16'h	2a2d;
945	:douta	=	16'h	3a6c;
946	:douta	=	16'h	21c9;
947	:douta	=	16'h	2989;
948	:douta	=	16'h	d657;
949	:douta	=	16'h	8c72;
950	:douta	=	16'h	cdd4;
951	:douta	=	16'h	9cf3;
952	:douta	=	16'h	bdb5;
953	:douta	=	16'h	2a4e;
954	:douta	=	16'h	5b0d;
955	:douta	=	16'h	2105;
956	:douta	=	16'h	10c4;
957	:douta	=	16'h	10c4;
958	:douta	=	16'h	10e5;
959	:douta	=	16'h	3a4c;
960	:douta	=	16'h	5b4f;
961	:douta	=	16'h	b594;
962	:douta	=	16'h	94b3;
963	:douta	=	16'h	52ce;
964	:douta	=	16'h	73b0;
965	:douta	=	16'h	6371;
966	:douta	=	16'h	4ace;
967	:douta	=	16'h	7bf1;
968	:douta	=	16'h	6bb1;
969	:douta	=	16'h	94b3;
970	:douta	=	16'h	9cb3;
971	:douta	=	16'h	9d37;
972	:douta	=	16'h	63d3;
973	:douta	=	16'h	530f;
974	:douta	=	16'h	5bd3;
975	:douta	=	16'h	2a2d;
976	:douta	=	16'h	6bd2;
977	:douta	=	16'h	7c32;
978	:douta	=	16'h	9c94;
979	:douta	=	16'h	bdb7;
980	:douta	=	16'h	7434;
981	:douta	=	16'h	6c56;
982	:douta	=	16'h	328f;
983	:douta	=	16'h	4b31;
984	:douta	=	16'h	3ad0;
985	:douta	=	16'h	9538;
986	:douta	=	16'h	8cf8;
987	:douta	=	16'h	6c34;
988	:douta	=	16'h	ce5a;
989	:douta	=	16'h	8cf9;
990	:douta	=	16'h	6436;
991	:douta	=	16'h	19ee;
992	:douta	=	16'h	3aaf;
993	:douta	=	16'h	2a90;
994	:douta	=	16'h	11ac;
995	:douta	=	16'h	4b31;
996	:douta	=	16'h	5bf5;
997	:douta	=	16'h	8d17;
998	:douta	=	16'h	8d19;
999	:douta	=	16'h	8d18;
1000	:douta	=	16'h	6457;
1001	:douta	=	16'h	7c76;
1002	:douta	=	16'h	9559;
1003	:douta	=	16'h	21ce;
1004	:douta	=	16'h	4b72;
1005	:douta	=	16'h	4374;
1006	:douta	=	16'h	8517;
1007	:douta	=	16'h	8d18;
1008	:douta	=	16'h	4b51;
1009	:douta	=	16'h	63f5;
1010	:douta	=	16'h	11ed;
1011	:douta	=	16'h	6435;
1012	:douta	=	16'h	5bd4;
1013	:douta	=	16'h	ae1c;
1014	:douta	=	16'h	9e1d;
1015	:douta	=	16'h	5c15;
1016	:douta	=	16'h	5c38;
1017	:douta	=	16'h	32d2;
1018	:douta	=	16'h	3ad2;
1019	:douta	=	16'h	53d5;
1020	:douta	=	16'h	5bb2;
1021	:douta	=	16'h	74d9;
1022	:douta	=	16'h	6436;
1023	:douta	=	16'h	5bf7;
1024	:douta	=	16'h	2a6f;
1025	:douta	=	16'h	3af1;
1026	:douta	=	16'h	32d1;
1027	:douta	=	16'h	4353;
1028	:douta	=	16'h	4b53;
1029	:douta	=	16'h	74b8;
1030	:douta	=	16'h	7cf9;
1031	:douta	=	16'h	7d3b;
1032	:douta	=	16'h	5352;
1033	:douta	=	16'h	4b10;
1034	:douta	=	16'h	7c56;
1035	:douta	=	16'h	7434;
1036	:douta	=	16'h	7435;
1037	:douta	=	16'h	a558;
1038	:douta	=	16'h	8d18;
1039	:douta	=	16'h	84b7;
1040	:douta	=	16'h	94d6;
1041	:douta	=	16'h	be3a;
1042	:douta	=	16'h	428e;
1043	:douta	=	16'h	6b91;
1044	:douta	=	16'h	a536;
1045	:douta	=	16'h	7413;
1046	:douta	=	16'h	94d6;
1047	:douta	=	16'h	ce38;
1048	:douta	=	16'h	adb8;
1049	:douta	=	16'h	d69b;
1050	:douta	=	16'h	7476;
1051	:douta	=	16'h	7c34;
1052	:douta	=	16'h	7455;
1053	:douta	=	16'h	73f3;
1054	:douta	=	16'h	8cd6;
1055	:douta	=	16'h	84b6;
1056	:douta	=	16'h	9516;
1057	:douta	=	16'h	c619;
1058	:douta	=	16'h	ef3c;
1059	:douta	=	16'h	ef5b;
1060	:douta	=	16'h	9d58;
1061	:douta	=	16'h	ad56;
1062	:douta	=	16'h	7cd7;
1063	:douta	=	16'h	6bb3;
1064	:douta	=	16'h	b5b8;
1065	:douta	=	16'h	8454;
1066	:douta	=	16'h	ce59;
1067	:douta	=	16'h	deba;
1068	:douta	=	16'h	e6da;
1069	:douta	=	16'h	c5f8;
1070	:douta	=	16'h	7475;
1071	:douta	=	16'h	7c12;
1072	:douta	=	16'h	c619;
1073	:douta	=	16'h	6371;
1074	:douta	=	16'h	8494;
1075	:douta	=	16'h	de58;
1076	:douta	=	16'h	ded9;
1077	:douta	=	16'h	bdd7;
1078	:douta	=	16'h	d6da;
1079	:douta	=	16'h	9cf7;
1080	:douta	=	16'h	8c93;
1081	:douta	=	16'h	a514;
1082	:douta	=	16'h	94f5;
1083	:douta	=	16'h	84b5;
1084	:douta	=	16'h	8474;
1085	:douta	=	16'h	f77b;
1086	:douta	=	16'h	e71b;
1087	:douta	=	16'h	ad98;
1088	:douta	=	16'h	6c36;
1089	:douta	=	16'h	3ad0;
1090	:douta	=	16'h	a4d4;
1091	:douta	=	16'h	b5f8;
1092	:douta	=	16'h	a577;
1093	:douta	=	16'h	7453;
1094	:douta	=	16'h	a556;
1095	:douta	=	16'h	deb9;
1096	:douta	=	16'h	9537;
1097	:douta	=	16'h	ff9c;
1098	:douta	=	16'h	63f4;
1099	:douta	=	16'h	6bf4;
1100	:douta	=	16'h	b5f9;
1101	:douta	=	16'h	4b72;
1102	:douta	=	16'h	9599;
1103	:douta	=	16'h	7bd0;
1104	:douta	=	16'h	ae19;
1105	:douta	=	16'h	9515;
1106	:douta	=	16'h	8cf6;
1107	:douta	=	16'h	be5b;
1108	:douta	=	16'h	adb8;
1109	:douta	=	16'h	d67b;
1110	:douta	=	16'h	9d98;
1111	:douta	=	16'h	7415;
1112	:douta	=	16'h	7477;
1113	:douta	=	16'h	7476;
1114	:douta	=	16'h	b5d8;
1115	:douta	=	16'h	7c74;
1116	:douta	=	16'h	c619;
1117	:douta	=	16'h	7477;
1118	:douta	=	16'h	b5f9;
1119	:douta	=	16'h	be19;
1120	:douta	=	16'h	32b1;
1121	:douta	=	16'h	7bf3;
1122	:douta	=	16'h	11ce;
1123	:douta	=	16'h	4b74;
1124	:douta	=	16'h	a596;
1125	:douta	=	16'h	5b93;
1126	:douta	=	16'h	bdd8;
1127	:douta	=	16'h	9dda;
1128	:douta	=	16'h	9518;
1129	:douta	=	16'h	6c77;
1130	:douta	=	16'h	defc;
1131	:douta	=	16'h	74f8;
1132	:douta	=	16'h	4b53;
1133	:douta	=	16'h	6414;
1134	:douta	=	16'h	6c55;
1135	:douta	=	16'h	9538;
1136	:douta	=	16'h	5bd5;
1137	:douta	=	16'h	c65b;
1138	:douta	=	16'h	e71b;
1139	:douta	=	16'h	9518;
1140	:douta	=	16'h	63d2;
1141	:douta	=	16'h	63b2;
1142	:douta	=	16'h	7c12;
1143	:douta	=	16'h	9d77;
1144	:douta	=	16'h	8473;
1145	:douta	=	16'h	6bd3;
1146	:douta	=	16'h	7c74;
1147	:douta	=	16'h	bdd7;
1148	:douta	=	16'h	ff7c;
1149	:douta	=	16'h	a598;
1150	:douta	=	16'h	5bf5;
1151	:douta	=	16'h	42d0;
1152	:douta	=	16'h	324e;
1153	:douta	=	16'h	5350;
1154	:douta	=	16'h	426d;
1155	:douta	=	16'h	ad96;
1156	:douta	=	16'h	8c94;
1157	:douta	=	16'h	8cb4;
1158	:douta	=	16'h	b596;
1159	:douta	=	16'h	632e;
1160	:douta	=	16'h	8474;
1161	:douta	=	16'h	42cf;
1162	:douta	=	16'h	52ec;
1163	:douta	=	16'h	5b4e;
1164	:douta	=	16'h	9cf3;
1165	:douta	=	16'h	ce78;
1166	:douta	=	16'h	8472;
1167	:douta	=	16'h	c5d6;
1168	:douta	=	16'h	7c31;
1169	:douta	=	16'h	ad15;
1170	:douta	=	16'h	0907;
1171	:douta	=	16'h	4a6a;
1172	:douta	=	16'h	9450;
1173	:douta	=	16'h	ad33;
1174	:douta	=	16'h	a470;
1175	:douta	=	16'h	9471;
1176	:douta	=	16'h	3a0b;
1177	:douta	=	16'h	9430;
1178	:douta	=	16'h	632e;
1179	:douta	=	16'h	8c50;
1180	:douta	=	16'h	3a0a;
1181	:douta	=	16'h	5b2e;
1182	:douta	=	16'h	7c31;
1183	:douta	=	16'h	7c11;
1184	:douta	=	16'h	ce77;
1185	:douta	=	16'h	6b8f;
1186	:douta	=	16'h	acf3;
1187	:douta	=	16'h	7c10;
1188	:douta	=	16'h	634f;
1189	:douta	=	16'h	428e;
1190	:douta	=	16'h	4aad;
1191	:douta	=	16'h	29ea;
1192	:douta	=	16'h	2187;
1193	:douta	=	16'h	7c31;
1194	:douta	=	16'h	6b8f;
1195	:douta	=	16'h	94d4;
1196	:douta	=	16'h	e6d8;
1197	:douta	=	16'h	5331;
1198	:douta	=	16'h	630d;
1199	:douta	=	16'h	9d16;
1200	:douta	=	16'h	6414;
1201	:douta	=	16'h	5b2f;
1202	:douta	=	16'h	0884;
1203	:douta	=	16'h	0043;
1204	:douta	=	16'h	5b2f;
1205	:douta	=	16'h	1128;
1206	:douta	=	16'h	8450;
1207	:douta	=	16'h	9cb2;
1208	:douta	=	16'h	c5b4;
1209	:douta	=	16'h	6350;
1210	:douta	=	16'h	9cd2;
1211	:douta	=	16'h	18c4;
1212	:douta	=	16'h	10c5;
1213	:douta	=	16'h	10c4;
1214	:douta	=	16'h	1926;
1215	:douta	=	16'h	1949;
1216	:douta	=	16'h	1149;
1217	:douta	=	16'h	a555;
1218	:douta	=	16'h	9d15;
1219	:douta	=	16'h	73d1;
1220	:douta	=	16'h	9493;
1221	:douta	=	16'h	8c52;
1222	:douta	=	16'h	4aae;
1223	:douta	=	16'h	5b4f;
1224	:douta	=	16'h	29a9;
1225	:douta	=	16'h	3a6c;
1226	:douta	=	16'h	9d14;
1227	:douta	=	16'h	6bd1;
1228	:douta	=	16'h	5b70;
1229	:douta	=	16'h	ad55;
1230	:douta	=	16'h	7c55;
1231	:douta	=	16'h	63d3;
1232	:douta	=	16'h	21cb;
1233	:douta	=	16'h	6370;
1234	:douta	=	16'h	ce58;
1235	:douta	=	16'h	9d37;
1236	:douta	=	16'h	de9a;
1237	:douta	=	16'h	74f9;
1238	:douta	=	16'h	6415;
1239	:douta	=	16'h	9d59;
1240	:douta	=	16'h	4b74;
1241	:douta	=	16'h	32d1;
1242	:douta	=	16'h	5373;
1243	:douta	=	16'h	7414;
1244	:douta	=	16'h	9d37;
1245	:douta	=	16'h	ad97;
1246	:douta	=	16'h	adda;
1247	:douta	=	16'h	52d0;
1248	:douta	=	16'h	84b7;
1249	:douta	=	16'h	3ad1;
1250	:douta	=	16'h	328f;
1251	:douta	=	16'h	222f;
1252	:douta	=	16'h	4353;
1253	:douta	=	16'h	2ab1;
1254	:douta	=	16'h	a5ba;
1255	:douta	=	16'h	9d79;
1256	:douta	=	16'h	84b7;
1257	:douta	=	16'h	63d3;
1258	:douta	=	16'h	6c77;
1259	:douta	=	16'h	3b53;
1260	:douta	=	16'h	53f7;
1261	:douta	=	16'h	4353;
1262	:douta	=	16'h	63d2;
1263	:douta	=	16'h	84f7;
1264	:douta	=	16'h	bdfa;
1265	:douta	=	16'h	959c;
1266	:douta	=	16'h	63f4;
1267	:douta	=	16'h	3af1;
1268	:douta	=	16'h	4311;
1269	:douta	=	16'h	3b33;
1270	:douta	=	16'h	3b74;
1271	:douta	=	16'h	a5da;
1272	:douta	=	16'h	53d6;
1273	:douta	=	16'h	7c97;
1274	:douta	=	16'h	6479;
1275	:douta	=	16'h	32f3;
1276	:douta	=	16'h	4b73;
1277	:douta	=	16'h	4b74;
1278	:douta	=	16'h	9559;
1279	:douta	=	16'h	53f6;
1280	:douta	=	16'h	7cfa;
1281	:douta	=	16'h	3b12;
1282	:douta	=	16'h	4b53;
1283	:douta	=	16'h	3b12;
1284	:douta	=	16'h	2a4e;
1285	:douta	=	16'h	32b0;
1286	:douta	=	16'h	7455;
1287	:douta	=	16'h	5bd5;
1288	:douta	=	16'h	63b3;
1289	:douta	=	16'h	6bf3;
1290	:douta	=	16'h	7455;
1291	:douta	=	16'h	6bf4;
1292	:douta	=	16'h	7c55;
1293	:douta	=	16'h	5372;
1294	:douta	=	16'h	7c13;
1295	:douta	=	16'h	6392;
1296	:douta	=	16'h	a577;
1297	:douta	=	16'h	bdf9;
1298	:douta	=	16'h	ad56;
1299	:douta	=	16'h	b5d9;
1300	:douta	=	16'h	7c76;
1301	:douta	=	16'h	a5ba;
1302	:douta	=	16'h	4312;
1303	:douta	=	16'h	94b6;
1304	:douta	=	16'h	8475;
1305	:douta	=	16'h	a557;
1306	:douta	=	16'h	7414;
1307	:douta	=	16'h	94b4;
1308	:douta	=	16'h	f77c;
1309	:douta	=	16'h	b5d9;
1310	:douta	=	16'h	e6b9;
1311	:douta	=	16'h	7476;
1312	:douta	=	16'h	94f6;
1313	:douta	=	16'h	94d5;
1314	:douta	=	16'h	5b93;
1315	:douta	=	16'h	7413;
1316	:douta	=	16'h	7413;
1317	:douta	=	16'h	adb8;
1318	:douta	=	16'h	defa;
1319	:douta	=	16'h	de79;
1320	:douta	=	16'h	ff7b;
1321	:douta	=	16'h	8cd6;
1322	:douta	=	16'h	8454;
1323	:douta	=	16'h	94d4;
1324	:douta	=	16'h	5330;
1325	:douta	=	16'h	de99;
1326	:douta	=	16'h	8c96;
1327	:douta	=	16'h	bdf8;
1328	:douta	=	16'h	c659;
1329	:douta	=	16'h	de79;
1330	:douta	=	16'h	be3a;
1331	:douta	=	16'h	6371;
1332	:douta	=	16'h	ad36;
1333	:douta	=	16'h	6370;
1334	:douta	=	16'h	84d5;
1335	:douta	=	16'h	7413;
1336	:douta	=	16'h	defa;
1337	:douta	=	16'h	ff7b;
1338	:douta	=	16'h	94d4;
1339	:douta	=	16'h	c6bb;
1340	:douta	=	16'h	53d4;
1341	:douta	=	16'h	b596;
1342	:douta	=	16'h	c67a;
1343	:douta	=	16'h	8c94;
1344	:douta	=	16'h	7c13;
1345	:douta	=	16'h	9d56;
1346	:douta	=	16'h	ff5b;
1347	:douta	=	16'h	e73c;
1348	:douta	=	16'h	d618;
1349	:douta	=	16'h	6c54;
1350	:douta	=	16'h	5b0f;
1351	:douta	=	16'h	c619;
1352	:douta	=	16'h	6bd2;
1353	:douta	=	16'h	9d58;
1354	:douta	=	16'h	6414;
1355	:douta	=	16'h	b5b8;
1356	:douta	=	16'h	b619;
1357	:douta	=	16'h	ce18;
1358	:douta	=	16'h	8d57;
1359	:douta	=	16'h	ce17;
1360	:douta	=	16'h	7bd3;
1361	:douta	=	16'h	defa;
1362	:douta	=	16'h	95bb;
1363	:douta	=	16'h	63b3;
1364	:douta	=	16'h	63d3;
1365	:douta	=	16'h	7c33;
1366	:douta	=	16'h	8495;
1367	:douta	=	16'h	c638;
1368	:douta	=	16'h	b619;
1369	:douta	=	16'h	ce39;
1370	:douta	=	16'h	b63a;
1371	:douta	=	16'h	d65b;
1372	:douta	=	16'h	a5fa;
1373	:douta	=	16'h	3aaf;
1374	:douta	=	16'h	5332;
1375	:douta	=	16'h	a5b8;
1376	:douta	=	16'h	9537;
1377	:douta	=	16'h	ce7a;
1378	:douta	=	16'h	8d39;
1379	:douta	=	16'h	adb9;
1380	:douta	=	16'h	e71d;
1381	:douta	=	16'h	63d4;
1382	:douta	=	16'h	a537;
1383	:douta	=	16'h	2a6f;
1384	:douta	=	16'h	9cd5;
1385	:douta	=	16'h	63f4;
1386	:douta	=	16'h	e73c;
1387	:douta	=	16'h	9579;
1388	:douta	=	16'h	959b;
1389	:douta	=	16'h	ce7b;
1390	:douta	=	16'h	8d59;
1391	:douta	=	16'h	be3a;
1392	:douta	=	16'h	6476;
1393	:douta	=	16'h	bdb8;
1394	:douta	=	16'h	a599;
1395	:douta	=	16'h	5b93;
1396	:douta	=	16'h	63f3;
1397	:douta	=	16'h	5bb2;
1398	:douta	=	16'h	e6da;
1399	:douta	=	16'h	b65a;
1400	:douta	=	16'h	b575;
1401	:douta	=	16'h	3aae;
1402	:douta	=	16'h	198a;
1403	:douta	=	16'h	9515;
1404	:douta	=	16'h	84f5;
1405	:douta	=	16'h	8cb6;
1406	:douta	=	16'h	7455;
1407	:douta	=	16'h	7c95;
1408	:douta	=	16'h	ffbc;
1409	:douta	=	16'h	b619;
1410	:douta	=	16'h	5ace;
1411	:douta	=	16'h	7c13;
1412	:douta	=	16'h	1969;
1413	:douta	=	16'h	634f;
1414	:douta	=	16'h	534f;
1415	:douta	=	16'h	63af;
1416	:douta	=	16'h	b5d6;
1417	:douta	=	16'h	a533;
1418	:douta	=	16'h	ce57;
1419	:douta	=	16'h	73d0;
1420	:douta	=	16'h	62ec;
1421	:douta	=	16'h	3a2c;
1422	:douta	=	16'h	21a9;
1423	:douta	=	16'h	6b90;
1424	:douta	=	16'h	a513;
1425	:douta	=	16'h	bd95;
1426	:douta	=	16'h	9c70;
1427	:douta	=	16'h	8bf0;
1428	:douta	=	16'h	9d13;
1429	:douta	=	16'h	4a8c;
1430	:douta	=	16'h	73ae;
1431	:douta	=	16'h	636e;
1432	:douta	=	16'h	8430;
1433	:douta	=	16'h	adb5;
1434	:douta	=	16'h	a513;
1435	:douta	=	16'h	ad35;
1436	:douta	=	16'h	4a6b;
1437	:douta	=	16'h	9c0f;
1438	:douta	=	16'h	3a4c;
1439	:douta	=	16'h	1905;
1440	:douta	=	16'h	4a6b;
1441	:douta	=	16'h	422a;
1442	:douta	=	16'h	8c71;
1443	:douta	=	16'h	94d4;
1444	:douta	=	16'h	ad76;
1445	:douta	=	16'h	8c94;
1446	:douta	=	16'h	73f1;
1447	:douta	=	16'h	6b90;
1448	:douta	=	16'h	7bf1;
1449	:douta	=	16'h	3a2b;
1450	:douta	=	16'h	2169;
1451	:douta	=	16'h	31ca;
1452	:douta	=	16'h	3af0;
1453	:douta	=	16'h	5b6f;
1454	:douta	=	16'h	c617;
1455	:douta	=	16'h	8473;
1456	:douta	=	16'h	530f;
1457	:douta	=	16'h	ce78;
1458	:douta	=	16'h	73f2;
1459	:douta	=	16'h	e658;
1460	:douta	=	16'h	5bb1;
1461	:douta	=	16'h	3a0b;
1462	:douta	=	16'h	428d;
1463	:douta	=	16'h	326c;
1464	:douta	=	16'h	21ca;
1465	:douta	=	16'h	5b2e;
1466	:douta	=	16'h	a533;
1467	:douta	=	16'h	18a3;
1468	:douta	=	16'h	10c4;
1469	:douta	=	16'h	10c4;
1470	:douta	=	16'h	2967;
1471	:douta	=	16'h	94b4;
1472	:douta	=	16'h	2989;
1473	:douta	=	16'h	29ca;
1474	:douta	=	16'h	29cb;
1475	:douta	=	16'h	8453;
1476	:douta	=	16'h	638f;
1477	:douta	=	16'h	636f;
1478	:douta	=	16'h	9d14;
1479	:douta	=	16'h	8452;
1480	:douta	=	16'h	9472;
1481	:douta	=	16'h	73f3;
1482	:douta	=	16'h	5b2f;
1483	:douta	=	16'h	21aa;
1484	:douta	=	16'h	1107;
1485	:douta	=	16'h	8493;
1486	:douta	=	16'h	ad55;
1487	:douta	=	16'h	7c34;
1488	:douta	=	16'h	8452;
1489	:douta	=	16'h	ce59;
1490	:douta	=	16'h	4b93;
1491	:douta	=	16'h	7414;
1492	:douta	=	16'h	32b1;
1493	:douta	=	16'h	2a2d;
1494	:douta	=	16'h	6bd2;
1495	:douta	=	16'h	a578;
1496	:douta	=	16'h	cebb;
1497	:douta	=	16'h	6456;
1498	:douta	=	16'h	6bf4;
1499	:douta	=	16'h	63f4;
1500	:douta	=	16'h	63f4;
1501	:douta	=	16'h	4b72;
1502	:douta	=	16'h	32d0;
1503	:douta	=	16'h	6412;
1504	:douta	=	16'h	a5d9;
1505	:douta	=	16'h	9d57;
1506	:douta	=	16'h	9558;
1507	:douta	=	16'h	7414;
1508	:douta	=	16'h	7477;
1509	:douta	=	16'h	7498;
1510	:douta	=	16'h	3b11;
1511	:douta	=	16'h	2250;
1512	:douta	=	16'h	32f1;
1513	:douta	=	16'h	6c35;
1514	:douta	=	16'h	a599;
1515	:douta	=	16'h	a59a;
1516	:douta	=	16'h	6c56;
1517	:douta	=	16'h	6435;
1518	:douta	=	16'h	21cd;
1519	:douta	=	16'h	2a2e;
1520	:douta	=	16'h	1a4f;
1521	:douta	=	16'h	19ed;
1522	:douta	=	16'h	9559;
1523	:douta	=	16'h	8d18;
1524	:douta	=	16'h	8d18;
1525	:douta	=	16'h	6499;
1526	:douta	=	16'h	4354;
1527	:douta	=	16'h	5c16;
1528	:douta	=	16'h	5bf5;
1529	:douta	=	16'h	6c77;
1530	:douta	=	16'h	4375;
1531	:douta	=	16'h	6c35;
1532	:douta	=	16'h	6cb9;
1533	:douta	=	16'h	53d6;
1534	:douta	=	16'h	2290;
1535	:douta	=	16'h	1a2e;
1536	:douta	=	16'h	4b73;
1537	:douta	=	16'h	4312;
1538	:douta	=	16'h	5bd4;
1539	:douta	=	16'h	6458;
1540	:douta	=	16'h	5373;
1541	:douta	=	16'h	6c77;
1542	:douta	=	16'h	7477;
1543	:douta	=	16'h	53b4;
1544	:douta	=	16'h	116a;
1545	:douta	=	16'h	6372;
1546	:douta	=	16'h	7c96;
1547	:douta	=	16'h	84b6;
1548	:douta	=	16'h	a579;
1549	:douta	=	16'h	8cd7;
1550	:douta	=	16'h	8495;
1551	:douta	=	16'h	9517;
1552	:douta	=	16'h	5b92;
1553	:douta	=	16'h	7475;
1554	:douta	=	16'h	ad56;
1555	:douta	=	16'h	a576;
1556	:douta	=	16'h	ad77;
1557	:douta	=	16'h	9538;
1558	:douta	=	16'h	6c36;
1559	:douta	=	16'h	8cf6;
1560	:douta	=	16'h	8433;
1561	:douta	=	16'h	ad76;
1562	:douta	=	16'h	63d3;
1563	:douta	=	16'h	42d0;
1564	:douta	=	16'h	9d36;
1565	:douta	=	16'h	9d15;
1566	:douta	=	16'h	c618;
1567	:douta	=	16'h	b5d9;
1568	:douta	=	16'h	a599;
1569	:douta	=	16'h	ef1c;
1570	:douta	=	16'h	9d36;
1571	:douta	=	16'h	bdd7;
1572	:douta	=	16'h	222e;
1573	:douta	=	16'h	5b31;
1574	:douta	=	16'h	add8;
1575	:douta	=	16'h	9d17;
1576	:douta	=	16'h	deda;
1577	:douta	=	16'h	d679;
1578	:douta	=	16'h	ce9a;
1579	:douta	=	16'h	b5b8;
1580	:douta	=	16'h	a516;
1581	:douta	=	16'h	d679;
1582	:douta	=	16'h	5392;
1583	:douta	=	16'h	8473;
1584	:douta	=	16'h	b5b7;
1585	:douta	=	16'h	deb9;
1586	:douta	=	16'h	d6b9;
1587	:douta	=	16'h	a4f5;
1588	:douta	=	16'h	f6fb;
1589	:douta	=	16'h	6bb2;
1590	:douta	=	16'h	8d16;
1591	:douta	=	16'h	2a8f;
1592	:douta	=	16'h	a576;
1593	:douta	=	16'h	ad97;
1594	:douta	=	16'h	b576;
1595	:douta	=	16'h	be59;
1596	:douta	=	16'h	a557;
1597	:douta	=	16'h	e6fa;
1598	:douta	=	16'h	be9a;
1599	:douta	=	16'h	8c53;
1600	:douta	=	16'h	5351;
1601	:douta	=	16'h	8434;
1602	:douta	=	16'h	ce37;
1603	:douta	=	16'h	c659;
1604	:douta	=	16'h	f77c;
1605	:douta	=	16'h	b5f9;
1606	:douta	=	16'h	9d15;
1607	:douta	=	16'h	be18;
1608	:douta	=	16'h	8495;
1609	:douta	=	16'h	b619;
1610	:douta	=	16'h	32d1;
1611	:douta	=	16'h	5bb3;
1612	:douta	=	16'h	8c95;
1613	:douta	=	16'h	9d57;
1614	:douta	=	16'h	a5d8;
1615	:douta	=	16'h	d679;
1616	:douta	=	16'h	e6fb;
1617	:douta	=	16'h	d6db;
1618	:douta	=	16'h	b5b9;
1619	:douta	=	16'h	8519;
1620	:douta	=	16'h	83f3;
1621	:douta	=	16'h	b5b7;
1622	:douta	=	16'h	5372;
1623	:douta	=	16'h	3a8f;
1624	:douta	=	16'h	84b6;
1625	:douta	=	16'h	ce9a;
1626	:douta	=	16'h	b5f8;
1627	:douta	=	16'h	ef1b;
1628	:douta	=	16'h	be9b;
1629	:douta	=	16'h	7c76;
1630	:douta	=	16'h	7c34;
1631	:douta	=	16'h	6415;
1632	:douta	=	16'h	4b0f;
1633	:douta	=	16'h	6c13;
1634	:douta	=	16'h	9578;
1635	:douta	=	16'h	a5da;
1636	:douta	=	16'h	84d6;
1637	:douta	=	16'h	ad98;
1638	:douta	=	16'h	d6bb;
1639	:douta	=	16'h	8496;
1640	:douta	=	16'h	c619;
1641	:douta	=	16'h	4af0;
1642	:douta	=	16'h	a5fb;
1643	:douta	=	16'h	5bf5;
1644	:douta	=	16'h	5353;
1645	:douta	=	16'h	94f6;
1646	:douta	=	16'h	84d7;
1647	:douta	=	16'h	be7b;
1648	:douta	=	16'h	6c77;
1649	:douta	=	16'h	ef3d;
1650	:douta	=	16'h	b65b;
1651	:douta	=	16'h	6393;
1652	:douta	=	16'h	21ab;
1653	:douta	=	16'h	1949;
1654	:douta	=	16'h	9d55;
1655	:douta	=	16'h	84b5;
1656	:douta	=	16'h	be18;
1657	:douta	=	16'h	8474;
1658	:douta	=	16'h	94b5;
1659	:douta	=	16'h	ce59;
1660	:douta	=	16'h	5bb2;
1661	:douta	=	16'h	7c94;
1662	:douta	=	16'h	322d;
1663	:douta	=	16'h	6bb3;
1664	:douta	=	16'h	9db8;
1665	:douta	=	16'h	7cb6;
1666	:douta	=	16'h	acd4;
1667	:douta	=	16'h	8473;
1668	:douta	=	16'h	5330;
1669	:douta	=	16'h	94b3;
1670	:douta	=	16'h	322b;
1671	:douta	=	16'h	632f;
1672	:douta	=	16'h	4aad;
1673	:douta	=	16'h	8471;
1674	:douta	=	16'h	8c72;
1675	:douta	=	16'h	a555;
1676	:douta	=	16'h	9cb3;
1677	:douta	=	16'h	52ee;
1678	:douta	=	16'h	630d;
1679	:douta	=	16'h	5b0e;
1680	:douta	=	16'h	73af;
1681	:douta	=	16'h	73af;
1682	:douta	=	16'h	736e;
1683	:douta	=	16'h	ad12;
1684	:douta	=	16'h	94b1;
1685	:douta	=	16'h	52ac;
1686	:douta	=	16'h	cdf5;
1687	:douta	=	16'h	1969;
1688	:douta	=	16'h	1107;
1689	:douta	=	16'h	6b90;
1690	:douta	=	16'h	9cd3;
1691	:douta	=	16'h	de99;
1692	:douta	=	16'h	9451;
1693	:douta	=	16'h	ff7b;
1694	:douta	=	16'h	530f;
1695	:douta	=	16'h	4a8d;
1696	:douta	=	16'h	6b8f;
1697	:douta	=	16'h	10e5;
1698	:douta	=	16'h	428b;
1699	:douta	=	16'h	5b6f;
1700	:douta	=	16'h	7c31;
1701	:douta	=	16'h	73d1;
1702	:douta	=	16'h	7c11;
1703	:douta	=	16'h	a514;
1704	:douta	=	16'h	5b0d;
1705	:douta	=	16'h	9453;
1706	:douta	=	16'h	39eb;
1707	:douta	=	16'h	9410;
1708	:douta	=	16'h	3a8e;
1709	:douta	=	16'h	29ea;
1710	:douta	=	16'h	530e;
1711	:douta	=	16'h	5b4f;
1712	:douta	=	16'h	8431;
1713	:douta	=	16'h	c618;
1714	:douta	=	16'h	73f1;
1715	:douta	=	16'h	ce36;
1716	:douta	=	16'h	5b71;
1717	:douta	=	16'h	9451;
1718	:douta	=	16'h	5b51;
1719	:douta	=	16'h	6bb1;
1720	:douta	=	16'h	320c;
1721	:douta	=	16'h	52cd;
1722	:douta	=	16'h	8472;
1723	:douta	=	16'h	18e4;
1724	:douta	=	16'h	10c4;
1725	:douta	=	16'h	10c4;
1726	:douta	=	16'h	29c8;
1727	:douta	=	16'h	94d2;
1728	:douta	=	16'h	8451;
1729	:douta	=	16'h	428d;
1730	:douta	=	16'h	52ce;
1731	:douta	=	16'h	5b51;
1732	:douta	=	16'h	1108;
1733	:douta	=	16'h	5b2f;
1734	:douta	=	16'h	6bd1;
1735	:douta	=	16'h	6b90;
1736	:douta	=	16'h	d636;
1737	:douta	=	16'h	6bb1;
1738	:douta	=	16'h	a555;
1739	:douta	=	16'h	52ef;
1740	:douta	=	16'h	9d15;
1741	:douta	=	16'h	218b;
1742	:douta	=	16'h	7411;
1743	:douta	=	16'h	322c;
1744	:douta	=	16'h	ad75;
1745	:douta	=	16'h	d69a;
1746	:douta	=	16'h	7c55;
1747	:douta	=	16'h	de9a;
1748	:douta	=	16'h	5c16;
1749	:douta	=	16'h	326d;
1750	:douta	=	16'h	4b31;
1751	:douta	=	16'h	84b5;
1752	:douta	=	16'h	7c95;
1753	:douta	=	16'h	63f5;
1754	:douta	=	16'h	ad77;
1755	:douta	=	16'h	9d58;
1756	:douta	=	16'h	9d58;
1757	:douta	=	16'h	84d9;
1758	:douta	=	16'h	3a8f;
1759	:douta	=	16'h	3290;
1760	:douta	=	16'h	19ee;
1761	:douta	=	16'h	3aaf;
1762	:douta	=	16'h	7c95;
1763	:douta	=	16'h	9536;
1764	:douta	=	16'h	adba;
1765	:douta	=	16'h	9d58;
1766	:douta	=	16'h	6cb9;
1767	:douta	=	16'h	32b1;
1768	:douta	=	16'h	6436;
1769	:douta	=	16'h	010b;
1770	:douta	=	16'h	3b53;
1771	:douta	=	16'h	4332;
1772	:douta	=	16'h	84f8;
1773	:douta	=	16'h	8d39;
1774	:douta	=	16'h	3b34;
1775	:douta	=	16'h	7455;
1776	:douta	=	16'h	222e;
1777	:douta	=	16'h	4b73;
1778	:douta	=	16'h	2a4f;
1779	:douta	=	16'h	a5b9;
1780	:douta	=	16'h	b65c;
1781	:douta	=	16'h	5c37;
1782	:douta	=	16'h	84b7;
1783	:douta	=	16'h	5c17;
1784	:douta	=	16'h	959b;
1785	:douta	=	16'h	4396;
1786	:douta	=	16'h	11ac;
1787	:douta	=	16'h	63f4;
1788	:douta	=	16'h	6c78;
1789	:douta	=	16'h	5c58;
1790	:douta	=	16'h	4355;
1791	:douta	=	16'h	5395;
1792	:douta	=	16'h	6c98;
1793	:douta	=	16'h	4bd6;
1794	:douta	=	16'h	5c17;
1795	:douta	=	16'h	4bf6;
1796	:douta	=	16'h	4b32;
1797	:douta	=	16'h	4b53;
1798	:douta	=	16'h	63d4;
1799	:douta	=	16'h	7cd8;
1800	:douta	=	16'h	6c56;
1801	:douta	=	16'h	6bd3;
1802	:douta	=	16'h	7c35;
1803	:douta	=	16'h	5351;
1804	:douta	=	16'h	4b31;
1805	:douta	=	16'h	6bd3;
1806	:douta	=	16'h	7c75;
1807	:douta	=	16'h	ad98;
1808	:douta	=	16'h	ce5a;
1809	:douta	=	16'h	d6bd;
1810	:douta	=	16'h	94f5;
1811	:douta	=	16'h	5bd3;
1812	:douta	=	16'h	428f;
1813	:douta	=	16'h	4332;
1814	:douta	=	16'h	3ad0;
1815	:douta	=	16'h	6bf1;
1816	:douta	=	16'h	c639;
1817	:douta	=	16'h	e6da;
1818	:douta	=	16'h	be3a;
1819	:douta	=	16'h	9d78;
1820	:douta	=	16'h	d6ba;
1821	:douta	=	16'h	9d79;
1822	:douta	=	16'h	a577;
1823	:douta	=	16'h	5372;
1824	:douta	=	16'h	6bd3;
1825	:douta	=	16'h	73f2;
1826	:douta	=	16'h	c639;
1827	:douta	=	16'h	e6da;
1828	:douta	=	16'h	9d36;
1829	:douta	=	16'h	eefa;
1830	:douta	=	16'h	ce7a;
1831	:douta	=	16'h	9495;
1832	:douta	=	16'h	e6bb;
1833	:douta	=	16'h	6bf3;
1834	:douta	=	16'h	7c54;
1835	:douta	=	16'h	ad97;
1836	:douta	=	16'h	eed9;
1837	:douta	=	16'h	eefa;
1838	:douta	=	16'h	a578;
1839	:douta	=	16'h	bdd8;
1840	:douta	=	16'h	ad98;
1841	:douta	=	16'h	8433;
1842	:douta	=	16'h	6bd2;
1843	:douta	=	16'h	7c53;
1844	:douta	=	16'h	a534;
1845	:douta	=	16'h	ad56;
1846	:douta	=	16'h	ce58;
1847	:douta	=	16'h	a4f5;
1848	:douta	=	16'h	f75a;
1849	:douta	=	16'h	bdf7;
1850	:douta	=	16'h	7bf0;
1851	:douta	=	16'h	6415;
1852	:douta	=	16'h	4312;
1853	:douta	=	16'h	ded9;
1854	:douta	=	16'h	deba;
1855	:douta	=	16'h	e73a;
1856	:douta	=	16'h	a557;
1857	:douta	=	16'h	7c55;
1858	:douta	=	16'h	f77d;
1859	:douta	=	16'h	5c36;
1860	:douta	=	16'h	9c93;
1861	:douta	=	16'h	220d;
1862	:douta	=	16'h	21ab;
1863	:douta	=	16'h	9515;
1864	:douta	=	16'h	bdd6;
1865	:douta	=	16'h	ce59;
1866	:douta	=	16'h	a578;
1867	:douta	=	16'h	ce7a;
1868	:douta	=	16'h	6c56;
1869	:douta	=	16'h	5b73;
1870	:douta	=	16'h	7495;
1871	:douta	=	16'h	63f3;
1872	:douta	=	16'h	426d;
1873	:douta	=	16'h	84f9;
1874	:douta	=	16'h	7474;
1875	:douta	=	16'h	a557;
1876	:douta	=	16'h	e6b9;
1877	:douta	=	16'h	ce9a;
1878	:douta	=	16'h	6bd3;
1879	:douta	=	16'h	eed9;
1880	:douta	=	16'h	53d5;
1881	:douta	=	16'h	4b11;
1882	:douta	=	16'h	5bb4;
1883	:douta	=	16'h	84f7;
1884	:douta	=	16'h	4b71;
1885	:douta	=	16'h	7cb6;
1886	:douta	=	16'h	ad98;
1887	:douta	=	16'h	8d38;
1888	:douta	=	16'h	d67a;
1889	:douta	=	16'h	be7c;
1890	:douta	=	16'h	32b0;
1891	:douta	=	16'h	7c14;
1892	:douta	=	16'h	7496;
1893	:douta	=	16'h	7c54;
1894	:douta	=	16'h	6414;
1895	:douta	=	16'h	7454;
1896	:douta	=	16'h	84b4;
1897	:douta	=	16'h	adb8;
1898	:douta	=	16'h	d6fb;
1899	:douta	=	16'h	6c98;
1900	:douta	=	16'h	df1d;
1901	:douta	=	16'h	df3e;
1902	:douta	=	16'h	8cf8;
1903	:douta	=	16'h	7434;
1904	:douta	=	16'h	63b4;
1905	:douta	=	16'h	8d59;
1906	:douta	=	16'h	84d7;
1907	:douta	=	16'h	9577;
1908	:douta	=	16'h	9517;
1909	:douta	=	16'h	b5f9;
1910	:douta	=	16'h	b5f8;
1911	:douta	=	16'h	5331;
1912	:douta	=	16'h	63b1;
1913	:douta	=	16'h	29aa;
1914	:douta	=	16'h	63b2;
1915	:douta	=	16'h	9536;
1916	:douta	=	16'h	7412;
1917	:douta	=	16'h	9d77;
1918	:douta	=	16'h	9d57;
1919	:douta	=	16'h	ad76;
1920	:douta	=	16'h	6c13;
1921	:douta	=	16'h	29cc;
1922	:douta	=	16'h	8c93;
1923	:douta	=	16'h	3a4c;
1924	:douta	=	16'h	3a8e;
1925	:douta	=	16'h	a597;
1926	:douta	=	16'h	5330;
1927	:douta	=	16'h	ef3a;
1928	:douta	=	16'h	3a4c;
1929	:douta	=	16'h	8bf0;
1930	:douta	=	16'h	4aac;
1931	:douta	=	16'h	0885;
1932	:douta	=	16'h	6b8e;
1933	:douta	=	16'h	b595;
1934	:douta	=	16'h	ce78;
1935	:douta	=	16'h	738f;
1936	:douta	=	16'h	cdf6;
1937	:douta	=	16'h	526b;
1938	:douta	=	16'h	944e;
1939	:douta	=	16'h	ce14;
1940	:douta	=	16'h	31ea;
1941	:douta	=	16'h	424a;
1942	:douta	=	16'h	638f;
1943	:douta	=	16'h	a512;
1944	:douta	=	16'h	e6b7;
1945	:douta	=	16'h	9431;
1946	:douta	=	16'h	b575;
1947	:douta	=	16'h	31ec;
1948	:douta	=	16'h	7bd0;
1949	:douta	=	16'h	428c;
1950	:douta	=	16'h	a4d3;
1951	:douta	=	16'h	ad75;
1952	:douta	=	16'h	73af;
1953	:douta	=	16'h	9c71;
1954	:douta	=	16'h	d698;
1955	:douta	=	16'h	8433;
1956	:douta	=	16'h	a516;
1957	:douta	=	16'h	1169;
1958	:douta	=	16'h	08a4;
1959	:douta	=	16'h	0063;
1960	:douta	=	16'h	73f1;
1961	:douta	=	16'h	7c32;
1962	:douta	=	16'h	8c52;
1963	:douta	=	16'h	a575;
1964	:douta	=	16'h	5b70;
1965	:douta	=	16'h	bd54;
1966	:douta	=	16'h	8453;
1967	:douta	=	16'h	21cb;
1968	:douta	=	16'h	322c;
1969	:douta	=	16'h	3a2c;
1970	:douta	=	16'h	5350;
1971	:douta	=	16'h	63f2;
1972	:douta	=	16'h	8454;
1973	:douta	=	16'h	7411;
1974	:douta	=	16'h	8c72;
1975	:douta	=	16'h	8473;
1976	:douta	=	16'h	5b2f;
1977	:douta	=	16'h	9471;
1978	:douta	=	16'h	94f5;
1979	:douta	=	16'h	18a3;
1980	:douta	=	16'h	08c4;
1981	:douta	=	16'h	10a4;
1982	:douta	=	16'h	1906;
1983	:douta	=	16'h	2189;
1984	:douta	=	16'h	6bb0;
1985	:douta	=	16'h	a514;
1986	:douta	=	16'h	b555;
1987	:douta	=	16'h	7c12;
1988	:douta	=	16'h	8453;
1989	:douta	=	16'h	3a2b;
1990	:douta	=	16'h	39e9;
1991	:douta	=	16'h	52cd;
1992	:douta	=	16'h	29ca;
1993	:douta	=	16'h	428c;
1994	:douta	=	16'h	530f;
1995	:douta	=	16'h	ff58;
1996	:douta	=	16'h	c5f6;
1997	:douta	=	16'h	9c93;
1998	:douta	=	16'h	a515;
1999	:douta	=	16'h	3a4c;
2000	:douta	=	16'h	5331;
2001	:douta	=	16'h	0129;
2002	:douta	=	16'h	b5d7;
2003	:douta	=	16'h	9d57;
2004	:douta	=	16'h	63b2;
2005	:douta	=	16'h	b598;
2006	:douta	=	16'h	5373;
2007	:douta	=	16'h	9539;
2008	:douta	=	16'h	32d2;
2009	:douta	=	16'h	63d3;
2010	:douta	=	16'h	224e;
2011	:douta	=	16'h	3aaf;
2012	:douta	=	16'h	84b4;
2013	:douta	=	16'h	42cf;
2014	:douta	=	16'h	be59;
2015	:douta	=	16'h	5bf5;
2016	:douta	=	16'h	2a2e;
2017	:douta	=	16'h	53b4;
2018	:douta	=	16'h	012b;
2019	:douta	=	16'h	3af0;
2020	:douta	=	16'h	4312;
2021	:douta	=	16'h	5bf5;
2022	:douta	=	16'h	6c56;
2023	:douta	=	16'h	c639;
2024	:douta	=	16'h	9518;
2025	:douta	=	16'h	53b4;
2026	:douta	=	16'h	5c16;
2027	:douta	=	16'h	32d2;
2028	:douta	=	16'h	222e;
2029	:douta	=	16'h	4b53;
2030	:douta	=	16'h	7c75;
2031	:douta	=	16'h	8d19;
2032	:douta	=	16'h	9538;
2033	:douta	=	16'h	9539;
2034	:douta	=	16'h	53f6;
2035	:douta	=	16'h	63f5;
2036	:douta	=	16'h	11ac;
2037	:douta	=	16'h	220d;
2038	:douta	=	16'h	2270;
2039	:douta	=	16'h	7497;
2040	:douta	=	16'h	8519;
2041	:douta	=	16'h	53f6;
2042	:douta	=	16'h	857c;
2043	:douta	=	16'h	5438;
2044	:douta	=	16'h	3312;
2045	:douta	=	16'h	2ab0;
2046	:douta	=	16'h	3ad0;
2047	:douta	=	16'h	a5da;
2048	:douta	=	16'h	6c78;
2049	:douta	=	16'h	5c57;
2050	:douta	=	16'h	74d9;
2051	:douta	=	16'h	43b5;
2052	:douta	=	16'h	4311;
2053	:douta	=	16'h	3af1;
2054	:douta	=	16'h	5bb3;
2055	:douta	=	16'h	5b94;
2056	:douta	=	16'h	5393;
2057	:douta	=	16'h	8cf8;
2058	:douta	=	16'h	9518;
2059	:douta	=	16'h	7c75;
2060	:douta	=	16'h	6bf4;
2061	:douta	=	16'h	42f0;
2062	:douta	=	16'h	6b92;
2063	:douta	=	16'h	84b7;
2064	:douta	=	16'h	94d6;
2065	:douta	=	16'h	7455;
2066	:douta	=	16'h	ce59;
2067	:douta	=	16'h	9d57;
2068	:douta	=	16'h	9d16;
2069	:douta	=	16'h	7cb6;
2070	:douta	=	16'h	63b2;
2071	:douta	=	16'h	5330;
2072	:douta	=	16'h	6bf3;
2073	:douta	=	16'h	a536;
2074	:douta	=	16'h	7cb6;
2075	:douta	=	16'h	8cd5;
2076	:douta	=	16'h	bdd8;
2077	:douta	=	16'h	c63a;
2078	:douta	=	16'h	ce18;
2079	:douta	=	16'h	7cb6;
2080	:douta	=	16'h	6bd2;
2081	:douta	=	16'h	5350;
2082	:douta	=	16'h	94f6;
2083	:douta	=	16'h	94d5;
2084	:douta	=	16'h	a576;
2085	:douta	=	16'h	c5f8;
2086	:douta	=	16'h	c679;
2087	:douta	=	16'h	de59;
2088	:douta	=	16'h	ff9b;
2089	:douta	=	16'h	7435;
2090	:douta	=	16'h	6bd3;
2091	:douta	=	16'h	8c95;
2092	:douta	=	16'h	d679;
2093	:douta	=	16'h	e6d9;
2094	:douta	=	16'h	9d15;
2095	:douta	=	16'h	de98;
2096	:douta	=	16'h	d6ba;
2097	:douta	=	16'h	e6b9;
2098	:douta	=	16'h	be58;
2099	:douta	=	16'h	6bb2;
2100	:douta	=	16'h	9493;
2101	:douta	=	16'h	5330;
2102	:douta	=	16'h	84b4;
2103	:douta	=	16'h	8c53;
2104	:douta	=	16'h	c657;
2105	:douta	=	16'h	deb8;
2106	:douta	=	16'h	ad55;
2107	:douta	=	16'h	959a;
2108	:douta	=	16'h	4313;
2109	:douta	=	16'h	ad96;
2110	:douta	=	16'h	9516;
2111	:douta	=	16'h	a534;
2112	:douta	=	16'h	9d16;
2113	:douta	=	16'h	c619;
2114	:douta	=	16'h	f7bd;
2115	:douta	=	16'h	7496;
2116	:douta	=	16'h	fefa;
2117	:douta	=	16'h	4331;
2118	:douta	=	16'h	2a2d;
2119	:douta	=	16'h	8433;
2120	:douta	=	16'h	9cd5;
2121	:douta	=	16'h	a598;
2122	:douta	=	16'h	9d58;
2123	:douta	=	16'h	ce59;
2124	:douta	=	16'h	add9;
2125	:douta	=	16'h	ad57;
2126	:douta	=	16'h	9558;
2127	:douta	=	16'h	42d0;
2128	:douta	=	16'h	9494;
2129	:douta	=	16'h	4395;
2130	:douta	=	16'h	3a6f;
2131	:douta	=	16'h	6414;
2132	:douta	=	16'h	def9;
2133	:douta	=	16'h	be39;
2134	:douta	=	16'h	c619;
2135	:douta	=	16'h	ffbb;
2136	:douta	=	16'h	63b4;
2137	:douta	=	16'h	bd97;
2138	:douta	=	16'h	6c76;
2139	:douta	=	16'h	9558;
2140	:douta	=	16'h	5bb3;
2141	:douta	=	16'h	7456;
2142	:douta	=	16'h	4b11;
2143	:douta	=	16'h	84f7;
2144	:douta	=	16'h	94d5;
2145	:douta	=	16'h	6c33;
2146	:douta	=	16'h	7476;
2147	:douta	=	16'h	b5b9;
2148	:douta	=	16'h	853a;
2149	:douta	=	16'h	ad57;
2150	:douta	=	16'h	84f7;
2151	:douta	=	16'h	9d37;
2152	:douta	=	16'h	6c34;
2153	:douta	=	16'h	5b92;
2154	:douta	=	16'h	a5fa;
2155	:douta	=	16'h	9559;
2156	:douta	=	16'h	9558;
2157	:douta	=	16'h	a5b9;
2158	:douta	=	16'h	be39;
2159	:douta	=	16'h	9538;
2160	:douta	=	16'h	7415;
2161	:douta	=	16'h	8517;
2162	:douta	=	16'h	5351;
2163	:douta	=	16'h	53d3;
2164	:douta	=	16'h	7413;
2165	:douta	=	16'h	8cb5;
2166	:douta	=	16'h	be18;
2167	:douta	=	16'h	ad56;
2168	:douta	=	16'h	7c75;
2169	:douta	=	16'h	8452;
2170	:douta	=	16'h	8c73;
2171	:douta	=	16'h	3aae;
2172	:douta	=	16'h	1128;
2173	:douta	=	16'h	5b50;
2174	:douta	=	16'h	7455;
2175	:douta	=	16'h	9d57;
2176	:douta	=	16'h	4312;
2177	:douta	=	16'h	4a8f;
2178	:douta	=	16'h	b596;
2179	:douta	=	16'h	3a2c;
2180	:douta	=	16'h	29eb;
2181	:douta	=	16'h	638f;
2182	:douta	=	16'h	3a2c;
2183	:douta	=	16'h	9d35;
2184	:douta	=	16'h	6b8f;
2185	:douta	=	16'h	b575;
2186	:douta	=	16'h	632e;
2187	:douta	=	16'h	83d0;
2188	:douta	=	16'h	6b6e;
2189	:douta	=	16'h	8451;
2190	:douta	=	16'h	3aab;
2191	:douta	=	16'h	4aab;
2192	:douta	=	16'h	8c90;
2193	:douta	=	16'h	630c;
2194	:douta	=	16'h	bd72;
2195	:douta	=	16'h	d614;
2196	:douta	=	16'h	7411;
2197	:douta	=	16'h	73b0;
2198	:douta	=	16'h	426d;
2199	:douta	=	16'h	634f;
2200	:douta	=	16'h	9513;
2201	:douta	=	16'h	ad34;
2202	:douta	=	16'h	ded9;
2203	:douta	=	16'h	634f;
2204	:douta	=	16'h	a514;
2205	:douta	=	16'h	322b;
2206	:douta	=	16'h	6b8f;
2207	:douta	=	16'h	63af;
2208	:douta	=	16'h	6b8f;
2209	:douta	=	16'h	ce36;
2210	:douta	=	16'h	a555;
2211	:douta	=	16'h	8c53;
2212	:douta	=	16'h	8c73;
2213	:douta	=	16'h	3a2c;
2214	:douta	=	16'h	39e9;
2215	:douta	=	16'h	4a6b;
2216	:douta	=	16'h	1128;
2217	:douta	=	16'h	3a4c;
2218	:douta	=	16'h	6370;
2219	:douta	=	16'h	7c32;
2220	:douta	=	16'h	6370;
2221	:douta	=	16'h	ff7a;
2222	:douta	=	16'h	94d4;
2223	:douta	=	16'h	52ee;
2224	:douta	=	16'h	734f;
2225	:douta	=	16'h	42af;
2226	:douta	=	16'h	5b51;
2227	:douta	=	16'h	2a0d;
2228	:douta	=	16'h	6390;
2229	:douta	=	16'h	4aef;
2230	:douta	=	16'h	c638;
2231	:douta	=	16'h	6b90;
2232	:douta	=	16'h	6bb1;
2233	:douta	=	16'h	e656;
2234	:douta	=	16'h	ad35;
2235	:douta	=	16'h	18c3;
2236	:douta	=	16'h	10e4;
2237	:douta	=	16'h	10a4;
2238	:douta	=	16'h	2168;
2239	:douta	=	16'h	1106;
2240	:douta	=	16'h	218a;
2241	:douta	=	16'h	8c51;
2242	:douta	=	16'h	a534;
2243	:douta	=	16'h	7c33;
2244	:douta	=	16'h	8c94;
2245	:douta	=	16'h	6370;
2246	:douta	=	16'h	7bf0;
2247	:douta	=	16'h	634f;
2248	:douta	=	16'h	00e6;
2249	:douta	=	16'h	1148;
2250	:douta	=	16'h	21ca;
2251	:douta	=	16'h	6c10;
2252	:douta	=	16'h	73f1;
2253	:douta	=	16'h	ce37;
2254	:douta	=	16'h	bdb6;
2255	:douta	=	16'h	b534;
2256	:douta	=	16'h	8c94;
2257	:douta	=	16'h	8c53;
2258	:douta	=	16'h	6c13;
2259	:douta	=	16'h	6bf4;
2260	:douta	=	16'h	42cf;
2261	:douta	=	16'h	9d16;
2262	:douta	=	16'h	a577;
2263	:douta	=	16'h	84b7;
2264	:douta	=	16'h	5b93;
2265	:douta	=	16'h	8495;
2266	:douta	=	16'h	2a91;
2267	:douta	=	16'h	5372;
2268	:douta	=	16'h	114a;
2269	:douta	=	16'h	220c;
2270	:douta	=	16'h	8cf6;
2271	:douta	=	16'h	7454;
2272	:douta	=	16'h	8c95;
2273	:douta	=	16'h	5394;
2274	:douta	=	16'h	6391;
2275	:douta	=	16'h	6458;
2276	:douta	=	16'h	5bd5;
2277	:douta	=	16'h	4b94;
2278	:douta	=	16'h	32f1;
2279	:douta	=	16'h	63f4;
2280	:douta	=	16'h	9538;
2281	:douta	=	16'h	8519;
2282	:douta	=	16'h	6499;
2283	:douta	=	16'h	2290;
2284	:douta	=	16'h	3aaf;
2285	:douta	=	16'h	222e;
2286	:douta	=	16'h	4333;
2287	:douta	=	16'h	4352;
2288	:douta	=	16'h	ce9a;
2289	:douta	=	16'h	be3b;
2290	:douta	=	16'h	5bb3;
2291	:douta	=	16'h	957b;
2292	:douta	=	16'h	4353;
2293	:douta	=	16'h	5373;
2294	:douta	=	16'h	3af2;
2295	:douta	=	16'h	32d1;
2296	:douta	=	16'h	5c36;
2297	:douta	=	16'h	4bb4;
2298	:douta	=	16'h	7cd8;
2299	:douta	=	16'h	6c36;
2300	:douta	=	16'h	5c58;
2301	:douta	=	16'h	224f;
2302	:douta	=	16'h	4b32;
2303	:douta	=	16'h	5bd5;
2304	:douta	=	16'h	4b53;
2305	:douta	=	16'h	53d5;
2306	:douta	=	16'h	326f;
2307	:douta	=	16'h	5436;
2308	:douta	=	16'h	3af1;
2309	:douta	=	16'h	53b4;
2310	:douta	=	16'h	7c77;
2311	:douta	=	16'h	84f8;
2312	:douta	=	16'h	8d19;
2313	:douta	=	16'h	3aaf;
2314	:douta	=	16'h	324d;
2315	:douta	=	16'h	6391;
2316	:douta	=	16'h	8495;
2317	:douta	=	16'h	7c56;
2318	:douta	=	16'h	c619;
2319	:douta	=	16'h	adfb;
2320	:douta	=	16'h	d65a;
2321	:douta	=	16'h	adda;
2322	:douta	=	16'h	7433;
2323	:douta	=	16'h	6b92;
2324	:douta	=	16'h	7413;
2325	:douta	=	16'h	a578;
2326	:douta	=	16'h	9516;
2327	:douta	=	16'h	ce59;
2328	:douta	=	16'h	c639;
2329	:douta	=	16'h	c618;
2330	:douta	=	16'h	6c55;
2331	:douta	=	16'h	63d3;
2332	:douta	=	16'h	8495;
2333	:douta	=	16'h	a536;
2334	:douta	=	16'h	ad56;
2335	:douta	=	16'h	a516;
2336	:douta	=	16'h	a537;
2337	:douta	=	16'h	d679;
2338	:douta	=	16'h	ad77;
2339	:douta	=	16'h	bdb7;
2340	:douta	=	16'h	9d16;
2341	:douta	=	16'h	b577;
2342	:douta	=	16'h	94d5;
2343	:douta	=	16'h	7c95;
2344	:douta	=	16'h	94f6;
2345	:douta	=	16'h	ce18;
2346	:douta	=	16'h	d69a;
2347	:douta	=	16'h	ce38;
2348	:douta	=	16'h	e6b9;
2349	:douta	=	16'h	d698;
2350	:douta	=	16'h	7c33;
2351	:douta	=	16'h	8c93;
2352	:douta	=	16'h	8494;
2353	:douta	=	16'h	8c73;
2354	:douta	=	16'h	8474;
2355	:douta	=	16'h	e6d9;
2356	:douta	=	16'h	d698;
2357	:douta	=	16'h	ce58;
2358	:douta	=	16'h	add7;
2359	:douta	=	16'h	7433;
2360	:douta	=	16'h	e699;
2361	:douta	=	16'h	add7;
2362	:douta	=	16'h	428e;
2363	:douta	=	16'h	8c93;
2364	:douta	=	16'h	c5f6;
2365	:douta	=	16'h	f77a;
2366	:douta	=	16'h	be38;
2367	:douta	=	16'h	ce17;
2368	:douta	=	16'h	7414;
2369	:douta	=	16'h	3ab0;
2370	:douta	=	16'h	94f4;
2371	:douta	=	16'h	7474;
2372	:douta	=	16'h	ef7a;
2373	:douta	=	16'h	9d37;
2374	:douta	=	16'h	cdf9;
2375	:douta	=	16'h	ad97;
2376	:douta	=	16'h	d69a;
2377	:douta	=	16'h	b619;
2378	:douta	=	16'h	7c13;
2379	:douta	=	16'h	a576;
2380	:douta	=	16'h	4b73;
2381	:douta	=	16'h	94d4;
2382	:douta	=	16'h	6c34;
2383	:douta	=	16'h	d69a;
2384	:douta	=	16'h	e73c;
2385	:douta	=	16'h	9d79;
2386	:douta	=	16'h	de78;
2387	:douta	=	16'h	6436;
2388	:douta	=	16'h	d659;
2389	:douta	=	16'h	8d58;
2390	:douta	=	16'h	5a8c;
2391	:douta	=	16'h	94f6;
2392	:douta	=	16'h	b5d9;
2393	:douta	=	16'h	9db8;
2394	:douta	=	16'h	8d17;
2395	:douta	=	16'h	c69b;
2396	:douta	=	16'h	5bd5;
2397	:douta	=	16'h	add9;
2398	:douta	=	16'h	c5f8;
2399	:douta	=	16'h	5416;
2400	:douta	=	16'h	a5b9;
2401	:douta	=	16'h	7498;
2402	:douta	=	16'h	5372;
2403	:douta	=	16'h	4aaf;
2404	:douta	=	16'h	84d7;
2405	:douta	=	16'h	4352;
2406	:douta	=	16'h	63d4;
2407	:douta	=	16'h	a597;
2408	:douta	=	16'h	add9;
2409	:douta	=	16'h	de99;
2410	:douta	=	16'h	53b5;
2411	:douta	=	16'h	6bd4;
2412	:douta	=	16'h	84f8;
2413	:douta	=	16'h	5bb4;
2414	:douta	=	16'h	add8;
2415	:douta	=	16'h	a599;
2416	:douta	=	16'h	9558;
2417	:douta	=	16'h	9dba;
2418	:douta	=	16'h	9d79;
2419	:douta	=	16'h	adfa;
2420	:douta	=	16'h	9d37;
2421	:douta	=	16'h	8c33;
2422	:douta	=	16'h	7c74;
2423	:douta	=	16'h	1169;
2424	:douta	=	16'h	5330;
2425	:douta	=	16'h	9493;
2426	:douta	=	16'h	deba;
2427	:douta	=	16'h	8474;
2428	:douta	=	16'h	d67a;
2429	:douta	=	16'h	6391;
2430	:douta	=	16'h	6391;
2431	:douta	=	16'h	52ef;
2432	:douta	=	16'h	29ca;
2433	:douta	=	16'h	428d;
2434	:douta	=	16'h	9515;
2435	:douta	=	16'h	6bd2;
2436	:douta	=	16'h	a536;
2437	:douta	=	16'h	8474;
2438	:douta	=	16'h	defc;
2439	:douta	=	16'h	6bb1;
2440	:douta	=	16'h	8430;
2441	:douta	=	16'h	320a;
2442	:douta	=	16'h	422a;
2443	:douta	=	16'h	2987;
2444	:douta	=	16'h	52aa;
2445	:douta	=	16'h	20a2;
2446	:douta	=	16'h	18a3;
2447	:douta	=	16'h	0862;
2448	:douta	=	16'h	0000;
2449	:douta	=	16'h	2127;
2450	:douta	=	16'h	7c32;
2451	:douta	=	16'h	21a9;
2452	:douta	=	16'h	29a9;
2453	:douta	=	16'h	6baf;
2454	:douta	=	16'h	5b0e;
2455	:douta	=	16'h	8c94;
2456	:douta	=	16'h	5b0e;
2457	:douta	=	16'h	8c94;
2458	:douta	=	16'h	21aa;
2459	:douta	=	16'h	9cb3;
2460	:douta	=	16'h	52ec;
2461	:douta	=	16'h	6b4f;
2462	:douta	=	16'h	a514;
2463	:douta	=	16'h	73d1;
2464	:douta	=	16'h	bdd6;
2465	:douta	=	16'h	530f;
2466	:douta	=	16'h	94d4;
2467	:douta	=	16'h	ad76;
2468	:douta	=	16'h	bdf7;
2469	:douta	=	16'h	4aad;
2470	:douta	=	16'h	8431;
2471	:douta	=	16'h	8452;
2472	:douta	=	16'h	8453;
2473	:douta	=	16'h	6b90;
2474	:douta	=	16'h	6b70;
2475	:douta	=	16'h	8c94;
2476	:douta	=	16'h	4ace;
2477	:douta	=	16'h	42cf;
2478	:douta	=	16'h	8411;
2479	:douta	=	16'h	b596;
2480	:douta	=	16'h	ce99;
2481	:douta	=	16'h	b535;
2482	:douta	=	16'h	5bd2;
2483	:douta	=	16'h	428e;
2484	:douta	=	16'h	5b71;
2485	:douta	=	16'h	2a2b;
2486	:douta	=	16'h	4acf;
2487	:douta	=	16'h	6bb1;
2488	:douta	=	16'h	426d;
2489	:douta	=	16'h	3aae;
2490	:douta	=	16'h	5310;
2491	:douta	=	16'h	18a3;
2492	:douta	=	16'h	18e4;
2493	:douta	=	16'h	10c4;
2494	:douta	=	16'h	29c9;
2495	:douta	=	16'h	7412;
2496	:douta	=	16'h	424c;
2497	:douta	=	16'h	7c75;
2498	:douta	=	16'h	42af;
2499	:douta	=	16'h	29c9;
2500	:douta	=	16'h	220c;
2501	:douta	=	16'h	5b0f;
2502	:douta	=	16'h	c5f5;
2503	:douta	=	16'h	8c52;
2504	:douta	=	16'h	b596;
2505	:douta	=	16'h	8495;
2506	:douta	=	16'h	52cd;
2507	:douta	=	16'h	5b51;
2508	:douta	=	16'h	29eb;
2509	:douta	=	16'h	21ca;
2510	:douta	=	16'h	4b0f;
2511	:douta	=	16'h	7c73;
2512	:douta	=	16'h	94d4;
2513	:douta	=	16'h	bdd7;
2514	:douta	=	16'h	5372;
2515	:douta	=	16'h	5bd3;
2516	:douta	=	16'h	ad36;
2517	:douta	=	16'h	5b92;
2518	:douta	=	16'h	2a90;
2519	:douta	=	16'h	7c95;
2520	:douta	=	16'h	432f;
2521	:douta	=	16'h	9536;
2522	:douta	=	16'h	de58;
2523	:douta	=	16'h	9517;
2524	:douta	=	16'h	b5b8;
2525	:douta	=	16'h	9538;
2526	:douta	=	16'h	6c15;
2527	:douta	=	16'h	5373;
2528	:douta	=	16'h	4312;
2529	:douta	=	16'h	5bd4;
2530	:douta	=	16'h	8d18;
2531	:douta	=	16'h	b5fa;
2532	:douta	=	16'h	95bb;
2533	:douta	=	16'h	5c17;
2534	:douta	=	16'h	ae3c;
2535	:douta	=	16'h	6c99;
2536	:douta	=	16'h	4353;
2537	:douta	=	16'h	4bb5;
2538	:douta	=	16'h	53f5;
2539	:douta	=	16'h	84b5;
2540	:douta	=	16'h	a5da;
2541	:douta	=	16'h	8d5a;
2542	:douta	=	16'h	63d3;
2543	:douta	=	16'h	5b94;
2544	:douta	=	16'h	222f;
2545	:douta	=	16'h	19ce;
2546	:douta	=	16'h	53d3;
2547	:douta	=	16'h	326f;
2548	:douta	=	16'h	7434;
2549	:douta	=	16'h	7456;
2550	:douta	=	16'h	6437;
2551	:douta	=	16'h	7d1c;
2552	:douta	=	16'h	09ac;
2553	:douta	=	16'h	2ad1;
2554	:douta	=	16'h	3312;
2555	:douta	=	16'h	5c15;
2556	:douta	=	16'h	4394;
2557	:douta	=	16'h	ce59;
2558	:douta	=	16'h	7cb7;
2559	:douta	=	16'h	857b;
2560	:douta	=	16'h	6c78;
2561	:douta	=	16'h	6cb9;
2562	:douta	=	16'h	53d6;
2563	:douta	=	16'h	6478;
2564	:douta	=	16'h	4b53;
2565	:douta	=	16'h	4b52;
2566	:douta	=	16'h	5b93;
2567	:douta	=	16'h	7cb7;
2568	:douta	=	16'h	5393;
2569	:douta	=	16'h	7cb7;
2570	:douta	=	16'h	5311;
2571	:douta	=	16'h	63f4;
2572	:douta	=	16'h	4af1;
2573	:douta	=	16'h	3acf;
2574	:douta	=	16'h	8cb5;
2575	:douta	=	16'h	7c96;
2576	:douta	=	16'h	c639;
2577	:douta	=	16'h	a557;
2578	:douta	=	16'h	bdd9;
2579	:douta	=	16'h	9d16;
2580	:douta	=	16'h	7413;
2581	:douta	=	16'h	a578;
2582	:douta	=	16'h	6bf4;
2583	:douta	=	16'h	94b4;
2584	:douta	=	16'h	c5f8;
2585	:douta	=	16'h	ce59;
2586	:douta	=	16'h	9d58;
2587	:douta	=	16'h	bdd7;
2588	:douta	=	16'h	9d16;
2589	:douta	=	16'h	ad77;
2590	:douta	=	16'h	ad76;
2591	:douta	=	16'h	7c34;
2592	:douta	=	16'h	9cd4;
2593	:douta	=	16'h	b5f8;
2594	:douta	=	16'h	bdb6;
2595	:douta	=	16'h	c618;
2596	:douta	=	16'h	c639;
2597	:douta	=	16'h	e71b;
2598	:douta	=	16'h	ce5a;
2599	:douta	=	16'h	c619;
2600	:douta	=	16'h	9d58;
2601	:douta	=	16'h	7c53;
2602	:douta	=	16'h	73f1;
2603	:douta	=	16'h	adb8;
2604	:douta	=	16'h	ff9b;
2605	:douta	=	16'h	f75b;
2606	:douta	=	16'h	bdf8;
2607	:douta	=	16'h	e6b9;
2608	:douta	=	16'h	b5d8;
2609	:douta	=	16'h	8433;
2610	:douta	=	16'h	5bb2;
2611	:douta	=	16'h	6b91;
2612	:douta	=	16'h	9d35;
2613	:douta	=	16'h	8c93;
2614	:douta	=	16'h	ce59;
2615	:douta	=	16'h	ad35;
2616	:douta	=	16'h	ffdb;
2617	:douta	=	16'h	d6b9;
2618	:douta	=	16'h	9cb3;
2619	:douta	=	16'h	3acf;
2620	:douta	=	16'h	52ef;
2621	:douta	=	16'h	b596;
2622	:douta	=	16'h	a555;
2623	:douta	=	16'h	de78;
2624	:douta	=	16'h	ad77;
2625	:douta	=	16'h	9cb4;
2626	:douta	=	16'h	be39;
2627	:douta	=	16'h	6371;
2628	:douta	=	16'h	9d16;
2629	:douta	=	16'h	5bb2;
2630	:douta	=	16'h	6bb2;
2631	:douta	=	16'h	c618;
2632	:douta	=	16'h	b596;
2633	:douta	=	16'h	adb7;
2634	:douta	=	16'h	be3a;
2635	:douta	=	16'h	bdf8;
2636	:douta	=	16'h	6c56;
2637	:douta	=	16'h	a4f6;
2638	:douta	=	16'h	8517;
2639	:douta	=	16'h	4b31;
2640	:douta	=	16'h	5b70;
2641	:douta	=	16'h	6c34;
2642	:douta	=	16'h	bdf7;
2643	:douta	=	16'h	9d18;
2644	:douta	=	16'h	f77b;
2645	:douta	=	16'h	b61a;
2646	:douta	=	16'h	c5d8;
2647	:douta	=	16'h	d71c;
2648	:douta	=	16'h	63b4;
2649	:douta	=	16'h	8cd5;
2650	:douta	=	16'h	5372;
2651	:douta	=	16'h	8495;
2652	:douta	=	16'h	6c55;
2653	:douta	=	16'h	c618;
2654	:douta	=	16'h	e6fa;
2655	:douta	=	16'h	74b8;
2656	:douta	=	16'h	9d98;
2657	:douta	=	16'h	5bf6;
2658	:douta	=	16'h	3291;
2659	:douta	=	16'h	9cb4;
2660	:douta	=	16'h	6456;
2661	:douta	=	16'h	7434;
2662	:douta	=	16'h	3af1;
2663	:douta	=	16'h	6bd3;
2664	:douta	=	16'h	5bb3;
2665	:douta	=	16'h	ffdb;
2666	:douta	=	16'h	9599;
2667	:douta	=	16'h	6457;
2668	:douta	=	16'h	d69b;
2669	:douta	=	16'h	84d7;
2670	:douta	=	16'h	9d79;
2671	:douta	=	16'h	8cf6;
2672	:douta	=	16'h	9517;
2673	:douta	=	16'h	63f4;
2674	:douta	=	16'h	63b3;
2675	:douta	=	16'h	84d6;
2676	:douta	=	16'h	9d77;
2677	:douta	=	16'h	eefa;
2678	:douta	=	16'h	9d57;
2679	:douta	=	16'h	5b10;
2680	:douta	=	16'h	5370;
2681	:douta	=	16'h	9cb3;
2682	:douta	=	16'h	a5d7;
2683	:douta	=	16'h	52ee;
2684	:douta	=	16'h	94d5;
2685	:douta	=	16'h	a557;
2686	:douta	=	16'h	a557;
2687	:douta	=	16'h	a557;
2688	:douta	=	16'h	5b2f;
2689	:douta	=	16'h	6370;
2690	:douta	=	16'h	5b0f;
2691	:douta	=	16'h	6b90;
2692	:douta	=	16'h	532f;
2693	:douta	=	16'h	7c13;
2694	:douta	=	16'h	8495;
2695	:douta	=	16'h	8cb5;
2696	:douta	=	16'h	c658;
2697	:douta	=	16'h	6bd0;
2698	:douta	=	16'h	8c31;
2699	:douta	=	16'h	738e;
2700	:douta	=	16'h	0000;
2701	:douta	=	16'h	2924;
2702	:douta	=	16'h	18e3;
2703	:douta	=	16'h	0861;
2704	:douta	=	16'h	10e3;
2705	:douta	=	16'h	2188;
2706	:douta	=	16'h	5351;
2707	:douta	=	16'h	426d;
2708	:douta	=	16'h	3a2b;
2709	:douta	=	16'h	08a6;
2710	:douta	=	16'h	636f;
2711	:douta	=	16'h	3a0a;
2712	:douta	=	16'h	7c12;
2713	:douta	=	16'h	9d36;
2714	:douta	=	16'h	532f;
2715	:douta	=	16'h	b596;
2716	:douta	=	16'h	630e;
2717	:douta	=	16'h	8432;
2718	:douta	=	16'h	636f;
2719	:douta	=	16'h	3a2a;
2720	:douta	=	16'h	c617;
2721	:douta	=	16'h	8c72;
2722	:douta	=	16'h	bdb7;
2723	:douta	=	16'h	5b51;
2724	:douta	=	16'h	73f2;
2725	:douta	=	16'h	5b0d;
2726	:douta	=	16'h	29a9;
2727	:douta	=	16'h	29a8;
2728	:douta	=	16'h	532e;
2729	:douta	=	16'h	4aed;
2730	:douta	=	16'h	b5b6;
2731	:douta	=	16'h	8474;
2732	:douta	=	16'h	7bd0;
2733	:douta	=	16'h	428f;
2734	:douta	=	16'h	5b2f;
2735	:douta	=	16'h	6bf1;
2736	:douta	=	16'h	5bb1;
2737	:douta	=	16'h	bdf7;
2738	:douta	=	16'h	8c94;
2739	:douta	=	16'h	7bf2;
2740	:douta	=	16'h	8473;
2741	:douta	=	16'h	73f2;
2742	:douta	=	16'h	7454;
2743	:douta	=	16'h	2168;
2744	:douta	=	16'h	6b8f;
2745	:douta	=	16'h	6391;
2746	:douta	=	16'h	4af0;
2747	:douta	=	16'h	2124;
2748	:douta	=	16'h	10e4;
2749	:douta	=	16'h	10c4;
2750	:douta	=	16'h	39e9;
2751	:douta	=	16'h	9494;
2752	:douta	=	16'h	738f;
2753	:douta	=	16'h	7455;
2754	:douta	=	16'h	3ab0;
2755	:douta	=	16'h	7c33;
2756	:douta	=	16'h	3a6e;
2757	:douta	=	16'h	1107;
2758	:douta	=	16'h	4aee;
2759	:douta	=	16'h	4acd;
2760	:douta	=	16'h	c617;
2761	:douta	=	16'h	6b70;
2762	:douta	=	16'h	d615;
2763	:douta	=	16'h	5352;
2764	:douta	=	16'h	6bb2;
2765	:douta	=	16'h	222d;
2766	:douta	=	16'h	1969;
2767	:douta	=	16'h	63d2;
2768	:douta	=	16'h	8cb5;
2769	:douta	=	16'h	9d16;
2770	:douta	=	16'h	6bd2;
2771	:douta	=	16'h	4aee;
2772	:douta	=	16'h	c63a;
2773	:douta	=	16'h	84d7;
2774	:douta	=	16'h	6c16;
2775	:douta	=	16'h	19ac;
2776	:douta	=	16'h	29ec;
2777	:douta	=	16'h	328e;
2778	:douta	=	16'h	9516;
2779	:douta	=	16'h	9517;
2780	:douta	=	16'h	d69a;
2781	:douta	=	16'h	b5b9;
2782	:douta	=	16'h	84d7;
2783	:douta	=	16'h	6416;
2784	:douta	=	16'h	4b54;
2785	:douta	=	16'h	84d6;
2786	:douta	=	16'h	4394;
2787	:douta	=	16'h	5bb3;
2788	:douta	=	16'h	4bd5;
2789	:douta	=	16'h	5bd4;
2790	:douta	=	16'h	b65c;
2791	:douta	=	16'h	959a;
2792	:douta	=	16'h	7477;
2793	:douta	=	16'h	6437;
2794	:douta	=	16'h	21ac;
2795	:douta	=	16'h	2a6f;
2796	:douta	=	16'h	222d;
2797	:douta	=	16'h	7cd7;
2798	:douta	=	16'h	9518;
2799	:douta	=	16'h	9518;
2800	:douta	=	16'h	5b94;
2801	:douta	=	16'h	7c77;
2802	:douta	=	16'h	2a4f;
2803	:douta	=	16'h	42f0;
2804	:douta	=	16'h	42f0;
2805	:douta	=	16'h	63b3;
2806	:douta	=	16'h	9517;
2807	:douta	=	16'h	7499;
2808	:douta	=	16'h	74b8;
2809	:douta	=	16'h	5c17;
2810	:douta	=	16'h	4375;
2811	:douta	=	16'h	3313;
2812	:douta	=	16'h	1a0d;
2813	:douta	=	16'h	7cb6;
2814	:douta	=	16'h	9d78;
2815	:douta	=	16'h	74d9;
2816	:douta	=	16'h	19ee;
2817	:douta	=	16'h	4bb5;
2818	:douta	=	16'h	32d1;
2819	:douta	=	16'h	53f6;
2820	:douta	=	16'h	7498;
2821	:douta	=	16'h	5352;
2822	:douta	=	16'h	63f5;
2823	:douta	=	16'h	6436;
2824	:douta	=	16'h	74b8;
2825	:douta	=	16'h	42d0;
2826	:douta	=	16'h	5b50;
2827	:douta	=	16'h	7414;
2828	:douta	=	16'h	a537;
2829	:douta	=	16'h	84d7;
2830	:douta	=	16'h	c61a;
2831	:douta	=	16'h	adfb;
2832	:douta	=	16'h	7c13;
2833	:douta	=	16'h	7c75;
2834	:douta	=	16'h	63b2;
2835	:douta	=	16'h	8452;
2836	:douta	=	16'h	7c14;
2837	:douta	=	16'h	ad77;
2838	:douta	=	16'h	8c95;
2839	:douta	=	16'h	ce59;
2840	:douta	=	16'h	194a;
2841	:douta	=	16'h	7350;
2842	:douta	=	16'h	8cd5;
2843	:douta	=	16'h	5352;
2844	:douta	=	16'h	9cf5;
2845	:douta	=	16'h	b577;
2846	:douta	=	16'h	e6d9;
2847	:douta	=	16'h	ad56;
2848	:douta	=	16'h	ce18;
2849	:douta	=	16'h	9d37;
2850	:douta	=	16'h	b597;
2851	:douta	=	16'h	8474;
2852	:douta	=	16'h	5b30;
2853	:douta	=	16'h	a515;
2854	:douta	=	16'h	b5d8;
2855	:douta	=	16'h	b598;
2856	:douta	=	16'h	bdd7;
2857	:douta	=	16'h	ad98;
2858	:douta	=	16'h	d65a;
2859	:douta	=	16'h	7413;
2860	:douta	=	16'h	8c94;
2861	:douta	=	16'h	b576;
2862	:douta	=	16'h	3aaf;
2863	:douta	=	16'h	83f2;
2864	:douta	=	16'h	9d35;
2865	:douta	=	16'h	d678;
2866	:douta	=	16'h	c5f7;
2867	:douta	=	16'h	e6ba;
2868	:douta	=	16'h	f77b;
2869	:douta	=	16'h	bd76;
2870	:douta	=	16'h	7413;
2871	:douta	=	16'h	4aee;
2872	:douta	=	16'h	83f0;
2873	:douta	=	16'h	b5d6;
2874	:douta	=	16'h	b596;
2875	:douta	=	16'h	bd95;
2876	:douta	=	16'h	eed8;
2877	:douta	=	16'h	de98;
2878	:douta	=	16'h	9473;
2879	:douta	=	16'h	ad75;
2880	:douta	=	16'h	426d;
2881	:douta	=	16'h	7bf2;
2882	:douta	=	16'h	6bf2;
2883	:douta	=	16'h	6370;
2884	:douta	=	16'h	f79a;
2885	:douta	=	16'h	9cd5;
2886	:douta	=	16'h	de79;
2887	:douta	=	16'h	b5b7;
2888	:douta	=	16'h	e71b;
2889	:douta	=	16'h	4b94;
2890	:douta	=	16'h	be19;
2891	:douta	=	16'h	be18;
2892	:douta	=	16'h	8cb4;
2893	:douta	=	16'h	be17;
2894	:douta	=	16'h	ad77;
2895	:douta	=	16'h	bdf9;
2896	:douta	=	16'h	ef1b;
2897	:douta	=	16'h	8cd8;
2898	:douta	=	16'h	bdf9;
2899	:douta	=	16'h	1a0e;
2900	:douta	=	16'h	7c33;
2901	:douta	=	16'h	9d78;
2902	:douta	=	16'h	be18;
2903	:douta	=	16'h	a5b9;
2904	:douta	=	16'h	be5a;
2905	:douta	=	16'h	e71c;
2906	:douta	=	16'h	7476;
2907	:douta	=	16'h	95ba;
2908	:douta	=	16'h	3b33;
2909	:douta	=	16'h	94d7;
2910	:douta	=	16'h	63f3;
2911	:douta	=	16'h	4b51;
2912	:douta	=	16'h	8495;
2913	:douta	=	16'h	9557;
2914	:douta	=	16'h	8d38;
2915	:douta	=	16'h	ad97;
2916	:douta	=	16'h	be1a;
2917	:douta	=	16'h	7496;
2918	:douta	=	16'h	94d6;
2919	:douta	=	16'h	6c96;
2920	:douta	=	16'h	6b93;
2921	:douta	=	16'h	8d99;
2922	:douta	=	16'h	5b72;
2923	:douta	=	16'h	9d78;
2924	:douta	=	16'h	5bf5;
2925	:douta	=	16'h	7c75;
2926	:douta	=	16'h	9538;
2927	:douta	=	16'h	b619;
2928	:douta	=	16'h	d6ba;
2929	:douta	=	16'h	84d8;
2930	:douta	=	16'h	9d78;
2931	:douta	=	16'h	4b74;
2932	:douta	=	16'h	8c95;
2933	:douta	=	16'h	7434;
2934	:douta	=	16'h	8c94;
2935	:douta	=	16'h	9d36;
2936	:douta	=	16'h	9cd6;
2937	:douta	=	16'h	a4f4;
2938	:douta	=	16'h	b596;
2939	:douta	=	16'h	6bd1;
2940	:douta	=	16'h	5b10;
2941	:douta	=	16'h	530f;
2942	:douta	=	16'h	7c53;
2943	:douta	=	16'h	7c53;
2944	:douta	=	16'h	a535;
2945	:douta	=	16'h	8473;
2946	:douta	=	16'h	a576;
2947	:douta	=	16'h	b5b8;
2948	:douta	=	16'h	7c33;
2949	:douta	=	16'h	a576;
2950	:douta	=	16'h	42ef;
2951	:douta	=	16'h	530e;
2952	:douta	=	16'h	1106;
2953	:douta	=	16'h	422b;
2954	:douta	=	16'h	426b;
2955	:douta	=	16'h	424a;
2956	:douta	=	16'h	a536;
2957	:douta	=	16'h	2104;
2958	:douta	=	16'h	2103;
2959	:douta	=	16'h	18e3;
2960	:douta	=	16'h	10a2;
2961	:douta	=	16'h	31c8;
2962	:douta	=	16'h	29a9;
2963	:douta	=	16'h	29a8;
2964	:douta	=	16'h	73d0;
2965	:douta	=	16'h	5aed;
2966	:douta	=	16'h	6b6f;
2967	:douta	=	16'h	a4f4;
2968	:douta	=	16'h	634f;
2969	:douta	=	16'h	2967;
2970	:douta	=	16'h	632e;
2971	:douta	=	16'h	320b;
2972	:douta	=	16'h	5b0d;
2973	:douta	=	16'h	8c93;
2974	:douta	=	16'h	526a;
2975	:douta	=	16'h	bd33;
2976	:douta	=	16'h	73b0;
2977	:douta	=	16'h	7412;
2978	:douta	=	16'h	532f;
2979	:douta	=	16'h	7c31;
2980	:douta	=	16'h	4a8c;
2981	:douta	=	16'h	6b8f;
2982	:douta	=	16'h	a4f4;
2983	:douta	=	16'h	ce37;
2984	:douta	=	16'h	5b0e;
2985	:douta	=	16'h	7baf;
2986	:douta	=	16'h	4ace;
2987	:douta	=	16'h	3a2c;
2988	:douta	=	16'h	9d14;
2989	:douta	=	16'h	7bf1;
2990	:douta	=	16'h	9472;
2991	:douta	=	16'h	a536;
2992	:douta	=	16'h	8c52;
2993	:douta	=	16'h	42d0;
2994	:douta	=	16'h	4ace;
2995	:douta	=	16'h	5b70;
2996	:douta	=	16'h	8c72;
2997	:douta	=	16'h	c638;
2998	:douta	=	16'h	6bd2;
2999	:douta	=	16'h	bdd7;
3000	:douta	=	16'h	9cf4;
3001	:douta	=	16'h	a4d5;
3002	:douta	=	16'h	9cf5;
3003	:douta	=	16'h	1083;
3004	:douta	=	16'h	10e5;
3005	:douta	=	16'h	08c4;
3006	:douta	=	16'h	29a9;
3007	:douta	=	16'h	7413;
3008	:douta	=	16'h	532f;
3009	:douta	=	16'h	7413;
3010	:douta	=	16'h	9cd5;
3011	:douta	=	16'h	73f3;
3012	:douta	=	16'h	5b70;
3013	:douta	=	16'h	7bf1;
3014	:douta	=	16'h	5b50;
3015	:douta	=	16'h	5350;
3016	:douta	=	16'h	0065;
3017	:douta	=	16'h	2a0b;
3018	:douta	=	16'h	7c31;
3019	:douta	=	16'h	94d4;
3020	:douta	=	16'h	ad75;
3021	:douta	=	16'h	7413;
3022	:douta	=	16'h	94d4;
3023	:douta	=	16'h	328f;
3024	:douta	=	16'h	326d;
3025	:douta	=	16'h	00c8;
3026	:douta	=	16'h	6bf3;
3027	:douta	=	16'h	42ad;
3028	:douta	=	16'h	6b90;
3029	:douta	=	16'h	63b1;
3030	:douta	=	16'h	63d3;
3031	:douta	=	16'h	9517;
3032	:douta	=	16'h	b61a;
3033	:douta	=	16'h	adb9;
3034	:douta	=	16'h	3a8f;
3035	:douta	=	16'h	6392;
3036	:douta	=	16'h	53b4;
3037	:douta	=	16'h	3ad1;
3038	:douta	=	16'h	4b52;
3039	:douta	=	16'h	7436;
3040	:douta	=	16'h	84b6;
3041	:douta	=	16'h	84d8;
3042	:douta	=	16'h	6c36;
3043	:douta	=	16'h	7cda;
3044	:douta	=	16'h	8455;
3045	:douta	=	16'h	9559;
3046	:douta	=	16'h	00e9;
3047	:douta	=	16'h	2a2d;
3048	:douta	=	16'h	5415;
3049	:douta	=	16'h	5373;
3050	:douta	=	16'h	b61a;
3051	:douta	=	16'h	84f9;
3052	:douta	=	16'h	9539;
3053	:douta	=	16'h	116a;
3054	:douta	=	16'h	6c35;
3055	:douta	=	16'h	5b93;
3056	:douta	=	16'h	9d38;
3057	:douta	=	16'h	9558;
3058	:douta	=	16'h	5310;
3059	:douta	=	16'h	5b52;
3060	:douta	=	16'h	2a6f;
3061	:douta	=	16'h	6436;
3062	:douta	=	16'h	2ad2;
3063	:douta	=	16'h	118b;
3064	:douta	=	16'h	6415;
3065	:douta	=	16'h	8d19;
3066	:douta	=	16'h	6459;
3067	:douta	=	16'h	5bb5;
3068	:douta	=	16'h	853b;
3069	:douta	=	16'h	5c38;
3070	:douta	=	16'h	5c36;
3071	:douta	=	16'h	3b33;
3072	:douta	=	16'h	4b73;
3073	:douta	=	16'h	4b94;
3074	:douta	=	16'h	53f6;
3075	:douta	=	16'h	4bd5;
3076	:douta	=	16'h	32b0;
3077	:douta	=	16'h	3af0;
3078	:douta	=	16'h	5b93;
3079	:douta	=	16'h	6bf5;
3080	:douta	=	16'h	7497;
3081	:douta	=	16'h	7c76;
3082	:douta	=	16'h	42cf;
3083	:douta	=	16'h	5393;
3084	:douta	=	16'h	4b31;
3085	:douta	=	16'h	4b11;
3086	:douta	=	16'h	ad97;
3087	:douta	=	16'h	a599;
3088	:douta	=	16'h	c5d8;
3089	:douta	=	16'h	ce5b;
3090	:douta	=	16'h	9d16;
3091	:douta	=	16'h	8454;
3092	:douta	=	16'h	63b2;
3093	:douta	=	16'h	7c33;
3094	:douta	=	16'h	5b6f;
3095	:douta	=	16'h	be19;
3096	:douta	=	16'h	73f3;
3097	:douta	=	16'h	b597;
3098	:douta	=	16'h	b5d9;
3099	:douta	=	16'h	9d37;
3100	:douta	=	16'h	9cf6;
3101	:douta	=	16'h	8454;
3102	:douta	=	16'h	bdd7;
3103	:douta	=	16'h	be17;
3104	:douta	=	16'h	bdd8;
3105	:douta	=	16'h	be18;
3106	:douta	=	16'h	c638;
3107	:douta	=	16'h	ded9;
3108	:douta	=	16'h	9d16;
3109	:douta	=	16'h	e6fb;
3110	:douta	=	16'h	9d37;
3111	:douta	=	16'h	9495;
3112	:douta	=	16'h	7c53;
3113	:douta	=	16'h	ad56;
3114	:douta	=	16'h	b5b7;
3115	:douta	=	16'h	b597;
3116	:douta	=	16'h	e699;
3117	:douta	=	16'h	f73a;
3118	:douta	=	16'h	7c13;
3119	:douta	=	16'h	ad35;
3120	:douta	=	16'h	94d4;
3121	:douta	=	16'h	7433;
3122	:douta	=	16'h	7c52;
3123	:douta	=	16'h	ce38;
3124	:douta	=	16'h	ce78;
3125	:douta	=	16'h	deb8;
3126	:douta	=	16'h	a556;
3127	:douta	=	16'h	8474;
3128	:douta	=	16'h	b575;
3129	:douta	=	16'h	94d4;
3130	:douta	=	16'h	7c11;
3131	:douta	=	16'h	8432;
3132	:douta	=	16'h	c5f6;
3133	:douta	=	16'h	c637;
3134	:douta	=	16'h	ad33;
3135	:douta	=	16'h	e6d9;
3136	:douta	=	16'h	cdf7;
3137	:douta	=	16'h	e71a;
3138	:douta	=	16'h	6bd2;
3139	:douta	=	16'h	0908;
3140	:douta	=	16'h	ad75;
3141	:douta	=	16'h	2a2b;
3142	:douta	=	16'h	ce37;
3143	:douta	=	16'h	c5f9;
3144	:douta	=	16'h	eefa;
3145	:douta	=	16'h	53d5;
3146	:douta	=	16'h	bdb9;
3147	:douta	=	16'h	ce7a;
3148	:douta	=	16'h	5b71;
3149	:douta	=	16'h	9494;
3150	:douta	=	16'h	63b3;
3151	:douta	=	16'h	b5d8;
3152	:douta	=	16'h	d6ba;
3153	:douta	=	16'h	ce5b;
3154	:douta	=	16'h	ef3b;
3155	:douta	=	16'h	7c56;
3156	:douta	=	16'h	ce38;
3157	:douta	=	16'h	9d58;
3158	:douta	=	16'h	84b7;
3159	:douta	=	16'h	7476;
3160	:douta	=	16'h	9579;
3161	:douta	=	16'h	8d37;
3162	:douta	=	16'h	8454;
3163	:douta	=	16'h	959a;
3164	:douta	=	16'h	7cb8;
3165	:douta	=	16'h	b5b8;
3166	:douta	=	16'h	c67a;
3167	:douta	=	16'h	5395;
3168	:douta	=	16'h	4b10;
3169	:douta	=	16'h	4b73;
3170	:douta	=	16'h	5b52;
3171	:douta	=	16'h	5351;
3172	:douta	=	16'h	63d2;
3173	:douta	=	16'h	6bd4;
3174	:douta	=	16'h	c65a;
3175	:douta	=	16'h	a599;
3176	:douta	=	16'h	94b6;
3177	:douta	=	16'h	a65c;
3178	:douta	=	16'h	7c56;
3179	:douta	=	16'h	8496;
3180	:douta	=	16'h	6434;
3181	:douta	=	16'h	5bb3;
3182	:douta	=	16'h	3ad1;
3183	:douta	=	16'h	9517;
3184	:douta	=	16'h	b5f9;
3185	:douta	=	16'h	7c76;
3186	:douta	=	16'h	adb8;
3187	:douta	=	16'h	7456;
3188	:douta	=	16'h	deba;
3189	:douta	=	16'h	a5d9;
3190	:douta	=	16'h	4a8d;
3191	:douta	=	16'h	636f;
3192	:douta	=	16'h	42ae;
3193	:douta	=	16'h	d658;
3194	:douta	=	16'h	ad76;
3195	:douta	=	16'h	ad98;
3196	:douta	=	16'h	7c13;
3197	:douta	=	16'h	7c54;
3198	:douta	=	16'h	8413;
3199	:douta	=	16'h	4aef;
3200	:douta	=	16'h	52ce;
3201	:douta	=	16'h	218a;
3202	:douta	=	16'h	a598;
3203	:douta	=	16'h	8cb5;
3204	:douta	=	16'h	7c95;
3205	:douta	=	16'h	be39;
3206	:douta	=	16'h	7455;
3207	:douta	=	16'h	b575;
3208	:douta	=	16'h	2a4d;
3209	:douta	=	16'h	6b6f;
3210	:douta	=	16'h	3a4a;
3211	:douta	=	16'h	10e5;
3212	:douta	=	16'h	8472;
3213	:douta	=	16'h	3166;
3214	:douta	=	16'h	2924;
3215	:douta	=	16'h	1903;
3216	:douta	=	16'h	0020;
3217	:douta	=	16'h	83cf;
3218	:douta	=	16'h	4a6a;
3219	:douta	=	16'h	424a;
3220	:douta	=	16'h	29a9;
3221	:douta	=	16'h	29e9;
3222	:douta	=	16'h	4aad;
3223	:douta	=	16'h	ad75;
3224	:douta	=	16'h	8c94;
3225	:douta	=	16'h	8c31;
3226	:douta	=	16'h	a4f3;
3227	:douta	=	16'h	62cc;
3228	:douta	=	16'h	2188;
3229	:douta	=	16'h	31c9;
3230	:douta	=	16'h	7bf0;
3231	:douta	=	16'h	94d3;
3232	:douta	=	16'h	ad55;
3233	:douta	=	16'h	6bb1;
3234	:douta	=	16'h	42ae;
3235	:douta	=	16'h	3a2b;
3236	:douta	=	16'h	5acd;
3237	:douta	=	16'h	3a6c;
3238	:douta	=	16'h	42ee;
3239	:douta	=	16'h	8472;
3240	:douta	=	16'h	a514;
3241	:douta	=	16'h	c5f6;
3242	:douta	=	16'h	73d1;
3243	:douta	=	16'h	7bd0;
3244	:douta	=	16'h	4acf;
3245	:douta	=	16'h	52ad;
3246	:douta	=	16'h	8431;
3247	:douta	=	16'h	73b0;
3248	:douta	=	16'h	c5f6;
3249	:douta	=	16'h	63d2;
3250	:douta	=	16'h	7bf1;
3251	:douta	=	16'h	8433;
3252	:douta	=	16'h	5b2f;
3253	:douta	=	16'h	7432;
3254	:douta	=	16'h	6bd1;
3255	:douta	=	16'h	b596;
3256	:douta	=	16'h	8c94;
3257	:douta	=	16'h	ad77;
3258	:douta	=	16'h	bdd7;
3259	:douta	=	16'h	0883;
3260	:douta	=	16'h	08c4;
3261	:douta	=	16'h	10c3;
3262	:douta	=	16'h	1127;
3263	:douta	=	16'h	3a6c;
3264	:douta	=	16'h	5330;
3265	:douta	=	16'h	322c;
3266	:douta	=	16'h	4b0f;
3267	:douta	=	16'h	7c11;
3268	:douta	=	16'h	9492;
3269	:douta	=	16'h	8c93;
3270	:douta	=	16'h	7bf2;
3271	:douta	=	16'h	73f2;
3272	:douta	=	16'h	31ec;
3273	:douta	=	16'h	6b70;
3274	:douta	=	16'h	21aa;
3275	:douta	=	16'h	19ab;
3276	:douta	=	16'h	4b51;
3277	:douta	=	16'h	ad76;
3278	:douta	=	16'h	ce58;
3279	:douta	=	16'h	73d2;
3280	:douta	=	16'h	63d3;
3281	:douta	=	16'h	3aaf;
3282	:douta	=	16'h	63b1;
3283	:douta	=	16'h	322c;
3284	:douta	=	16'h	6390;
3285	:douta	=	16'h	2a4e;
3286	:douta	=	16'h	2a4e;
3287	:douta	=	16'h	9d78;
3288	:douta	=	16'h	84f7;
3289	:douta	=	16'h	b5f9;
3290	:douta	=	16'h	94f7;
3291	:douta	=	16'h	c67b;
3292	:douta	=	16'h	6436;
3293	:douta	=	16'h	63f4;
3294	:douta	=	16'h	32d1;
3295	:douta	=	16'h	63f5;
3296	:douta	=	16'h	2a8f;
3297	:douta	=	16'h	7476;
3298	:douta	=	16'h	7cf8;
3299	:douta	=	16'h	6c56;
3300	:douta	=	16'h	b61b;
3301	:douta	=	16'h	ae5d;
3302	:douta	=	16'h	5b93;
3303	:douta	=	16'h	63f4;
3304	:douta	=	16'h	2270;
3305	:douta	=	16'h	3ad0;
3306	:douta	=	16'h	4332;
3307	:douta	=	16'h	8d17;
3308	:douta	=	16'h	84d8;
3309	:douta	=	16'h	9518;
3310	:douta	=	16'h	7456;
3311	:douta	=	16'h	4b52;
3312	:douta	=	16'h	5bd3;
3313	:douta	=	16'h	4b73;
3314	:douta	=	16'h	73f3;
3315	:douta	=	16'h	8495;
3316	:douta	=	16'h	7bd2;
3317	:douta	=	16'h	7d1a;
3318	:douta	=	16'h	3b33;
3319	:douta	=	16'h	19cc;
3320	:douta	=	16'h	222e;
3321	:douta	=	16'h	4332;
3322	:douta	=	16'h	3b96;
3323	:douta	=	16'h	8cd6;
3324	:douta	=	16'h	74b7;
3325	:douta	=	16'h	8d3a;
3326	:douta	=	16'h	7d3b;
3327	:douta	=	16'h	6478;
3328	:douta	=	16'h	222f;
3329	:douta	=	16'h	6c77;
3330	:douta	=	16'h	6436;
3331	:douta	=	16'h	7d1a;
3332	:douta	=	16'h	53d4;
3333	:douta	=	16'h	42d0;
3334	:douta	=	16'h	42f1;
3335	:douta	=	16'h	5393;
3336	:douta	=	16'h	5394;
3337	:douta	=	16'h	3aaf;
3338	:douta	=	16'h	6b92;
3339	:douta	=	16'h	7434;
3340	:douta	=	16'h	9d38;
3341	:douta	=	16'h	9538;
3342	:douta	=	16'h	8453;
3343	:douta	=	16'h	9d37;
3344	:douta	=	16'h	5b92;
3345	:douta	=	16'h	6bd2;
3346	:douta	=	16'h	6c14;
3347	:douta	=	16'h	8453;
3348	:douta	=	16'h	a536;
3349	:douta	=	16'h	e6fb;
3350	:douta	=	16'h	a5b9;
3351	:douta	=	16'h	8c94;
3352	:douta	=	16'h	a578;
3353	:douta	=	16'h	5352;
3354	:douta	=	16'h	7c13;
3355	:douta	=	16'h	324e;
3356	:douta	=	16'h	c618;
3357	:douta	=	16'h	a536;
3358	:douta	=	16'h	c5d7;
3359	:douta	=	16'h	9d15;
3360	:douta	=	16'h	94d4;
3361	:douta	=	16'h	9cf6;
3362	:douta	=	16'h	7413;
3363	:douta	=	16'h	7413;
3364	:douta	=	16'h	8432;
3365	:douta	=	16'h	a555;
3366	:douta	=	16'h	bdf8;
3367	:douta	=	16'h	de98;
3368	:douta	=	16'h	d6fb;
3369	:douta	=	16'h	ce38;
3370	:douta	=	16'h	b619;
3371	:douta	=	16'h	9493;
3372	:douta	=	16'h	8c73;
3373	:douta	=	16'h	a576;
3374	:douta	=	16'h	8cb3;
3375	:douta	=	16'h	bdd7;
3376	:douta	=	16'h	ef3a;
3377	:douta	=	16'h	de98;
3378	:douta	=	16'h	ce7a;
3379	:douta	=	16'h	bd96;
3380	:douta	=	16'h	deba;
3381	:douta	=	16'h	83f1;
3382	:douta	=	16'h	63d1;
3383	:douta	=	16'h	5aee;
3384	:douta	=	16'h	ce56;
3385	:douta	=	16'h	c616;
3386	:douta	=	16'h	ff5a;
3387	:douta	=	16'h	8c93;
3388	:douta	=	16'h	acd4;
3389	:douta	=	16'h	9d35;
3390	:douta	=	16'h	530f;
3391	:douta	=	16'h	8c93;
3392	:douta	=	16'h	73b1;
3393	:douta	=	16'h	c5f7;
3394	:douta	=	16'h	9d36;
3395	:douta	=	16'h	9d15;
3396	:douta	=	16'h	e6f9;
3397	:douta	=	16'h	94f6;
3398	:douta	=	16'h	6372;
3399	:douta	=	16'h	8cb4;
3400	:douta	=	16'h	4b0e;
3401	:douta	=	16'h	a577;
3402	:douta	=	16'h	d6ba;
3403	:douta	=	16'h	deba;
3404	:douta	=	16'h	bdf9;
3405	:douta	=	16'h	e6fb;
3406	:douta	=	16'h	8496;
3407	:douta	=	16'h	e71c;
3408	:douta	=	16'h	7cf8;
3409	:douta	=	16'h	39c9;
3410	:douta	=	16'h	94d4;
3411	:douta	=	16'h	8cf7;
3412	:douta	=	16'h	ce79;
3413	:douta	=	16'h	adf9;
3414	:douta	=	16'h	f75b;
3415	:douta	=	16'h	8538;
3416	:douta	=	16'h	ce5a;
3417	:douta	=	16'h	ceba;
3418	:douta	=	16'h	a578;
3419	:douta	=	16'h	3af0;
3420	:douta	=	16'h	5bd3;
3421	:douta	=	16'h	73f2;
3422	:douta	=	16'h	b5d8;
3423	:douta	=	16'h	8c94;
3424	:douta	=	16'h	6415;
3425	:douta	=	16'h	b5b9;
3426	:douta	=	16'h	df1b;
3427	:douta	=	16'h	b69c;
3428	:douta	=	16'h	8454;
3429	:douta	=	16'h	42f1;
3430	:douta	=	16'h	6bd3;
3431	:douta	=	16'h	3af0;
3432	:douta	=	16'h	220c;
3433	:douta	=	16'h	5373;
3434	:douta	=	16'h	c65b;
3435	:douta	=	16'h	a5b8;
3436	:douta	=	16'h	6c76;
3437	:douta	=	16'h	a578;
3438	:douta	=	16'h	4354;
3439	:douta	=	16'h	d69b;
3440	:douta	=	16'h	8559;
3441	:douta	=	16'h	7c75;
3442	:douta	=	16'h	7c97;
3443	:douta	=	16'h	63f4;
3444	:douta	=	16'h	5bb2;
3445	:douta	=	16'h	3a2c;
3446	:douta	=	16'h	9d14;
3447	:douta	=	16'h	6c12;
3448	:douta	=	16'h	ad77;
3449	:douta	=	16'h	adb7;
3450	:douta	=	16'h	9494;
3451	:douta	=	16'h	5350;
3452	:douta	=	16'h	4ace;
3453	:douta	=	16'h	5b2f;
3454	:douta	=	16'h	9557;
3455	:douta	=	16'h	7c53;
3456	:douta	=	16'h	be19;
3457	:douta	=	16'h	8c74;
3458	:douta	=	16'h	8c72;
3459	:douta	=	16'h	324b;
3460	:douta	=	16'h	2947;
3461	:douta	=	16'h	430e;
3462	:douta	=	16'h	84d6;
3463	:douta	=	16'h	4aef;
3464	:douta	=	16'h	94b3;
3465	:douta	=	16'h	de98;
3466	:douta	=	16'h	a536;
3467	:douta	=	16'h	8c32;
3468	:douta	=	16'h	83f1;
3469	:douta	=	16'h	528a;
3470	:douta	=	16'h	2925;
3471	:douta	=	16'h	2104;
3472	:douta	=	16'h	18c3;
3473	:douta	=	16'h	5b0c;
3474	:douta	=	16'h	b594;
3475	:douta	=	16'h	73d0;
3476	:douta	=	16'h	ad34;
3477	:douta	=	16'h	c637;
3478	:douta	=	16'h	83f0;
3479	:douta	=	16'h	29ca;
3480	:douta	=	16'h	0085;
3481	:douta	=	16'h	5b2d;
3482	:douta	=	16'h	6bb0;
3483	:douta	=	16'h	73d1;
3484	:douta	=	16'h	73b0;
3485	:douta	=	16'h	9c92;
3486	:douta	=	16'h	73d0;
3487	:douta	=	16'h	31ea;
3488	:douta	=	16'h	52ed;
3489	:douta	=	16'h	52ed;
3490	:douta	=	16'h	7c31;
3491	:douta	=	16'h	5b4e;
3492	:douta	=	16'h	7c51;
3493	:douta	=	16'h	73d1;
3494	:douta	=	16'h	7c32;
3495	:douta	=	16'h	8c11;
3496	:douta	=	16'h	8cb5;
3497	:douta	=	16'h	0928;
3498	:douta	=	16'h	8473;
3499	:douta	=	16'h	6bd2;
3500	:douta	=	16'h	9493;
3501	:douta	=	16'h	be77;
3502	:douta	=	16'h	8cd4;
3503	:douta	=	16'h	8cb3;
3504	:douta	=	16'h	4b50;
3505	:douta	=	16'h	4aac;
3506	:douta	=	16'h	4b0e;
3507	:douta	=	16'h	428c;
3508	:douta	=	16'h	536e;
3509	:douta	=	16'h	328c;
3510	:douta	=	16'h	29c9;
3511	:douta	=	16'h	08e6;
3512	:douta	=	16'h	1988;
3513	:douta	=	16'h	08e6;
3514	:douta	=	16'h	1127;
3515	:douta	=	16'h	10a3;
3516	:douta	=	16'h	08a4;
3517	:douta	=	16'h	10a3;
3518	:douta	=	16'h	29e9;
3519	:douta	=	16'h	8cf4;
3520	:douta	=	16'h	4acf;
3521	:douta	=	16'h	84d5;
3522	:douta	=	16'h	5bb4;
3523	:douta	=	16'h	63b1;
3524	:douta	=	16'h	5b70;
3525	:douta	=	16'h	8493;
3526	:douta	=	16'h	73f2;
3527	:douta	=	16'h	5b70;
3528	:douta	=	16'h	bdb5;
3529	:douta	=	16'h	9cb2;
3530	:douta	=	16'h	6350;
3531	:douta	=	16'h	2a4d;
3532	:douta	=	16'h	00c6;
3533	:douta	=	16'h	4aef;
3534	:douta	=	16'h	0949;
3535	:douta	=	16'h	7474;
3536	:douta	=	16'h	6c35;
3537	:douta	=	16'h	7434;
3538	:douta	=	16'h	c5f8;
3539	:douta	=	16'h	8474;
3540	:douta	=	16'h	9d36;
3541	:douta	=	16'h	29ec;
3542	:douta	=	16'h	326e;
3543	:douta	=	16'h	29ed;
3544	:douta	=	16'h	21cd;
3545	:douta	=	16'h	5bd5;
3546	:douta	=	16'h	5351;
3547	:douta	=	16'h	5bd4;
3548	:douta	=	16'h	9517;
3549	:douta	=	16'h	9d78;
3550	:douta	=	16'h	6c56;
3551	:douta	=	16'h	a5da;
3552	:douta	=	16'h	8d59;
3553	:douta	=	16'h	6c35;
3554	:douta	=	16'h	4b53;
3555	:douta	=	16'h	4b31;
3556	:douta	=	16'h	2ab0;
3557	:douta	=	16'h	5373;
3558	:douta	=	16'h	7cd7;
3559	:douta	=	16'h	8519;
3560	:douta	=	16'h	8cb6;
3561	:douta	=	16'h	53b5;
3562	:douta	=	16'h	84b7;
3563	:douta	=	16'h	118c;
3564	:douta	=	16'h	2a2d;
3565	:douta	=	16'h	7455;
3566	:douta	=	16'h	84f8;
3567	:douta	=	16'h	84d7;
3568	:douta	=	16'h	4b73;
3569	:douta	=	16'h	3aaf;
3570	:douta	=	16'h	5bb4;
3571	:douta	=	16'h	5bd3;
3572	:douta	=	16'h	4372;
3573	:douta	=	16'h	6414;
3574	:douta	=	16'h	9d79;
3575	:douta	=	16'h	4353;
3576	:douta	=	16'h	7cd9;
3577	:douta	=	16'h	4bf7;
3578	:douta	=	16'h	4312;
3579	:douta	=	16'h	4373;
3580	:douta	=	16'h	1a50;
3581	:douta	=	16'h	8d5b;
3582	:douta	=	16'h	6458;
3583	:douta	=	16'h	9ddc;
3584	:douta	=	16'h	2a90;
3585	:douta	=	16'h	4b94;
3586	:douta	=	16'h	5c16;
3587	:douta	=	16'h	4332;
3588	:douta	=	16'h	3ad1;
3589	:douta	=	16'h	4b11;
3590	:douta	=	16'h	6c36;
3591	:douta	=	16'h	6c36;
3592	:douta	=	16'h	74b9;
3593	:douta	=	16'h	5352;
3594	:douta	=	16'h	63b3;
3595	:douta	=	16'h	116a;
3596	:douta	=	16'h	5b30;
3597	:douta	=	16'h	5bb3;
3598	:douta	=	16'h	b577;
3599	:douta	=	16'h	ce7b;
3600	:douta	=	16'h	9d37;
3601	:douta	=	16'h	c63a;
3602	:douta	=	16'h	7414;
3603	:douta	=	16'h	29eb;
3604	:douta	=	16'h	428d;
3605	:douta	=	16'h	9d16;
3606	:douta	=	16'h	9d17;
3607	:douta	=	16'h	ce79;
3608	:douta	=	16'h	ad97;
3609	:douta	=	16'h	9d17;
3610	:douta	=	16'h	b5d8;
3611	:douta	=	16'h	7414;
3612	:douta	=	16'h	a516;
3613	:douta	=	16'h	428e;
3614	:douta	=	16'h	73f1;
3615	:douta	=	16'h	bdd7;
3616	:douta	=	16'h	bdb6;
3617	:douta	=	16'h	bdd7;
3618	:douta	=	16'h	a536;
3619	:douta	=	16'h	bdf7;
3620	:douta	=	16'h	9493;
3621	:douta	=	16'h	b597;
3622	:douta	=	16'h	8cf6;
3623	:douta	=	16'h	bd95;
3624	:douta	=	16'h	c639;
3625	:douta	=	16'h	bdd7;
3626	:douta	=	16'h	ce59;
3627	:douta	=	16'h	ce38;
3628	:douta	=	16'h	acf5;
3629	:douta	=	16'h	e6b9;
3630	:douta	=	16'h	6bf1;
3631	:douta	=	16'h	de99;
3632	:douta	=	16'h	9cd5;
3633	:douta	=	16'h	a4f3;
3634	:douta	=	16'h	8cd4;
3635	:douta	=	16'h	ffbc;
3636	:douta	=	16'h	ef5b;
3637	:douta	=	16'h	c5d6;
3638	:douta	=	16'h	63b1;
3639	:douta	=	16'h	9c73;
3640	:douta	=	16'h	9492;
3641	:douta	=	16'h	b5b6;
3642	:douta	=	16'h	7bef;
3643	:douta	=	16'h	9cb3;
3644	:douta	=	16'h	de77;
3645	:douta	=	16'h	c657;
3646	:douta	=	16'h	a4f3;
3647	:douta	=	16'h	7c12;
3648	:douta	=	16'h	9452;
3649	:douta	=	16'h	a556;
3650	:douta	=	16'h	5b91;
3651	:douta	=	16'h	5b2f;
3652	:douta	=	16'h	ce78;
3653	:douta	=	16'h	9d15;
3654	:douta	=	16'h	ce18;
3655	:douta	=	16'h	a5b8;
3656	:douta	=	16'h	9473;
3657	:douta	=	16'h	5bb3;
3658	:douta	=	16'h	7433;
3659	:douta	=	16'h	a577;
3660	:douta	=	16'h	8c52;
3661	:douta	=	16'h	adf7;
3662	:douta	=	16'h	d659;
3663	:douta	=	16'h	e75c;
3664	:douta	=	16'h	ae1b;
3665	:douta	=	16'h	c5f9;
3666	:douta	=	16'h	a599;
3667	:douta	=	16'h	6414;
3668	:douta	=	16'h	84b5;
3669	:douta	=	16'h	4331;
3670	:douta	=	16'h	d6da;
3671	:douta	=	16'h	be5b;
3672	:douta	=	16'h	e6fb;
3673	:douta	=	16'h	be9a;
3674	:douta	=	16'h	be1a;
3675	:douta	=	16'h	6435;
3676	:douta	=	16'h	5bb4;
3677	:douta	=	16'h	322e;
3678	:douta	=	16'h	8473;
3679	:douta	=	16'h	3ab0;
3680	:douta	=	16'h	2a0e;
3681	:douta	=	16'h	7c76;
3682	:douta	=	16'h	a5b8;
3683	:douta	=	16'h	84f8;
3684	:douta	=	16'h	deba;
3685	:douta	=	16'h	7c97;
3686	:douta	=	16'h	b5d9;
3687	:douta	=	16'h	5bf5;
3688	:douta	=	16'h	5374;
3689	:douta	=	16'h	5bb4;
3690	:douta	=	16'h	9d98;
3691	:douta	=	16'h	5bb4;
3692	:douta	=	16'h	4b10;
3693	:douta	=	16'h	8cf7;
3694	:douta	=	16'h	8497;
3695	:douta	=	16'h	c639;
3696	:douta	=	16'h	8d39;
3697	:douta	=	16'h	ad98;
3698	:douta	=	16'h	8d18;
3699	:douta	=	16'h	42cf;
3700	:douta	=	16'h	7454;
3701	:douta	=	16'h	21aa;
3702	:douta	=	16'h	422a;
3703	:douta	=	16'h	4aad;
3704	:douta	=	16'h	8454;
3705	:douta	=	16'h	be3a;
3706	:douta	=	16'h	b5b8;
3707	:douta	=	16'h	5371;
3708	:douta	=	16'h	6330;
3709	:douta	=	16'h	2188;
3710	:douta	=	16'h	8495;
3711	:douta	=	16'h	52ee;
3712	:douta	=	16'h	8452;
3713	:douta	=	16'h	9cd5;
3714	:douta	=	16'h	bdf8;
3715	:douta	=	16'h	8c73;
3716	:douta	=	16'h	b575;
3717	:douta	=	16'h	19ed;
3718	:douta	=	16'h	322d;
3719	:douta	=	16'h	3a2b;
3720	:douta	=	16'h	3a4c;
3721	:douta	=	16'h	94f4;
3722	:douta	=	16'h	8cb5;
3723	:douta	=	16'h	9d15;
3724	:douta	=	16'h	8452;
3725	:douta	=	16'h	8c52;
3726	:douta	=	16'h	2925;
3727	:douta	=	16'h	2124;
3728	:douta	=	16'h	2104;
3729	:douta	=	16'h	39a6;
3730	:douta	=	16'h	6b8f;
3731	:douta	=	16'h	424a;
3732	:douta	=	16'h	5acc;
3733	:douta	=	16'h	7410;
3734	:douta	=	16'h	de37;
3735	:douta	=	16'h	7370;
3736	:douta	=	16'h	52cd;
3737	:douta	=	16'h	4aad;
3738	:douta	=	16'h	39ca;
3739	:douta	=	16'h	1948;
3740	:douta	=	16'h	73f0;
3741	:douta	=	16'h	7c10;
3742	:douta	=	16'h	94b3;
3743	:douta	=	16'h	8c11;
3744	:douta	=	16'h	6b70;
3745	:douta	=	16'h	4aad;
3746	:douta	=	16'h	31a9;
3747	:douta	=	16'h	31cb;
3748	:douta	=	16'h	00c6;
3749	:douta	=	16'h	5b4f;
3750	:douta	=	16'h	73f1;
3751	:douta	=	16'h	c617;
3752	:douta	=	16'h	6c13;
3753	:douta	=	16'h	8432;
3754	:douta	=	16'h	7453;
3755	:douta	=	16'h	32ae;
3756	:douta	=	16'h	5b90;
3757	:douta	=	16'h	19c9;
3758	:douta	=	16'h	19a8;
3759	:douta	=	16'h	1147;
3760	:douta	=	16'h	0084;
3761	:douta	=	16'h	08e5;
3762	:douta	=	16'h	0002;
3763	:douta	=	16'h	0002;
3764	:douta	=	16'h	0022;
3765	:douta	=	16'h	0001;
3766	:douta	=	16'h	0042;
3767	:douta	=	16'h	0042;
3768	:douta	=	16'h	0022;
3769	:douta	=	16'h	0042;
3770	:douta	=	16'h	0001;
3771	:douta	=	16'h	0063;
3772	:douta	=	16'h	0062;
3773	:douta	=	16'h	0063;
3774	:douta	=	16'h	0022;
3775	:douta	=	16'h	0002;
3776	:douta	=	16'h	0043;
3777	:douta	=	16'h	21a8;
3778	:douta	=	16'h	2188;
3779	:douta	=	16'h	08e6;
3780	:douta	=	16'h	322b;
3781	:douta	=	16'h	2a2b;
3782	:douta	=	16'h	5371;
3783	:douta	=	16'h	7434;
3784	:douta	=	16'h	c637;
3785	:douta	=	16'h	bdd7;
3786	:douta	=	16'h	c596;
3787	:douta	=	16'h	5b30;
3788	:douta	=	16'h	426d;
3789	:douta	=	16'h	8474;
3790	:douta	=	16'h	19cb;
3791	:douta	=	16'h	19cd;
3792	:douta	=	16'h	6c34;
3793	:douta	=	16'h	42f0;
3794	:douta	=	16'h	ad97;
3795	:douta	=	16'h	9d36;
3796	:douta	=	16'h	8494;
3797	:douta	=	16'h	ad77;
3798	:douta	=	16'h	a557;
3799	:douta	=	16'h	63f4;
3800	:douta	=	16'h	7435;
3801	:douta	=	16'h	0129;
3802	:douta	=	16'h	3ab0;
3803	:douta	=	16'h	11ac;
3804	:douta	=	16'h	32b0;
3805	:douta	=	16'h	5bf5;
3806	:douta	=	16'h	4bb4;
3807	:douta	=	16'h	9d9a;
3808	:douta	=	16'h	8cd7;
3809	:douta	=	16'h	7cd8;
3810	:douta	=	16'h	3af1;
3811	:douta	=	16'h	7455;
3812	:douta	=	16'h	3b32;
3813	:douta	=	16'h	4b53;
3814	:douta	=	16'h	6414;
3815	:douta	=	16'h	63f5;
3816	:douta	=	16'h	b5d8;
3817	:douta	=	16'h	9d37;
3818	:douta	=	16'h	8cf6;
3819	:douta	=	16'h	3ad1;
3820	:douta	=	16'h	6c35;
3821	:douta	=	16'h	3af1;
3822	:douta	=	16'h	3a90;
3823	:douta	=	16'h	7456;
3824	:douta	=	16'h	7c55;
3825	:douta	=	16'h	ad77;
3826	:douta	=	16'h	5b93;
3827	:douta	=	16'h	53b4;
3828	:douta	=	16'h	1a2e;
3829	:douta	=	16'h	4311;
3830	:douta	=	16'h	4b53;
3831	:douta	=	16'h	7c76;
3832	:douta	=	16'h	7498;
3833	:douta	=	16'h	53f6;
3834	:douta	=	16'h	6c57;
3835	:douta	=	16'h	53f6;
3836	:douta	=	16'h	4bf7;
3837	:douta	=	16'h	5c58;
3838	:douta	=	16'h	3b53;
3839	:douta	=	16'h	6cb8;
3840	:douta	=	16'h	32b0;
3841	:douta	=	16'h	5b93;
3842	:douta	=	16'h	6c77;
3843	:douta	=	16'h	6498;
3844	:douta	=	16'h	6478;
3845	:douta	=	16'h	5bf5;
3846	:douta	=	16'h	2a6e;
3847	:douta	=	16'h	4352;
3848	:douta	=	16'h	4311;
3849	:douta	=	16'h	63d3;
3850	:douta	=	16'h	94f6;
3851	:douta	=	16'h	8518;
3852	:douta	=	16'h	9d58;
3853	:douta	=	16'h	4b31;
3854	:douta	=	16'h	42ef;
3855	:douta	=	16'h	426e;
3856	:douta	=	16'h	42ef;
3857	:douta	=	16'h	6392;
3858	:douta	=	16'h	bdd8;
3859	:douta	=	16'h	c5d7;
3860	:douta	=	16'h	ce5a;
3861	:douta	=	16'h	ad55;
3862	:douta	=	16'h	7c54;
3863	:douta	=	16'h	8cb4;
3864	:douta	=	16'h	8c74;
3865	:douta	=	16'h	5352;
3866	:douta	=	16'h	7bf3;
3867	:douta	=	16'h	6bd2;
3868	:douta	=	16'h	94b5;
3869	:douta	=	16'h	be39;
3870	:douta	=	16'h	ad37;
3871	:douta	=	16'h	be38;
3872	:douta	=	16'h	ad57;
3873	:douta	=	16'h	8c95;
3874	:douta	=	16'h	7454;
3875	:douta	=	16'h	5b30;
3876	:douta	=	16'h	9cf5;
3877	:douta	=	16'h	bdf7;
3878	:douta	=	16'h	adb8;
3879	:douta	=	16'h	f75a;
3880	:douta	=	16'h	e6db;
3881	:douta	=	16'h	84b5;
3882	:douta	=	16'h	9d15;
3883	:douta	=	16'h	9493;
3884	:douta	=	16'h	c617;
3885	:douta	=	16'h	ce78;
3886	:douta	=	16'h	bd75;
3887	:douta	=	16'h	deb9;
3888	:douta	=	16'h	ce59;
3889	:douta	=	16'h	e6dc;
3890	:douta	=	16'h	7476;
3891	:douta	=	16'h	8c11;
3892	:douta	=	16'h	94d2;
3893	:douta	=	16'h	4acd;
3894	:douta	=	16'h	a534;
3895	:douta	=	16'h	8c30;
3896	:douta	=	16'h	ff7b;
3897	:douta	=	16'h	bd95;
3898	:douta	=	16'h	f75b;
3899	:douta	=	16'h	83f2;
3900	:douta	=	16'h	94b3;
3901	:douta	=	16'h	9d15;
3902	:douta	=	16'h	8c92;
3903	:douta	=	16'h	8451;
3904	:douta	=	16'h	b596;
3905	:douta	=	16'h	f75a;
3906	:douta	=	16'h	b576;
3907	:douta	=	16'h	d657;
3908	:douta	=	16'h	8493;
3909	:douta	=	16'h	4a8e;
3910	:douta	=	16'h	73b0;
3911	:douta	=	16'h	4350;
3912	:douta	=	16'h	84b5;
3913	:douta	=	16'h	ad77;
3914	:douta	=	16'h	ff9c;
3915	:douta	=	16'h	9d98;
3916	:douta	=	16'h	bd75;
3917	:douta	=	16'h	c619;
3918	:douta	=	16'h	328f;
3919	:douta	=	16'h	9517;
3920	:douta	=	16'h	6c76;
3921	:douta	=	16'h	8432;
3922	:douta	=	16'h	a5d9;
3923	:douta	=	16'h	d67a;
3924	:douta	=	16'h	9578;
3925	:douta	=	16'h	9cd6;
3926	:douta	=	16'h	6cd9;
3927	:douta	=	16'h	32f3;
3928	:douta	=	16'h	ce9a;
3929	:douta	=	16'h	be5a;
3930	:douta	=	16'h	9537;
3931	:douta	=	16'h	84d7;
3932	:douta	=	16'h	84b6;
3933	:douta	=	16'h	ad98;
3934	:douta	=	16'h	d6dc;
3935	:douta	=	16'h	ce7b;
3936	:douta	=	16'h	5373;
3937	:douta	=	16'h	8475;
3938	:douta	=	16'h	b5f9;
3939	:douta	=	16'h	6c77;
3940	:douta	=	16'h	5b72;
3941	:douta	=	16'h	4b32;
3942	:douta	=	16'h	8cb5;
3943	:douta	=	16'h	8495;
3944	:douta	=	16'h	defa;
3945	:douta	=	16'h	6c98;
3946	:douta	=	16'h	d679;
3947	:douta	=	16'h	be9c;
3948	:douta	=	16'h	8d39;
3949	:douta	=	16'h	7497;
3950	:douta	=	16'h	a557;
3951	:douta	=	16'h	be5b;
3952	:douta	=	16'h	a5da;
3953	:douta	=	16'h	326f;
3954	:douta	=	16'h	5373;
3955	:douta	=	16'h	c639;
3956	:douta	=	16'h	7455;
3957	:douta	=	16'h	8c52;
3958	:douta	=	16'h	b5d7;
3959	:douta	=	16'h	6bd2;
3960	:douta	=	16'h	ad34;
3961	:douta	=	16'h	4aef;
3962	:douta	=	16'h	42ae;
3963	:douta	=	16'h	6391;
3964	:douta	=	16'h	8d17;
3965	:douta	=	16'h	deda;
3966	:douta	=	16'h	5b30;
3967	:douta	=	16'h	d5f8;
3968	:douta	=	16'h	4aae;
3969	:douta	=	16'h	52ce;
3970	:douta	=	16'h	630e;
3971	:douta	=	16'h	8473;
3972	:douta	=	16'h	b619;
3973	:douta	=	16'h	9d15;
3974	:douta	=	16'h	d658;
3975	:douta	=	16'h	5b70;
3976	:douta	=	16'h	9c72;
3977	:douta	=	16'h	8c93;
3978	:douta	=	16'h	2167;
3979	:douta	=	16'h	1926;
3980	:douta	=	16'h	1926;
3981	:douta	=	16'h	a576;
3982	:douta	=	16'h	5acb;
3983	:douta	=	16'h	2124;
3984	:douta	=	16'h	20e4;
3985	:douta	=	16'h	1082;
3986	:douta	=	16'h	ad75;
3987	:douta	=	16'h	5b0e;
3988	:douta	=	16'h	b554;
3989	:douta	=	16'h	4aac;
3990	:douta	=	16'h	5b0e;
3991	:douta	=	16'h	634e;
3992	:douta	=	16'h	5b4e;
3993	:douta	=	16'h	8451;
3994	:douta	=	16'h	a534;
3995	:douta	=	16'h	9492;
3996	:douta	=	16'h	9430;
3997	:douta	=	16'h	b533;
3998	:douta	=	16'h	634f;
3999	:douta	=	16'h	8cb3;
4000	:douta	=	16'h	4aad;
4001	:douta	=	16'h	6b6f;
4002	:douta	=	16'h	b5f6;
4003	:douta	=	16'h	6370;
4004	:douta	=	16'h	73f2;
4005	:douta	=	16'h	1148;
4006	:douta	=	16'h	428c;
4007	:douta	=	16'h	1127;
4008	:douta	=	16'h	0083;
4009	:douta	=	16'h	0022;
4010	:douta	=	16'h	0842;
4011	:douta	=	16'h	0863;
4012	:douta	=	16'h	0063;
4013	:douta	=	16'h	0884;
4014	:douta	=	16'h	08a4;
4015	:douta	=	16'h	08a4;
4016	:douta	=	16'h	08a4;
4017	:douta	=	16'h	08a4;
4018	:douta	=	16'h	0884;
4019	:douta	=	16'h	10c4;
4020	:douta	=	16'h	08a4;
4021	:douta	=	16'h	08a4;
4022	:douta	=	16'h	08c4;
4023	:douta	=	16'h	0884;
4024	:douta	=	16'h	0884;
4025	:douta	=	16'h	0884;
4026	:douta	=	16'h	08a4;
4027	:douta	=	16'h	0883;
4028	:douta	=	16'h	0883;
4029	:douta	=	16'h	0883;
4030	:douta	=	16'h	0063;
4031	:douta	=	16'h	0863;
4032	:douta	=	16'h	0863;
4033	:douta	=	16'h	0883;
4034	:douta	=	16'h	0883;
4035	:douta	=	16'h	0062;
4036	:douta	=	16'h	0062;
4037	:douta	=	16'h	0062;
4038	:douta	=	16'h	0021;
4039	:douta	=	16'h	0001;
4040	:douta	=	16'h	0022;
4041	:douta	=	16'h	0022;
4042	:douta	=	16'h	1167;
4043	:douta	=	16'h	42ad;
4044	:douta	=	16'h	9d34;
4045	:douta	=	16'h	9517;
4046	:douta	=	16'h	c63a;
4047	:douta	=	16'h	6436;
4048	:douta	=	16'h	6371;
4049	:douta	=	16'h	5bb3;
4050	:douta	=	16'h	322d;
4051	:douta	=	16'h	2a2d;
4052	:douta	=	16'h	9d36;
4053	:douta	=	16'h	5b51;
4054	:douta	=	16'h	7c74;
4055	:douta	=	16'h	d67a;
4056	:douta	=	16'h	7c55;
4057	:douta	=	16'h	84b6;
4058	:douta	=	16'h	7498;
4059	:douta	=	16'h	3af2;
4060	:douta	=	16'h	2a4f;
4061	:douta	=	16'h	222e;
4062	:douta	=	16'h	32af;
4063	:douta	=	16'h	222e;
4064	:douta	=	16'h	4b53;
4065	:douta	=	16'h	4b53;
4066	:douta	=	16'h	63f4;
4067	:douta	=	16'h	7476;
4068	:douta	=	16'h	b5ba;
4069	:douta	=	16'h	7c55;
4070	:douta	=	16'h	5351;
4071	:douta	=	16'h	5351;
4072	:douta	=	16'h	326e;
4073	:douta	=	16'h	3af1;
4074	:douta	=	16'h	5352;
4075	:douta	=	16'h	9517;
4076	:douta	=	16'h	a578;
4077	:douta	=	16'h	6415;
4078	:douta	=	16'h	7498;
4079	:douta	=	16'h	32f1;
4080	:douta	=	16'h	4b31;
4081	:douta	=	16'h	11ac;
4082	:douta	=	16'h	8cd6;
4083	:douta	=	16'h	6416;
4084	:douta	=	16'h	6c14;
4085	:douta	=	16'h	6457;
4086	:douta	=	16'h	5bf6;
4087	:douta	=	16'h	3b13;
4088	:douta	=	16'h	3b32;
4089	:douta	=	16'h	5bf6;
4090	:douta	=	16'h	8518;
4091	:douta	=	16'h	959c;
4092	:douta	=	16'h	5c38;
4093	:douta	=	16'h	6c78;
4094	:douta	=	16'h	74da;
4095	:douta	=	16'h	2ad2;
4096	:douta	=	16'h	1a0d;
4097	:douta	=	16'h	5332;
4098	:douta	=	16'h	7478;
4099	:douta	=	16'h	53f5;
4100	:douta	=	16'h	74d9;
4101	:douta	=	16'h	6498;
4102	:douta	=	16'h	5b93;
4103	:douta	=	16'h	328f;
4104	:douta	=	16'h	6c56;
4105	:douta	=	16'h	3aaf;
4106	:douta	=	16'h	6bb2;
4107	:douta	=	16'h	7c34;
4108	:douta	=	16'h	8c94;
4109	:douta	=	16'h	6bf4;
4110	:douta	=	16'h	94d5;
4111	:douta	=	16'h	a557;
4112	:douta	=	16'h	5bd3;
4113	:douta	=	16'h	42f0;
4114	:douta	=	16'h	5351;
4115	:douta	=	16'h	73d1;
4116	:douta	=	16'h	7413;
4117	:douta	=	16'h	e6b9;
4118	:douta	=	16'h	add9;
4119	:douta	=	16'h	d679;
4120	:douta	=	16'h	b597;
4121	:douta	=	16'h	7c54;
4122	:douta	=	16'h	ad97;
4123	:douta	=	16'h	a577;
4124	:douta	=	16'h	8453;
4125	:douta	=	16'h	8cb6;
4126	:douta	=	16'h	6b91;
4127	:douta	=	16'h	ad96;
4128	:douta	=	16'h	b5b8;
4129	:douta	=	16'h	b5b8;
4130	:douta	=	16'h	b5b8;
4131	:douta	=	16'h	a516;
4132	:douta	=	16'h	73d2;
4133	:douta	=	16'h	ad56;
4134	:douta	=	16'h	8cb6;
4135	:douta	=	16'h	ce38;
4136	:douta	=	16'h	deb9;
4137	:douta	=	16'h	9d16;
4138	:douta	=	16'h	c639;
4139	:douta	=	16'h	c617;
4140	:douta	=	16'h	b555;
4141	:douta	=	16'h	9d35;
4142	:douta	=	16'h	7c12;
4143	:douta	=	16'h	b5b6;
4144	:douta	=	16'h	d6b9;
4145	:douta	=	16'h	e6fa;
4146	:douta	=	16'h	8cd5;
4147	:douta	=	16'h	e6d9;
4148	:douta	=	16'h	c637;
4149	:douta	=	16'h	5b0e;
4150	:douta	=	16'h	5350;
4151	:douta	=	16'h	42ad;
4152	:douta	=	16'h	b594;
4153	:douta	=	16'h	bdb5;
4154	:douta	=	16'h	bdd6;
4155	:douta	=	16'h	d658;
4156	:douta	=	16'h	bd96;
4157	:douta	=	16'h	ad77;
4158	:douta	=	16'h	7390;
4159	:douta	=	16'h	8cd4;
4160	:douta	=	16'h	6b0e;
4161	:douta	=	16'h	eefa;
4162	:douta	=	16'h	b533;
4163	:douta	=	16'h	ffba;
4164	:douta	=	16'h	9cd4;
4165	:douta	=	16'h	7c33;
4166	:douta	=	16'h	bdd6;
4167	:douta	=	16'h	42cf;
4168	:douta	=	16'h	6b50;
4169	:douta	=	16'h	5b50;
4170	:douta	=	16'h	9d56;
4171	:douta	=	16'h	9516;
4172	:douta	=	16'h	e6d8;
4173	:douta	=	16'h	e75b;
4174	:douta	=	16'h	8cb5;
4175	:douta	=	16'h	d71c;
4176	:douta	=	16'h	859a;
4177	:douta	=	16'h	9453;
4178	:douta	=	16'h	6c55;
4179	:douta	=	16'h	63d3;
4180	:douta	=	16'h	94d5;
4181	:douta	=	16'h	ce38;
4182	:douta	=	16'h	9518;
4183	:douta	=	16'h	9538;
4184	:douta	=	16'h	ce9b;
4185	:douta	=	16'h	be7b;
4186	:douta	=	16'h	9d38;
4187	:douta	=	16'h	6c35;
4188	:douta	=	16'h	84d6;
4189	:douta	=	16'h	63f3;
4190	:douta	=	16'h	84b6;
4191	:douta	=	16'h	7c75;
4192	:douta	=	16'h	8d18;
4193	:douta	=	16'h	bdd9;
4194	:douta	=	16'h	be5a;
4195	:douta	=	16'h	6477;
4196	:douta	=	16'h	84b6;
4197	:douta	=	16'h	4acf;
4198	:douta	=	16'h	6bf2;
4199	:douta	=	16'h	7413;
4200	:douta	=	16'h	8517;
4201	:douta	=	16'h	84b7;
4202	:douta	=	16'h	be5a;
4203	:douta	=	16'h	957a;
4204	:douta	=	16'h	be3b;
4205	:douta	=	16'h	ae1c;
4206	:douta	=	16'h	7c56;
4207	:douta	=	16'h	8d59;
4208	:douta	=	16'h	6bf5;
4209	:douta	=	16'h	6435;
4210	:douta	=	16'h	32b0;
4211	:douta	=	16'h	63d2;
4212	:douta	=	16'h	63d2;
4213	:douta	=	16'h	8c72;
4214	:douta	=	16'h	8cb4;
4215	:douta	=	16'h	8cb5;
4216	:douta	=	16'h	de98;
4217	:douta	=	16'h	9d37;
4218	:douta	=	16'h	84d6;
4219	:douta	=	16'h	3a0c;
4220	:douta	=	16'h	530f;
4221	:douta	=	16'h	adfa;
4222	:douta	=	16'h	6391;
4223	:douta	=	16'h	94d4;
4224	:douta	=	16'h	9d15;
4225	:douta	=	16'h	8cb4;
4226	:douta	=	16'h	ad54;
4227	:douta	=	16'h	6b90;
4228	:douta	=	16'h	6bf2;
4229	:douta	=	16'h	7433;
4230	:douta	=	16'h	94d4;
4231	:douta	=	16'h	7454;
4232	:douta	=	16'h	f73b;
4233	:douta	=	16'h	c618;
4234	:douta	=	16'h	63d2;
4235	:douta	=	16'h	8453;
4236	:douta	=	16'h	3189;
4237	:douta	=	16'h	320a;
4238	:douta	=	16'h	3167;
4239	:douta	=	16'h	2924;
4240	:douta	=	16'h	20e3;
4241	:douta	=	16'h	1883;
4242	:douta	=	16'h	6b8f;
4243	:douta	=	16'h	7bd0;
4244	:douta	=	16'h	bdd6;
4245	:douta	=	16'h	9471;
4246	:douta	=	16'h	a533;
4247	:douta	=	16'h	2988;
4248	:douta	=	16'h	632e;
4249	:douta	=	16'h	0001;
4250	:douta	=	16'h	31c8;
4251	:douta	=	16'h	8c92;
4252	:douta	=	16'h	b574;
4253	:douta	=	16'h	d6b8;
4254	:douta	=	16'h	a556;
4255	:douta	=	16'h	a577;
4256	:douta	=	16'h	3a4c;
4257	:douta	=	16'h	21a8;
4258	:douta	=	16'h	3acc;
4259	:douta	=	16'h	2168;
4260	:douta	=	16'h	1126;
4261	:douta	=	16'h	08a4;
4262	:douta	=	16'h	0002;
4263	:douta	=	16'h	0042;
4264	:douta	=	16'h	0883;
4265	:douta	=	16'h	0884;
4266	:douta	=	16'h	08a4;
4267	:douta	=	16'h	08a4;
4268	:douta	=	16'h	10c5;
4269	:douta	=	16'h	08c4;
4270	:douta	=	16'h	0884;
4271	:douta	=	16'h	08a4;
4272	:douta	=	16'h	08c4;
4273	:douta	=	16'h	08a4;
4274	:douta	=	16'h	08a4;
4275	:douta	=	16'h	08a4;
4276	:douta	=	16'h	0884;
4277	:douta	=	16'h	08a4;
4278	:douta	=	16'h	08a4;
4279	:douta	=	16'h	08a4;
4280	:douta	=	16'h	08a4;
4281	:douta	=	16'h	0884;
4282	:douta	=	16'h	0884;
4283	:douta	=	16'h	0884;
4284	:douta	=	16'h	0884;
4285	:douta	=	16'h	0884;
4286	:douta	=	16'h	0883;
4287	:douta	=	16'h	0883;
4288	:douta	=	16'h	0883;
4289	:douta	=	16'h	0883;
4290	:douta	=	16'h	0883;
4291	:douta	=	16'h	0883;
4292	:douta	=	16'h	0883;
4293	:douta	=	16'h	0883;
4294	:douta	=	16'h	0883;
4295	:douta	=	16'h	08a4;
4296	:douta	=	16'h	0843;
4297	:douta	=	16'h	1083;
4298	:douta	=	16'h	0001;
4299	:douta	=	16'h	0002;
4300	:douta	=	16'h	0063;
4301	:douta	=	16'h	2a0a;
4302	:douta	=	16'h	63f1;
4303	:douta	=	16'h	53b5;
4304	:douta	=	16'h	ad98;
4305	:douta	=	16'h	8cb6;
4306	:douta	=	16'h	7414;
4307	:douta	=	16'h	4b31;
4308	:douta	=	16'h	3a8e;
4309	:douta	=	16'h	196a;
4310	:douta	=	16'h	3a8e;
4311	:douta	=	16'h	7474;
4312	:douta	=	16'h	7cb7;
4313	:douta	=	16'h	b597;
4314	:douta	=	16'h	84b8;
4315	:douta	=	16'h	6415;
4316	:douta	=	16'h	4394;
4317	:douta	=	16'h	2a90;
4318	:douta	=	16'h	7cf9;
4319	:douta	=	16'h	3ab0;
4320	:douta	=	16'h	4311;
4321	:douta	=	16'h	3ad1;
4322	:douta	=	16'h	3ad0;
4323	:douta	=	16'h	3ad0;
4324	:douta	=	16'h	6c35;
4325	:douta	=	16'h	8cd6;
4326	:douta	=	16'h	8cb6;
4327	:douta	=	16'h	9559;
4328	:douta	=	16'h	7414;
4329	:douta	=	16'h	2a4d;
4330	:douta	=	16'h	6bf4;
4331	:douta	=	16'h	5bb3;
4332	:douta	=	16'h	7cb6;
4333	:douta	=	16'h	8cb6;
4334	:douta	=	16'h	5bd4;
4335	:douta	=	16'h	7c96;
4336	:douta	=	16'h	5bd3;
4337	:douta	=	16'h	3ad1;
4338	:douta	=	16'h	5bb4;
4339	:douta	=	16'h	114a;
4340	:douta	=	16'h	4310;
4341	:douta	=	16'h	8d5a;
4342	:douta	=	16'h	9579;
4343	:douta	=	16'h	5417;
4344	:douta	=	16'h	63f5;
4345	:douta	=	16'h	4394;
4346	:douta	=	16'h	0a0e;
4347	:douta	=	16'h	3b53;
4348	:douta	=	16'h	3b54;
4349	:douta	=	16'h	8d5a;
4350	:douta	=	16'h	74da;
4351	:douta	=	16'h	853a;
4352	:douta	=	16'h	6cba;
4353	:douta	=	16'h	6c98;
4354	:douta	=	16'h	6cb8;
4355	:douta	=	16'h	4b33;
4356	:douta	=	16'h	2a70;
4357	:douta	=	16'h	4332;
4358	:douta	=	16'h	5351;
4359	:douta	=	16'h	6c15;
4360	:douta	=	16'h	84d8;
4361	:douta	=	16'h	5bb4;
4362	:douta	=	16'h	6bf3;
4363	:douta	=	16'h	8495;
4364	:douta	=	16'h	5b71;
4365	:douta	=	16'h	63d3;
4366	:douta	=	16'h	5371;
4367	:douta	=	16'h	6bd2;
4368	:douta	=	16'h	ad56;
4369	:douta	=	16'h	9d36;
4370	:douta	=	16'h	ce39;
4371	:douta	=	16'h	9d36;
4372	:douta	=	16'h	9d57;
4373	:douta	=	16'h	9cd4;
4374	:douta	=	16'h	7413;
4375	:douta	=	16'h	6bf4;
4376	:douta	=	16'h	8c72;
4377	:douta	=	16'h	ad56;
4378	:douta	=	16'h	b5b7;
4379	:douta	=	16'h	9d16;
4380	:douta	=	16'h	c5f7;
4381	:douta	=	16'h	ce59;
4382	:douta	=	16'h	b577;
4383	:douta	=	16'h	be19;
4384	:douta	=	16'h	7c14;
4385	:douta	=	16'h	94f5;
4386	:douta	=	16'h	7c74;
4387	:douta	=	16'h	63d2;
4388	:douta	=	16'h	a536;
4389	:douta	=	16'h	d699;
4390	:douta	=	16'h	b5d9;
4391	:douta	=	16'h	f77c;
4392	:douta	=	16'h	8cb5;
4393	:douta	=	16'h	9cd4;
4394	:douta	=	16'h	8453;
4395	:douta	=	16'h	a515;
4396	:douta	=	16'h	d678;
4397	:douta	=	16'h	d6b9;
4398	:douta	=	16'h	c5f6;
4399	:douta	=	16'h	ef3b;
4400	:douta	=	16'h	8455;
4401	:douta	=	16'h	94d4;
4402	:douta	=	16'h	4acf;
4403	:douta	=	16'h	cdf6;
4404	:douta	=	16'h	c5d5;
4405	:douta	=	16'h	d657;
4406	:douta	=	16'h	bdd5;
4407	:douta	=	16'h	cdf6;
4408	:douta	=	16'h	deb8;
4409	:douta	=	16'h	7c32;
4410	:douta	=	16'h	8c94;
4411	:douta	=	16'h	7bb0;
4412	:douta	=	16'h	c5f6;
4413	:douta	=	16'h	8492;
4414	:douta	=	16'h	73d0;
4415	:douta	=	16'h	b595;
4416	:douta	=	16'h	ef3a;
4417	:douta	=	16'h	ef3a;
4418	:douta	=	16'h	6bd2;
4419	:douta	=	16'h	83d0;
4420	:douta	=	16'h	534f;
4421	:douta	=	16'h	6b6f;
4422	:douta	=	16'h	ce37;
4423	:douta	=	16'h	9472;
4424	:douta	=	16'h	ff7b;
4425	:douta	=	16'h	7413;
4426	:douta	=	16'h	d6ba;
4427	:douta	=	16'h	6c35;
4428	:douta	=	16'h	9c92;
4429	:douta	=	16'h	7c94;
4430	:douta	=	16'h	530f;
4431	:douta	=	16'h	8cf5;
4432	:douta	=	16'h	63b2;
4433	:douta	=	16'h	c698;
4434	:douta	=	16'h	9517;
4435	:douta	=	16'h	d67a;
4436	:douta	=	16'h	7cb6;
4437	:douta	=	16'h	8cd6;
4438	:douta	=	16'h	4bd4;
4439	:douta	=	16'h	5c36;
4440	:douta	=	16'h	a577;
4441	:douta	=	16'h	7c95;
4442	:douta	=	16'h	84b6;
4443	:douta	=	16'h	7435;
4444	:douta	=	16'h	9d58;
4445	:douta	=	16'h	cedd;
4446	:douta	=	16'h	6c56;
4447	:douta	=	16'h	6c55;
4448	:douta	=	16'h	5372;
4449	:douta	=	16'h	94d5;
4450	:douta	=	16'h	4b73;
4451	:douta	=	16'h	428e;
4452	:douta	=	16'h	63f3;
4453	:douta	=	16'h	adfa;
4454	:douta	=	16'h	a599;
4455	:douta	=	16'h	d6bb;
4456	:douta	=	16'h	ae1c;
4457	:douta	=	16'h	5b73;
4458	:douta	=	16'h	9518;
4459	:douta	=	16'h	7435;
4460	:douta	=	16'h	4b73;
4461	:douta	=	16'h	4353;
4462	:douta	=	16'h	a578;
4463	:douta	=	16'h	8d39;
4464	:douta	=	16'h	8d38;
4465	:douta	=	16'h	53d5;
4466	:douta	=	16'h	74b7;
4467	:douta	=	16'h	deba;
4468	:douta	=	16'h	8cd7;
4469	:douta	=	16'h	6b91;
4470	:douta	=	16'h	3a6e;
4471	:douta	=	16'h	420a;
4472	:douta	=	16'h	7433;
4473	:douta	=	16'h	7433;
4474	:douta	=	16'h	5b91;
4475	:douta	=	16'h	7433;
4476	:douta	=	16'h	73f3;
4477	:douta	=	16'h	adda;
4478	:douta	=	16'h	bdb7;
4479	:douta	=	16'h	8474;
4480	:douta	=	16'h	6390;
4481	:douta	=	16'h	73b1;
4482	:douta	=	16'h	8cd5;
4483	:douta	=	16'h	b619;
4484	:douta	=	16'h	a598;
4485	:douta	=	16'h	a4d4;
4486	:douta	=	16'h	ce38;
4487	:douta	=	16'h	7b6e;
4488	:douta	=	16'h	4aad;
4489	:douta	=	16'h	426d;
4490	:douta	=	16'h	4ace;
4491	:douta	=	16'h	6391;
4492	:douta	=	16'h	b5d7;
4493	:douta	=	16'h	428d;
4494	:douta	=	16'h	a536;
4495	:douta	=	16'h	18c3;
4496	:douta	=	16'h	2104;
4497	:douta	=	16'h	18c4;
4498	:douta	=	16'h	52cd;
4499	:douta	=	16'h	2988;
4500	:douta	=	16'h	29c9;
4501	:douta	=	16'h	4a8b;
4502	:douta	=	16'h	6baf;
4503	:douta	=	16'h	8c51;
4504	:douta	=	16'h	eefa;
4505	:douta	=	16'h	8c10;
4506	:douta	=	16'h	cdf6;
4507	:douta	=	16'h	3a6b;
4508	:douta	=	16'h	42cc;
4509	:douta	=	16'h	0083;
4510	:douta	=	16'h	08a3;
4511	:douta	=	16'h	0062;
4512	:douta	=	16'h	0883;
4513	:douta	=	16'h	08a3;
4514	:douta	=	16'h	08a4;
4515	:douta	=	16'h	08a5;
4516	:douta	=	16'h	10c5;
4517	:douta	=	16'h	08a4;
4518	:douta	=	16'h	10e5;
4519	:douta	=	16'h	08c4;
4520	:douta	=	16'h	10c5;
4521	:douta	=	16'h	10c5;
4522	:douta	=	16'h	08c4;
4523	:douta	=	16'h	10c5;
4524	:douta	=	16'h	0884;
4525	:douta	=	16'h	0063;
4526	:douta	=	16'h	0042;
4527	:douta	=	16'h	0042;
4528	:douta	=	16'h	0042;
4529	:douta	=	16'h	0022;
4530	:douta	=	16'h	0863;
4531	:douta	=	16'h	0883;
4532	:douta	=	16'h	10a4;
4533	:douta	=	16'h	10c5;
4534	:douta	=	16'h	10e5;
4535	:douta	=	16'h	1906;
4536	:douta	=	16'h	1905;
4537	:douta	=	16'h	1906;
4538	:douta	=	16'h	2127;
4539	:douta	=	16'h	1906;
4540	:douta	=	16'h	10a4;
4541	:douta	=	16'h	08a4;
4542	:douta	=	16'h	0883;
4543	:douta	=	16'h	0862;
4544	:douta	=	16'h	0022;
4545	:douta	=	16'h	0001;
4546	:douta	=	16'h	0021;
4547	:douta	=	16'h	0041;
4548	:douta	=	16'h	0882;
4549	:douta	=	16'h	0883;
4550	:douta	=	16'h	0884;
4551	:douta	=	16'h	0884;
4552	:douta	=	16'h	0884;
4553	:douta	=	16'h	10a4;
4554	:douta	=	16'h	0884;
4555	:douta	=	16'h	0884;
4556	:douta	=	16'h	0884;
4557	:douta	=	16'h	0883;
4558	:douta	=	16'h	0883;
4559	:douta	=	16'h	0862;
4560	:douta	=	16'h	0001;
4561	:douta	=	16'h	0043;
4562	:douta	=	16'h	220a;
4563	:douta	=	16'h	326c;
4564	:douta	=	16'h	b5b8;
4565	:douta	=	16'h	8495;
4566	:douta	=	16'h	a557;
4567	:douta	=	16'h	09ac;
4568	:douta	=	16'h	1948;
4569	:douta	=	16'h	4b74;
4570	:douta	=	16'h	21ec;
4571	:douta	=	16'h	5393;
4572	:douta	=	16'h	3b12;
4573	:douta	=	16'h	6c56;
4574	:douta	=	16'h	be1b;
4575	:douta	=	16'h	7497;
4576	:douta	=	16'h	3af1;
4577	:douta	=	16'h	9559;
4578	:douta	=	16'h	2a6f;
4579	:douta	=	16'h	4b31;
4580	:douta	=	16'h	2a4e;
4581	:douta	=	16'h	21cc;
4582	:douta	=	16'h	7c54;
4583	:douta	=	16'h	324d;
4584	:douta	=	16'h	7454;
4585	:douta	=	16'h	63f4;
4586	:douta	=	16'h	8d16;
4587	:douta	=	16'h	5bd3;
4588	:douta	=	16'h	5bd3;
4589	:douta	=	16'h	4332;
4590	:douta	=	16'h	42ae;
4591	:douta	=	16'h	7cb6;
4592	:douta	=	16'h	7c75;
4593	:douta	=	16'h	b5f8;
4594	:douta	=	16'h	4b52;
4595	:douta	=	16'h	7cd9;
4596	:douta	=	16'h	222f;
4597	:douta	=	16'h	224f;
4598	:douta	=	16'h	2ab1;
4599	:douta	=	16'h	5bb4;
4600	:douta	=	16'h	ae1c;
4601	:douta	=	16'h	7cb9;
4602	:douta	=	16'h	a63f;
4603	:douta	=	16'h	53d6;
4604	:douta	=	16'h	5c17;
4605	:douta	=	16'h	1a4f;
4606	:douta	=	16'h	6436;
4607	:douta	=	16'h	5c37;
4608	:douta	=	16'h	32f2;
4609	:douta	=	16'h	5332;
4610	:douta	=	16'h	6436;
4611	:douta	=	16'h	6437;
4612	:douta	=	16'h	6c98;
4613	:douta	=	16'h	4b94;
4614	:douta	=	16'h	21ac;
4615	:douta	=	16'h	5393;
4616	:douta	=	16'h	4b32;
4617	:douta	=	16'h	4b32;
4618	:douta	=	16'h	4aef;
4619	:douta	=	16'h	9d58;
4620	:douta	=	16'h	7c75;
4621	:douta	=	16'h	a579;
4622	:douta	=	16'h	5b72;
4623	:douta	=	16'h	6bd2;
4624	:douta	=	16'h	5393;
4625	:douta	=	16'h	6392;
4626	:douta	=	16'h	8476;
4627	:douta	=	16'h	b5b8;
4628	:douta	=	16'h	a577;
4629	:douta	=	16'h	de99;
4630	:douta	=	16'h	be3a;
4631	:douta	=	16'h	ad77;
4632	:douta	=	16'h	5b2f;
4633	:douta	=	16'h	8434;
4634	:douta	=	16'h	73f2;
4635	:douta	=	16'h	7c74;
4636	:douta	=	16'h	a536;
4637	:douta	=	16'h	63d2;
4638	:douta	=	16'h	a536;
4639	:douta	=	16'h	bdf7;
4640	:douta	=	16'h	c5f7;
4641	:douta	=	16'h	d659;
4642	:douta	=	16'h	a577;
4643	:douta	=	16'h	7c33;
4644	:douta	=	16'h	5b51;
4645	:douta	=	16'h	9cf6;
4646	:douta	=	16'h	9d57;
4647	:douta	=	16'h	eefa;
4648	:douta	=	16'h	deb9;
4649	:douta	=	16'h	ce17;
4650	:douta	=	16'h	94f5;
4651	:douta	=	16'h	a514;
4652	:douta	=	16'h	a4f4;
4653	:douta	=	16'h	8453;
4654	:douta	=	16'h	9cb4;
4655	:douta	=	16'h	e719;
4656	:douta	=	16'h	b576;
4657	:douta	=	16'h	ef7b;
4658	:douta	=	16'h	5b71;
4659	:douta	=	16'h	cdf5;
4660	:douta	=	16'h	bdd7;
4661	:douta	=	16'h	9492;
4662	:douta	=	16'h	7c52;
4663	:douta	=	16'h	a4d3;
4664	:douta	=	16'h	ef19;
4665	:douta	=	16'h	ad54;
4666	:douta	=	16'h	ce77;
4667	:douta	=	16'h	c5d6;
4668	:douta	=	16'h	ce77;
4669	:douta	=	16'h	328e;
4670	:douta	=	16'h	0085;
4671	:douta	=	16'h	532e;
4672	:douta	=	16'h	bdd5;
4673	:douta	=	16'h	e6d9;
4674	:douta	=	16'h	cdb5;
4675	:douta	=	16'h	ff19;
4676	:douta	=	16'h	4b0f;
4677	:douta	=	16'h	6b0e;
4678	:douta	=	16'h	b556;
4679	:douta	=	16'h	39ea;
4680	:douta	=	16'h	ad13;
4681	:douta	=	16'h	8cb4;
4682	:douta	=	16'h	d6b9;
4683	:douta	=	16'h	9536;
4684	:douta	=	16'h	ff9b;
4685	:douta	=	16'h	a598;
4686	:douta	=	16'h	6371;
4687	:douta	=	16'h	7c95;
4688	:douta	=	16'h	42d0;
4689	:douta	=	16'h	84d5;
4690	:douta	=	16'h	5351;
4691	:douta	=	16'h	b5b7;
4692	:douta	=	16'h	c659;
4693	:douta	=	16'h	c638;
4694	:douta	=	16'h	5394;
4695	:douta	=	16'h	5b93;
4696	:douta	=	16'h	6c14;
4697	:douta	=	16'h	32af;
4698	:douta	=	16'h	4331;
4699	:douta	=	16'h	8495;
4700	:douta	=	16'h	84f7;
4701	:douta	=	16'h	9599;
4702	:douta	=	16'h	9d99;
4703	:douta	=	16'h	7cd7;
4704	:douta	=	16'h	8d17;
4705	:douta	=	16'h	ce39;
4706	:douta	=	16'h	64d9;
4707	:douta	=	16'h	3a2f;
4708	:douta	=	16'h	5bd3;
4709	:douta	=	16'h	7455;
4710	:douta	=	16'h	6bf3;
4711	:douta	=	16'h	be1a;
4712	:douta	=	16'h	8d18;
4713	:douta	=	16'h	7497;
4714	:douta	=	16'h	cedc;
4715	:douta	=	16'h	9579;
4716	:douta	=	16'h	74b8;
4717	:douta	=	16'h	2ad2;
4718	:douta	=	16'h	ce59;
4719	:douta	=	16'h	8d18;
4720	:douta	=	16'h	4310;
4721	:douta	=	16'h	4b52;
4722	:douta	=	16'h	5332;
4723	:douta	=	16'h	a576;
4724	:douta	=	16'h	94b5;
4725	:douta	=	16'h	b597;
4726	:douta	=	16'h	7414;
4727	:douta	=	16'h	9452;
4728	:douta	=	16'h	9537;
4729	:douta	=	16'h	84b4;
4730	:douta	=	16'h	42cf;
4731	:douta	=	16'h	5b2f;
4732	:douta	=	16'h	6b90;
4733	:douta	=	16'h	8495;
4734	:douta	=	16'h	a576;
4735	:douta	=	16'h	73f3;
4736	:douta	=	16'h	8cb4;
4737	:douta	=	16'h	94b4;
4738	:douta	=	16'h	5b2f;
4739	:douta	=	16'h	94d5;
4740	:douta	=	16'h	532f;
4741	:douta	=	16'h	b5d7;
4742	:douta	=	16'h	b5f7;
4743	:douta	=	16'h	de99;
4744	:douta	=	16'h	6391;
4745	:douta	=	16'h	29eb;
4746	:douta	=	16'h	6371;
4747	:douta	=	16'h	29ea;
4748	:douta	=	16'h	6370;
4749	:douta	=	16'h	5b50;
4750	:douta	=	16'h	5b2f;
4751	:douta	=	16'h	3986;
4752	:douta	=	16'h	18e3;
4753	:douta	=	16'h	20e5;
4754	:douta	=	16'h	528c;
4755	:douta	=	16'h	a4d4;
4756	:douta	=	16'h	422b;
4757	:douta	=	16'h	5aed;
4758	:douta	=	16'h	3a4b;
4759	:douta	=	16'h	4aac;
4760	:douta	=	16'h	7c72;
4761	:douta	=	16'h	6baf;
4762	:douta	=	16'h	8cb2;
4763	:douta	=	16'h	29c8;
4764	:douta	=	16'h	0083;
4765	:douta	=	16'h	10a4;
4766	:douta	=	16'h	08a4;
4767	:douta	=	16'h	10a4;
4768	:douta	=	16'h	10a4;
4769	:douta	=	16'h	18c5;
4770	:douta	=	16'h	10e4;
4771	:douta	=	16'h	10c5;
4772	:douta	=	16'h	10a5;
4773	:douta	=	16'h	10c5;
4774	:douta	=	16'h	08a4;
4775	:douta	=	16'h	08a4;
4776	:douta	=	16'h	0883;
4777	:douta	=	16'h	0883;
4778	:douta	=	16'h	0062;
4779	:douta	=	16'h	0042;
4780	:douta	=	16'h	10a4;
4781	:douta	=	16'h	1926;
4782	:douta	=	16'h	2168;
4783	:douta	=	16'h	29a9;
4784	:douta	=	16'h	31ca;
4785	:douta	=	16'h	3a0c;
4786	:douta	=	16'h	3a4c;
4787	:douta	=	16'h	3a6c;
4788	:douta	=	16'h	4aef;
4789	:douta	=	16'h	42ae;
4790	:douta	=	16'h	4aaf;
4791	:douta	=	16'h	428f;
4792	:douta	=	16'h	428f;
4793	:douta	=	16'h	3a6d;
4794	:douta	=	16'h	42ae;
4795	:douta	=	16'h	426d;
4796	:douta	=	16'h	3a2c;
4797	:douta	=	16'h	322c;
4798	:douta	=	16'h	3a2b;
4799	:douta	=	16'h	320b;
4800	:douta	=	16'h	31ca;
4801	:douta	=	16'h	29ca;
4802	:douta	=	16'h	29a9;
4803	:douta	=	16'h	1926;
4804	:douta	=	16'h	10e5;
4805	:douta	=	16'h	0843;
4806	:douta	=	16'h	0062;
4807	:douta	=	16'h	0041;
4808	:douta	=	16'h	0882;
4809	:douta	=	16'h	0883;
4810	:douta	=	16'h	0884;
4811	:douta	=	16'h	08c3;
4812	:douta	=	16'h	08a3;
4813	:douta	=	16'h	0884;
4814	:douta	=	16'h	08a4;
4815	:douta	=	16'h	08a4;
4816	:douta	=	16'h	0883;
4817	:douta	=	16'h	0883;
4818	:douta	=	16'h	0000;
4819	:douta	=	16'h	0000;
4820	:douta	=	16'h	21ea;
4821	:douta	=	16'h	8cd5;
4822	:douta	=	16'h	8518;
4823	:douta	=	16'h	4b30;
4824	:douta	=	16'h	94f6;
4825	:douta	=	16'h	3af1;
4826	:douta	=	16'h	19ac;
4827	:douta	=	16'h	19cd;
4828	:douta	=	16'h	2a90;
4829	:douta	=	16'h	094b;
4830	:douta	=	16'h	7475;
4831	:douta	=	16'h	3b11;
4832	:douta	=	16'h	6c14;
4833	:douta	=	16'h	7435;
4834	:douta	=	16'h	5352;
4835	:douta	=	16'h	63f4;
4836	:douta	=	16'h	324e;
4837	:douta	=	16'h	3aaf;
4838	:douta	=	16'h	3a6e;
4839	:douta	=	16'h	4b2f;
4840	:douta	=	16'h	21ec;
4841	:douta	=	16'h	5331;
4842	:douta	=	16'h	6c34;
4843	:douta	=	16'h	9d79;
4844	:douta	=	16'h	9d79;
4845	:douta	=	16'h	4b32;
4846	:douta	=	16'h	3ad0;
4847	:douta	=	16'h	224f;
4848	:douta	=	16'h	4b32;
4849	:douta	=	16'h	5bd3;
4850	:douta	=	16'h	63d3;
4851	:douta	=	16'h	4b53;
4852	:douta	=	16'h	4b73;
4853	:douta	=	16'h	4b95;
4854	:douta	=	16'h	2250;
4855	:douta	=	16'h	3312;
4856	:douta	=	16'h	6c56;
4857	:douta	=	16'h	9dba;
4858	:douta	=	16'h	6cdb;
4859	:douta	=	16'h	6c57;
4860	:douta	=	16'h	6cdb;
4861	:douta	=	16'h	6457;
4862	:douta	=	16'h	5c58;
4863	:douta	=	16'h	1a0e;
4864	:douta	=	16'h	7d5c;
4865	:douta	=	16'h	326f;
4866	:douta	=	16'h	6c57;
4867	:douta	=	16'h	3af1;
4868	:douta	=	16'h	4332;
4869	:douta	=	16'h	2a4f;
4870	:douta	=	16'h	6c35;
4871	:douta	=	16'h	84f9;
4872	:douta	=	16'h	74b7;
4873	:douta	=	16'h	7435;
4874	:douta	=	16'h	8495;
4875	:douta	=	16'h	5331;
4876	:douta	=	16'h	4b30;
4877	:douta	=	16'h	63b2;
4878	:douta	=	16'h	5330;
4879	:douta	=	16'h	6350;
4880	:douta	=	16'h	9d37;
4881	:douta	=	16'h	a578;
4882	:douta	=	16'h	84d7;
4883	:douta	=	16'h	a555;
4884	:douta	=	16'h	94d5;
4885	:douta	=	16'h	8433;
4886	:douta	=	16'h	8454;
4887	:douta	=	16'h	7413;
4888	:douta	=	16'h	8c73;
4889	:douta	=	16'h	9d15;
4890	:douta	=	16'h	b597;
4891	:douta	=	16'h	a576;
4892	:douta	=	16'h	de99;
4893	:douta	=	16'h	be1a;
4894	:douta	=	16'h	9cf5;
4895	:douta	=	16'h	9516;
4896	:douta	=	16'h	6bb2;
4897	:douta	=	16'h	9d35;
4898	:douta	=	16'h	a4f4;
4899	:douta	=	16'h	9cf3;
4900	:douta	=	16'h	bdd8;
4901	:douta	=	16'h	e6da;
4902	:douta	=	16'h	94d5;
4903	:douta	=	16'h	d699;
4904	:douta	=	16'h	94f4;
4905	:douta	=	16'h	bd96;
4906	:douta	=	16'h	b5d7;
4907	:douta	=	16'h	a514;
4908	:douta	=	16'h	b595;
4909	:douta	=	16'h	de99;
4910	:douta	=	16'h	ce38;
4911	:douta	=	16'h	ded9;
4912	:douta	=	16'h	ad55;
4913	:douta	=	16'h	6bf1;
4914	:douta	=	16'h	4ace;
4915	:douta	=	16'h	ce16;
4916	:douta	=	16'h	c5f6;
4917	:douta	=	16'h	eed7;
4918	:douta	=	16'h	9d15;
4919	:douta	=	16'h	8411;
4920	:douta	=	16'h	bdb5;
4921	:douta	=	16'h	9d14;
4922	:douta	=	16'h	3aae;
4923	:douta	=	16'h	c5d4;
4924	:douta	=	16'h	e6d8;
4925	:douta	=	16'h	bd73;
4926	:douta	=	16'h	d617;
4927	:douta	=	16'h	8431;
4928	:douta	=	16'h	eeb8;
4929	:douta	=	16'h	7432;
4930	:douta	=	16'h	9471;
4931	:douta	=	16'h	94b2;
4932	:douta	=	16'h	5b0b;
4933	:douta	=	16'h	bd95;
4934	:douta	=	16'h	f77a;
4935	:douta	=	16'h	bd75;
4936	:douta	=	16'h	fffc;
4937	:douta	=	16'h	6370;
4938	:douta	=	16'h	a514;
4939	:douta	=	16'h	4b50;
4940	:douta	=	16'h	8452;
4941	:douta	=	16'h	9515;
4942	:douta	=	16'h	bdf8;
4943	:douta	=	16'h	a5b8;
4944	:douta	=	16'h	8475;
4945	:douta	=	16'h	ce78;
4946	:douta	=	16'h	7474;
4947	:douta	=	16'h	b577;
4948	:douta	=	16'h	52ce;
4949	:douta	=	16'h	7c74;
4950	:douta	=	16'h	9537;
4951	:douta	=	16'h	b63b;
4952	:douta	=	16'h	9579;
4953	:douta	=	16'h	5bd5;
4954	:douta	=	16'h	ae1a;
4955	:douta	=	16'h	7497;
4956	:douta	=	16'h	94f6;
4957	:douta	=	16'h	5c15;
4958	:douta	=	16'h	3a8f;
4959	:douta	=	16'h	32b0;
4960	:douta	=	16'h	6c14;
4961	:douta	=	16'h	9d78;
4962	:douta	=	16'h	63f4;
4963	:douta	=	16'h	9578;
4964	:douta	=	16'h	6c56;
4965	:douta	=	16'h	c67b;
4966	:douta	=	16'h	7476;
4967	:douta	=	16'h	a61b;
4968	:douta	=	16'h	53d4;
4969	:douta	=	16'h	6c35;
4970	:douta	=	16'h	5b93;
4971	:douta	=	16'h	7c96;
4972	:douta	=	16'h	2a6f;
4973	:douta	=	16'h	7476;
4974	:douta	=	16'h	c65a;
4975	:douta	=	16'h	8518;
4976	:douta	=	16'h	957a;
4977	:douta	=	16'h	3b33;
4978	:douta	=	16'h	9cd6;
4979	:douta	=	16'h	adfa;
4980	:douta	=	16'h	a556;
4981	:douta	=	16'h	9d56;
4982	:douta	=	16'h	3a4c;
4983	:douta	=	16'h	9cd3;
4984	:douta	=	16'h	5350;
4985	:douta	=	16'h	5b92;
4986	:douta	=	16'h	42f0;
4987	:douta	=	16'h	8d37;
4988	:douta	=	16'h	9d16;
4989	:douta	=	16'h	7c95;
4990	:douta	=	16'h	bdd8;
4991	:douta	=	16'h	5330;
4992	:douta	=	16'h	73b0;
4993	:douta	=	16'h	8473;
4994	:douta	=	16'h	7413;
4995	:douta	=	16'h	8d77;
4996	:douta	=	16'h	84d6;
4997	:douta	=	16'h	b595;
4998	:douta	=	16'h	7413;
4999	:douta	=	16'h	7cb5;
5000	:douta	=	16'h	6bf2;
5001	:douta	=	16'h	6bf2;
5002	:douta	=	16'h	9d56;
5003	:douta	=	16'h	5b72;
5004	:douta	=	16'h	be5b;
5005	:douta	=	16'h	8474;
5006	:douta	=	16'h	6bd1;
5007	:douta	=	16'h	6b4d;
5008	:douta	=	16'h	20e4;
5009	:douta	=	16'h	20e4;
5010	:douta	=	16'h	2145;
5011	:douta	=	16'h	5b0d;
5012	:douta	=	16'h	9d34;
5013	:douta	=	16'h	ce58;
5014	:douta	=	16'h	7411;
5015	:douta	=	16'h	4aac;
5016	:douta	=	16'h	10c5;
5017	:douta	=	16'h	08c3;
5018	:douta	=	16'h	0884;
5019	:douta	=	16'h	10e4;
5020	:douta	=	16'h	10c4;
5021	:douta	=	16'h	10e4;
5022	:douta	=	16'h	10c5;
5023	:douta	=	16'h	10e5;
5024	:douta	=	16'h	10e4;
5025	:douta	=	16'h	08a4;
5026	:douta	=	16'h	0063;
5027	:douta	=	16'h	0862;
5028	:douta	=	16'h	1084;
5029	:douta	=	16'h	2967;
5030	:douta	=	16'h	29c9;
5031	:douta	=	16'h	3a2b;
5032	:douta	=	16'h	4a8e;
5033	:douta	=	16'h	6331;
5034	:douta	=	16'h	4ace;
5035	:douta	=	16'h	5b72;
5036	:douta	=	16'h	4b51;
5037	:douta	=	16'h	5bb4;
5038	:douta	=	16'h	6415;
5039	:douta	=	16'h	63f6;
5040	:douta	=	16'h	6c56;
5041	:douta	=	16'h	6437;
5042	:douta	=	16'h	6415;
5043	:douta	=	16'h	6c57;
5044	:douta	=	16'h	6c57;
5045	:douta	=	16'h	6c78;
5046	:douta	=	16'h	74d9;
5047	:douta	=	16'h	6c98;
5048	:douta	=	16'h	7d1a;
5049	:douta	=	16'h	853b;
5050	:douta	=	16'h	7d1a;
5051	:douta	=	16'h	7cf9;
5052	:douta	=	16'h	853a;
5053	:douta	=	16'h	74b9;
5054	:douta	=	16'h	6456;
5055	:douta	=	16'h	6c57;
5056	:douta	=	16'h	6416;
5057	:douta	=	16'h	6c36;
5058	:douta	=	16'h	63f5;
5059	:douta	=	16'h	5b93;
5060	:douta	=	16'h	5372;
5061	:douta	=	16'h	4b10;
5062	:douta	=	16'h	426e;
5063	:douta	=	16'h	322d;
5064	:douta	=	16'h	3aae;
5065	:douta	=	16'h	2a0b;
5066	:douta	=	16'h	21a9;
5067	:douta	=	16'h	10e5;
5068	:douta	=	16'h	1084;
5069	:douta	=	16'h	0062;
5070	:douta	=	16'h	0042;
5071	:douta	=	16'h	0883;
5072	:douta	=	16'h	08a3;
5073	:douta	=	16'h	0884;
5074	:douta	=	16'h	08a4;
5075	:douta	=	16'h	08c4;
5076	:douta	=	16'h	08a4;
5077	:douta	=	16'h	0022;
5078	:douta	=	16'h	0001;
5079	:douta	=	16'h	29e9;
5080	:douta	=	16'h	42cf;
5081	:douta	=	16'h	6c76;
5082	:douta	=	16'h	6415;
5083	:douta	=	16'h	6c54;
5084	:douta	=	16'h	9538;
5085	:douta	=	16'h	6416;
5086	:douta	=	16'h	6415;
5087	:douta	=	16'h	1128;
5088	:douta	=	16'h	42d1;
5089	:douta	=	16'h	2a4e;
5090	:douta	=	16'h	42ce;
5091	:douta	=	16'h	63f3;
5092	:douta	=	16'h	ad56;
5093	:douta	=	16'h	a536;
5094	:douta	=	16'h	7c34;
5095	:douta	=	16'h	5b72;
5096	:douta	=	16'h	3a6f;
5097	:douta	=	16'h	3a8e;
5098	:douta	=	16'h	3ad0;
5099	:douta	=	16'h	116a;
5100	:douta	=	16'h	4310;
5101	:douta	=	16'h	63d3;
5102	:douta	=	16'h	6c34;
5103	:douta	=	16'h	7455;
5104	:douta	=	16'h	5bf5;
5105	:douta	=	16'h	224f;
5106	:douta	=	16'h	222e;
5107	:douta	=	16'h	5b92;
5108	:douta	=	16'h	7455;
5109	:douta	=	16'h	53b4;
5110	:douta	=	16'h	8cd6;
5111	:douta	=	16'h	5c58;
5112	:douta	=	16'h	7d1a;
5113	:douta	=	16'h	3355;
5114	:douta	=	16'h	5bf6;
5115	:douta	=	16'h	6cb9;
5116	:douta	=	16'h	3b33;
5117	:douta	=	16'h	7d19;
5118	:douta	=	16'h	6458;
5119	:douta	=	16'h	959b;
5120	:douta	=	16'h	6478;
5121	:douta	=	16'h	3a8f;
5122	:douta	=	16'h	6c36;
5123	:douta	=	16'h	5c16;
5124	:douta	=	16'h	4312;
5125	:douta	=	16'h	3af1;
5126	:douta	=	16'h	5371;
5127	:douta	=	16'h	3a8e;
5128	:douta	=	16'h	84d8;
5129	:douta	=	16'h	5331;
5130	:douta	=	16'h	8d17;
5131	:douta	=	16'h	8495;
5132	:douta	=	16'h	6bf4;
5133	:douta	=	16'h	7434;
5134	:douta	=	16'h	428d;
5135	:douta	=	16'h	6370;
5136	:douta	=	16'h	5351;
5137	:douta	=	16'h	63d2;
5138	:douta	=	16'h	8497;
5139	:douta	=	16'h	deba;
5140	:douta	=	16'h	be19;
5141	:douta	=	16'h	de99;
5142	:douta	=	16'h	c67a;
5143	:douta	=	16'h	8454;
5144	:douta	=	16'h	9452;
5145	:douta	=	16'h	a515;
5146	:douta	=	16'h	42d0;
5147	:douta	=	16'h	32ae;
5148	:douta	=	16'h	94f5;
5149	:douta	=	16'h	d6ba;
5150	:douta	=	16'h	c5f8;
5151	:douta	=	16'h	c639;
5152	:douta	=	16'h	b577;
5153	:douta	=	16'h	b5d8;
5154	:douta	=	16'h	8453;
5155	:douta	=	16'h	73d1;
5156	:douta	=	16'h	94d5;
5157	:douta	=	16'h	bdb7;
5158	:douta	=	16'h	ce37;
5159	:douta	=	16'h	ef5b;
5160	:douta	=	16'h	d679;
5161	:douta	=	16'h	d678;
5162	:douta	=	16'h	a556;
5163	:douta	=	16'h	a535;
5164	:douta	=	16'h	9473;
5165	:douta	=	16'h	bdf7;
5166	:douta	=	16'h	ce38;
5167	:douta	=	16'h	ef1a;
5168	:douta	=	16'h	de78;
5169	:douta	=	16'h	d698;
5170	:douta	=	16'h	6391;
5171	:douta	=	16'h	ad13;
5172	:douta	=	16'h	8cb3;
5173	:douta	=	16'h	deb8;
5174	:douta	=	16'h	b574;
5175	:douta	=	16'h	ce15;
5176	:douta	=	16'h	d678;
5177	:douta	=	16'h	8451;
5178	:douta	=	16'h	9d35;
5179	:douta	=	16'h	734e;
5180	:douta	=	16'h	9c70;
5181	:douta	=	16'h	bdd5;
5182	:douta	=	16'h	52a9;
5183	:douta	=	16'h	c5f4;
5184	:douta	=	16'h	f75a;
5185	:douta	=	16'h	ad33;
5186	:douta	=	16'h	c5d4;
5187	:douta	=	16'h	5aed;
5188	:douta	=	16'h	5aeb;
5189	:douta	=	16'h	6b8e;
5190	:douta	=	16'h	bdd5;
5191	:douta	=	16'h	73af;
5192	:douta	=	16'h	bdd5;
5193	:douta	=	16'h	b555;
5194	:douta	=	16'h	deb9;
5195	:douta	=	16'h	6c34;
5196	:douta	=	16'h	bdb6;
5197	:douta	=	16'h	5bb2;
5198	:douta	=	16'h	8493;
5199	:douta	=	16'h	84d5;
5200	:douta	=	16'h	6390;
5201	:douta	=	16'h	c637;
5202	:douta	=	16'h	9d56;
5203	:douta	=	16'h	e71a;
5204	:douta	=	16'h	a4f5;
5205	:douta	=	16'h	d6ba;
5206	:douta	=	16'h	3b11;
5207	:douta	=	16'h	5373;
5208	:douta	=	16'h	8517;
5209	:douta	=	16'h	3a90;
5210	:douta	=	16'h	9db9;
5211	:douta	=	16'h	6c56;
5212	:douta	=	16'h	ce7b;
5213	:douta	=	16'h	6c77;
5214	:douta	=	16'h	7c75;
5215	:douta	=	16'h	4b73;
5216	:douta	=	16'h	9d37;
5217	:douta	=	16'h	be7b;
5218	:douta	=	16'h	222d;
5219	:douta	=	16'h	42d0;
5220	:douta	=	16'h	7455;
5221	:douta	=	16'h	5bd4;
5222	:douta	=	16'h	7455;
5223	:douta	=	16'h	a61b;
5224	:douta	=	16'h	6c98;
5225	:douta	=	16'h	84f7;
5226	:douta	=	16'h	8d19;
5227	:douta	=	16'h	9d99;
5228	:douta	=	16'h	222f;
5229	:douta	=	16'h	5bb3;
5230	:douta	=	16'h	7cd7;
5231	:douta	=	16'h	42f0;
5232	:douta	=	16'h	7476;
5233	:douta	=	16'h	5bb4;
5234	:douta	=	16'h	94d6;
5235	:douta	=	16'h	9d77;
5236	:douta	=	16'h	a558;
5237	:douta	=	16'h	8d37;
5238	:douta	=	16'h	73f2;
5239	:douta	=	16'h	c5f7;
5240	:douta	=	16'h	3a2c;
5241	:douta	=	16'h	42f0;
5242	:douta	=	16'h	320d;
5243	:douta	=	16'h	326d;
5244	:douta	=	16'h	6bf2;
5245	:douta	=	16'h	7c12;
5246	:douta	=	16'h	9d56;
5247	:douta	=	16'h	6c13;
5248	:douta	=	16'h	d679;
5249	:douta	=	16'h	b5d8;
5250	:douta	=	16'h	8494;
5251	:douta	=	16'h	6c14;
5252	:douta	=	16'h	5330;
5253	:douta	=	16'h	add8;
5254	:douta	=	16'h	8cd5;
5255	:douta	=	16'h	9537;
5256	:douta	=	16'h	4b2f;
5257	:douta	=	16'h	8453;
5258	:douta	=	16'h	4acf;
5259	:douta	=	16'h	31ca;
5260	:douta	=	16'h	5b71;
5261	:douta	=	16'h	7434;
5262	:douta	=	16'h	9d15;
5263	:douta	=	16'h	8431;
5264	:douta	=	16'h	2925;
5265	:douta	=	16'h	10e3;
5266	:douta	=	16'h	18e4;
5267	:douta	=	16'h	426b;
5268	:douta	=	16'h	638f;
5269	:douta	=	16'h	534e;
5270	:douta	=	16'h	2167;
5271	:douta	=	16'h	0042;
5272	:douta	=	16'h	10a4;
5273	:douta	=	16'h	18e5;
5274	:douta	=	16'h	10a5;
5275	:douta	=	16'h	10e5;
5276	:douta	=	16'h	10e5;
5277	:douta	=	16'h	10e5;
5278	:douta	=	16'h	10c4;
5279	:douta	=	16'h	0884;
5280	:douta	=	16'h	0843;
5281	:douta	=	16'h	2126;
5282	:douta	=	16'h	2988;
5283	:douta	=	16'h	39eb;
5284	:douta	=	16'h	426c;
5285	:douta	=	16'h	5aef;
5286	:douta	=	16'h	5310;
5287	:douta	=	16'h	5332;
5288	:douta	=	16'h	63d4;
5289	:douta	=	16'h	7476;
5290	:douta	=	16'h	6c15;
5291	:douta	=	16'h	63d4;
5292	:douta	=	16'h	74d9;
5293	:douta	=	16'h	6c79;
5294	:douta	=	16'h	74fa;
5295	:douta	=	16'h	7d1b;
5296	:douta	=	16'h	74b9;
5297	:douta	=	16'h	6c78;
5298	:douta	=	16'h	5c37;
5299	:douta	=	16'h	6c98;
5300	:douta	=	16'h	6c78;
5301	:douta	=	16'h	6457;
5302	:douta	=	16'h	6cb9;
5303	:douta	=	16'h	6457;
5304	:douta	=	16'h	6c77;
5305	:douta	=	16'h	7cf9;
5306	:douta	=	16'h	8d5b;
5307	:douta	=	16'h	7d1a;
5308	:douta	=	16'h	7d1a;
5309	:douta	=	16'h	7d3a;
5310	:douta	=	16'h	5bf6;
5311	:douta	=	16'h	6437;
5312	:douta	=	16'h	6cb9;
5313	:douta	=	16'h	6498;
5314	:douta	=	16'h	753b;
5315	:douta	=	16'h	7cfa;
5316	:douta	=	16'h	74f9;
5317	:douta	=	16'h	6415;
5318	:douta	=	16'h	6c56;
5319	:douta	=	16'h	4b52;
5320	:douta	=	16'h	5bb4;
5321	:douta	=	16'h	5bb4;
5322	:douta	=	16'h	4310;
5323	:douta	=	16'h	3a4c;
5324	:douta	=	16'h	29ca;
5325	:douta	=	16'h	2168;
5326	:douta	=	16'h	2147;
5327	:douta	=	16'h	0042;
5328	:douta	=	16'h	0062;
5329	:douta	=	16'h	0883;
5330	:douta	=	16'h	1084;
5331	:douta	=	16'h	08c4;
5332	:douta	=	16'h	08a4;
5333	:douta	=	16'h	08a4;
5334	:douta	=	16'h	10a4;
5335	:douta	=	16'h	0002;
5336	:douta	=	16'h	0001;
5337	:douta	=	16'h	1968;
5338	:douta	=	16'h	3af0;
5339	:douta	=	16'h	6c54;
5340	:douta	=	16'h	9d99;
5341	:douta	=	16'h	9d58;
5342	:douta	=	16'h	63f5;
5343	:douta	=	16'h	8473;
5344	:douta	=	16'h	7c76;
5345	:douta	=	16'h	220d;
5346	:douta	=	16'h	0149;
5347	:douta	=	16'h	328f;
5348	:douta	=	16'h	5b92;
5349	:douta	=	16'h	7c74;
5350	:douta	=	16'h	8cb5;
5351	:douta	=	16'h	4b11;
5352	:douta	=	16'h	a557;
5353	:douta	=	16'h	4b51;
5354	:douta	=	16'h	4b31;
5355	:douta	=	16'h	21ab;
5356	:douta	=	16'h	21aa;
5357	:douta	=	16'h	4b52;
5358	:douta	=	16'h	6c14;
5359	:douta	=	16'h	8cf6;
5360	:douta	=	16'h	7477;
5361	:douta	=	16'h	63f4;
5362	:douta	=	16'h	3af1;
5363	:douta	=	16'h	3ad1;
5364	:douta	=	16'h	4352;
5365	:douta	=	16'h	53b4;
5366	:douta	=	16'h	9d9a;
5367	:douta	=	16'h	6cb8;
5368	:douta	=	16'h	9e1d;
5369	:douta	=	16'h	4bf7;
5370	:douta	=	16'h	74fa;
5371	:douta	=	16'h	4b96;
5372	:douta	=	16'h	4375;
5373	:douta	=	16'h	1a0e;
5374	:douta	=	16'h	4374;
5375	:douta	=	16'h	74b8;
5376	:douta	=	16'h	3b33;
5377	:douta	=	16'h	4b74;
5378	:douta	=	16'h	6c37;
5379	:douta	=	16'h	6436;
5380	:douta	=	16'h	6c77;
5381	:douta	=	16'h	6c98;
5382	:douta	=	16'h	42b0;
5383	:douta	=	16'h	8498;
5384	:douta	=	16'h	5b93;
5385	:douta	=	16'h	7477;
5386	:douta	=	16'h	5b93;
5387	:douta	=	16'h	6b91;
5388	:douta	=	16'h	8cd6;
5389	:douta	=	16'h	8434;
5390	:douta	=	16'h	6b91;
5391	:douta	=	16'h	bdf8;
5392	:douta	=	16'h	8cd6;
5393	:douta	=	16'h	9d37;
5394	:douta	=	16'h	6c16;
5395	:douta	=	16'h	4aac;
5396	:douta	=	16'h	5b50;
5397	:douta	=	16'h	6391;
5398	:douta	=	16'h	6bd2;
5399	:douta	=	16'h	c618;
5400	:douta	=	16'h	c5d7;
5401	:douta	=	16'h	eefa;
5402	:douta	=	16'h	c5d7;
5403	:douta	=	16'h	deba;
5404	:douta	=	16'h	9d16;
5405	:douta	=	16'h	5b92;
5406	:douta	=	16'h	94d5;
5407	:douta	=	16'h	4b72;
5408	:douta	=	16'h	6330;
5409	:douta	=	16'h	a556;
5410	:douta	=	16'h	d678;
5411	:douta	=	16'h	bdd8;
5412	:douta	=	16'h	d699;
5413	:douta	=	16'h	ad55;
5414	:douta	=	16'h	b619;
5415	:douta	=	16'h	acd3;
5416	:douta	=	16'h	add7;
5417	:douta	=	16'h	b575;
5418	:douta	=	16'h	ad75;
5419	:douta	=	16'h	d658;
5420	:douta	=	16'h	ff9b;
5421	:douta	=	16'h	c618;
5422	:douta	=	16'h	83af;
5423	:douta	=	16'h	ce37;
5424	:douta	=	16'h	636e;
5425	:douta	=	16'h	6b90;
5426	:douta	=	16'h	7bef;
5427	:douta	=	16'h	ded9;
5428	:douta	=	16'h	c5d5;
5429	:douta	=	16'h	eef9;
5430	:douta	=	16'h	3a8f;
5431	:douta	=	16'h	6b2e;
5432	:douta	=	16'h	b5f5;
5433	:douta	=	16'h	9451;
5434	:douta	=	16'h	ad12;
5435	:douta	=	16'h	bd73;
5436	:douta	=	16'h	f75a;
5437	:douta	=	16'h	6baf;
5438	:douta	=	16'h	acd2;
5439	:douta	=	16'h	5b6f;
5440	:douta	=	16'h	9c91;
5441	:douta	=	16'h	c636;
5442	:douta	=	16'h	ce15;
5443	:douta	=	16'h	ad32;
5444	:douta	=	16'h	ce15;
5445	:douta	=	16'h	de57;
5446	:douta	=	16'h	c637;
5447	:douta	=	16'h	62ed;
5448	:douta	=	16'h	c5f7;
5449	:douta	=	16'h	42ae;
5450	:douta	=	16'h	8431;
5451	:douta	=	16'h	8432;
5452	:douta	=	16'h	c658;
5453	:douta	=	16'h	9d15;
5454	:douta	=	16'h	c5d6;
5455	:douta	=	16'h	5bf4;
5456	:douta	=	16'h	a4b4;
5457	:douta	=	16'h	5392;
5458	:douta	=	16'h	4b51;
5459	:douta	=	16'h	632f;
5460	:douta	=	16'h	8c72;
5461	:douta	=	16'h	c679;
5462	:douta	=	16'h	7454;
5463	:douta	=	16'h	ad97;
5464	:douta	=	16'h	7d18;
5465	:douta	=	16'h	5bb4;
5466	:douta	=	16'h	9dfb;
5467	:douta	=	16'h	5b92;
5468	:douta	=	16'h	84d6;
5469	:douta	=	16'h	322e;
5470	:douta	=	16'h	8495;
5471	:douta	=	16'h	5394;
5472	:douta	=	16'h	be3a;
5473	:douta	=	16'h	8d38;
5474	:douta	=	16'h	6bf5;
5475	:douta	=	16'h	8d38;
5476	:douta	=	16'h	7476;
5477	:douta	=	16'h	8d18;
5478	:douta	=	16'h	6c36;
5479	:douta	=	16'h	6c76;
5480	:douta	=	16'h	2a4f;
5481	:douta	=	16'h	7cb8;
5482	:douta	=	16'h	6c76;
5483	:douta	=	16'h	7476;
5484	:douta	=	16'h	7477;
5485	:douta	=	16'h	8518;
5486	:douta	=	16'h	8539;
5487	:douta	=	16'h	c6de;
5488	:douta	=	16'h	6457;
5489	:douta	=	16'h	73f3;
5490	:douta	=	16'h	6bd2;
5491	:douta	=	16'h	4b31;
5492	:douta	=	16'h	5330;
5493	:douta	=	16'h	21aa;
5494	:douta	=	16'h	8454;
5495	:douta	=	16'h	a555;
5496	:douta	=	16'h	7c95;
5497	:douta	=	16'h	7c95;
5498	:douta	=	16'h	7455;
5499	:douta	=	16'h	8474;
5500	:douta	=	16'h	deba;
5501	:douta	=	16'h	a536;
5502	:douta	=	16'h	5b72;
5503	:douta	=	16'h	428d;
5504	:douta	=	16'h	7c32;
5505	:douta	=	16'h	8454;
5506	:douta	=	16'h	7c54;
5507	:douta	=	16'h	63f3;
5508	:douta	=	16'h	bdd8;
5509	:douta	=	16'h	6bf2;
5510	:douta	=	16'h	7bf1;
5511	:douta	=	16'h	324e;
5512	:douta	=	16'h	94b6;
5513	:douta	=	16'h	9517;
5514	:douta	=	16'h	9cd6;
5515	:douta	=	16'h	c69a;
5516	:douta	=	16'h	7435;
5517	:douta	=	16'h	9cd4;
5518	:douta	=	16'h	7c12;
5519	:douta	=	16'h	8454;
5520	:douta	=	16'h	528c;
5521	:douta	=	16'h	1905;
5522	:douta	=	16'h	2966;
5523	:douta	=	16'h	2167;
5524	:douta	=	16'h	0883;
5525	:douta	=	16'h	18e4;
5526	:douta	=	16'h	18e5;
5527	:douta	=	16'h	10c5;
5528	:douta	=	16'h	18e5;
5529	:douta	=	16'h	18e5;
5530	:douta	=	16'h	10e4;
5531	:douta	=	16'h	0863;
5532	:douta	=	16'h	18e4;
5533	:douta	=	16'h	3147;
5534	:douta	=	16'h	4a4b;
5535	:douta	=	16'h	5aee;
5536	:douta	=	16'h	73d3;
5537	:douta	=	16'h	5351;
5538	:douta	=	16'h	5373;
5539	:douta	=	16'h	7499;
5540	:douta	=	16'h	7499;
5541	:douta	=	16'h	855a;
5542	:douta	=	16'h	7d19;
5543	:douta	=	16'h	74d9;
5544	:douta	=	16'h	74da;
5545	:douta	=	16'h	74d9;
5546	:douta	=	16'h	6cb9;
5547	:douta	=	16'h	6457;
5548	:douta	=	16'h	6cba;
5549	:douta	=	16'h	7d3a;
5550	:douta	=	16'h	74d9;
5551	:douta	=	16'h	6cb8;
5552	:douta	=	16'h	74f9;
5553	:douta	=	16'h	74fa;
5554	:douta	=	16'h	74d9;
5555	:douta	=	16'h	855a;
5556	:douta	=	16'h	7cfa;
5557	:douta	=	16'h	7cda;
5558	:douta	=	16'h	7498;
5559	:douta	=	16'h	7d3a;
5560	:douta	=	16'h	74d9;
5561	:douta	=	16'h	6c77;
5562	:douta	=	16'h	6c77;
5563	:douta	=	16'h	74d9;
5564	:douta	=	16'h	74d9;
5565	:douta	=	16'h	6c98;
5566	:douta	=	16'h	855c;
5567	:douta	=	16'h	855c;
5568	:douta	=	16'h	6cd9;
5569	:douta	=	16'h	7d3b;
5570	:douta	=	16'h	74da;
5571	:douta	=	16'h	74b8;
5572	:douta	=	16'h	855a;
5573	:douta	=	16'h	6cd9;
5574	:douta	=	16'h	7d1a;
5575	:douta	=	16'h	74fa;
5576	:douta	=	16'h	6c98;
5577	:douta	=	16'h	5c37;
5578	:douta	=	16'h	6458;
5579	:douta	=	16'h	7d5b;
5580	:douta	=	16'h	7d3b;
5581	:douta	=	16'h	6416;
5582	:douta	=	16'h	5b93;
5583	:douta	=	16'h	42af;
5584	:douta	=	16'h	42af;
5585	:douta	=	16'h	322c;
5586	:douta	=	16'h	29a9;
5587	:douta	=	16'h	10e5;
5588	:douta	=	16'h	0042;
5589	:douta	=	16'h	0883;
5590	:douta	=	16'h	08c4;
5591	:douta	=	16'h	10a4;
5592	:douta	=	16'h	08a5;
5593	:douta	=	16'h	08a4;
5594	:douta	=	16'h	08a4;
5595	:douta	=	16'h	0043;
5596	:douta	=	16'h	0927;
5597	:douta	=	16'h	11aa;
5598	:douta	=	16'h	7c96;
5599	:douta	=	16'h	7c54;
5600	:douta	=	16'h	7414;
5601	:douta	=	16'h	8cb6;
5602	:douta	=	16'h	6bf4;
5603	:douta	=	16'h	5330;
5604	:douta	=	16'h	32af;
5605	:douta	=	16'h	2a4d;
5606	:douta	=	16'h	3acf;
5607	:douta	=	16'h	7c75;
5608	:douta	=	16'h	9d16;
5609	:douta	=	16'h	9516;
5610	:douta	=	16'h	a557;
5611	:douta	=	16'h	42f0;
5612	:douta	=	16'h	4b31;
5613	:douta	=	16'h	2a6f;
5614	:douta	=	16'h	220e;
5615	:douta	=	16'h	2a6f;
5616	:douta	=	16'h	3b32;
5617	:douta	=	16'h	53d3;
5618	:douta	=	16'h	6c35;
5619	:douta	=	16'h	4b95;
5620	:douta	=	16'h	4b94;
5621	:douta	=	16'h	7499;
5622	:douta	=	16'h	3b33;
5623	:douta	=	16'h	4bb6;
5624	:douta	=	16'h	3b54;
5625	:douta	=	16'h	7cf9;
5626	:douta	=	16'h	8d3b;
5627	:douta	=	16'h	959c;
5628	:douta	=	16'h	6457;
5629	:douta	=	16'h	7d7b;
5630	:douta	=	16'h	5c38;
5631	:douta	=	16'h	7c77;
5632	:douta	=	16'h	74fa;
5633	:douta	=	16'h	4333;
5634	:douta	=	16'h	6c78;
5635	:douta	=	16'h	7d1a;
5636	:douta	=	16'h	4b95;
5637	:douta	=	16'h	4b53;
5638	:douta	=	16'h	5bb4;
5639	:douta	=	16'h	5331;
5640	:douta	=	16'h	63b3;
5641	:douta	=	16'h	8519;
5642	:douta	=	16'h	7456;
5643	:douta	=	16'h	6371;
5644	:douta	=	16'h	5b72;
5645	:douta	=	16'h	5330;
5646	:douta	=	16'h	42ae;
5647	:douta	=	16'h	7c34;
5648	:douta	=	16'h	b5b8;
5649	:douta	=	16'h	de99;
5650	:douta	=	16'h	9538;
5651	:douta	=	16'h	b576;
5652	:douta	=	16'h	a577;
5653	:douta	=	16'h	530f;
5654	:douta	=	16'h	8454;
5655	:douta	=	16'h	5b0f;
5656	:douta	=	16'h	7bf2;
5657	:douta	=	16'h	9cf4;
5658	:douta	=	16'h	b597;
5659	:douta	=	16'h	9d56;
5660	:douta	=	16'h	b5d8;
5661	:douta	=	16'h	cebb;
5662	:douta	=	16'h	bdd8;
5663	:douta	=	16'h	8c95;
5664	:douta	=	16'h	bd76;
5665	:douta	=	16'h	94b5;
5666	:douta	=	16'h	a576;
5667	:douta	=	16'h	7c53;
5668	:douta	=	16'h	bdb7;
5669	:douta	=	16'h	eefa;
5670	:douta	=	16'h	d6ba;
5671	:douta	=	16'h	e657;
5672	:douta	=	16'h	b65a;
5673	:douta	=	16'h	9473;
5674	:douta	=	16'h	7c53;
5675	:douta	=	16'h	8432;
5676	:douta	=	16'h	c616;
5677	:douta	=	16'h	d637;
5678	:douta	=	16'h	d617;
5679	:douta	=	16'h	d698;
5680	:douta	=	16'h	ad34;
5681	:douta	=	16'h	7412;
5682	:douta	=	16'h	3a8d;
5683	:douta	=	16'h	c616;
5684	:douta	=	16'h	a514;
5685	:douta	=	16'h	f759;
5686	:douta	=	16'h	ad33;
5687	:douta	=	16'h	de57;
5688	:douta	=	16'h	6bcf;
5689	:douta	=	16'h	3a0a;
5690	:douta	=	16'h	6bf0;
5691	:douta	=	16'h	b512;
5692	:douta	=	16'h	bdd4;
5693	:douta	=	16'h	ad12;
5694	:douta	=	16'h	de57;
5695	:douta	=	16'h	8c71;
5696	:douta	=	16'h	ce57;
5697	:douta	=	16'h	a513;
5698	:douta	=	16'h	9491;
5699	:douta	=	16'h	8c71;
5700	:douta	=	16'h	6b4b;
5701	:douta	=	16'h	ef39;
5702	:douta	=	16'h	ce76;
5703	:douta	=	16'h	9c0f;
5704	:douta	=	16'h	e6d7;
5705	:douta	=	16'h	5b2f;
5706	:douta	=	16'h	a576;
5707	:douta	=	16'h	6bb1;
5708	:douta	=	16'h	6bd1;
5709	:douta	=	16'h	7bf2;
5710	:douta	=	16'h	d637;
5711	:douta	=	16'h	6413;
5712	:douta	=	16'h	8c52;
5713	:douta	=	16'h	7495;
5714	:douta	=	16'h	5372;
5715	:douta	=	16'h	deba;
5716	:douta	=	16'h	52cd;
5717	:douta	=	16'h	a557;
5718	:douta	=	16'h	3acf;
5719	:douta	=	16'h	9d16;
5720	:douta	=	16'h	5bb2;
5721	:douta	=	16'h	8c53;
5722	:douta	=	16'h	ae3b;
5723	:douta	=	16'h	9cd7;
5724	:douta	=	16'h	d6dc;
5725	:douta	=	16'h	42f1;
5726	:douta	=	16'h	ad98;
5727	:douta	=	16'h	220e;
5728	:douta	=	16'h	7c34;
5729	:douta	=	16'h	8d38;
5730	:douta	=	16'h	5c15;
5731	:douta	=	16'h	32d2;
5732	:douta	=	16'h	8d38;
5733	:douta	=	16'h	7497;
5734	:douta	=	16'h	9518;
5735	:douta	=	16'h	859b;
5736	:douta	=	16'h	4bf6;
5737	:douta	=	16'h	8cb6;
5738	:douta	=	16'h	6c56;
5739	:douta	=	16'h	5bb4;
5740	:douta	=	16'h	84b8;
5741	:douta	=	16'h	9559;
5742	:douta	=	16'h	5415;
5743	:douta	=	16'h	6c76;
5744	:douta	=	16'h	5bf5;
5745	:douta	=	16'h	8cb5;
5746	:douta	=	16'h	94f6;
5747	:douta	=	16'h	5b92;
5748	:douta	=	16'h	6c76;
5749	:douta	=	16'h	7414;
5750	:douta	=	16'h	632f;
5751	:douta	=	16'h	9d15;
5752	:douta	=	16'h	3a4d;
5753	:douta	=	16'h	322c;
5754	:douta	=	16'h	5351;
5755	:douta	=	16'h	6bd2;
5756	:douta	=	16'h	6c13;
5757	:douta	=	16'h	a577;
5758	:douta	=	16'h	7434;
5759	:douta	=	16'h	8cf6;
5760	:douta	=	16'h	9d57;
5761	:douta	=	16'h	84b5;
5762	:douta	=	16'h	a577;
5763	:douta	=	16'h	324e;
5764	:douta	=	16'h	63b2;
5765	:douta	=	16'h	8c94;
5766	:douta	=	16'h	c618;
5767	:douta	=	16'h	7454;
5768	:douta	=	16'h	9d17;
5769	:douta	=	16'h	9559;
5770	:douta	=	16'h	7413;
5771	:douta	=	16'h	84d7;
5772	:douta	=	16'h	6c14;
5773	:douta	=	16'h	a598;
5774	:douta	=	16'h	9536;
5775	:douta	=	16'h	bdf9;
5776	:douta	=	16'h	63b1;
5777	:douta	=	16'h	2987;
5778	:douta	=	16'h	2125;
5779	:douta	=	16'h	18e5;
5780	:douta	=	16'h	18e5;
5781	:douta	=	16'h	18e5;
5782	:douta	=	16'h	10e5;
5783	:douta	=	16'h	18e5;
5784	:douta	=	16'h	10e4;
5785	:douta	=	16'h	0863;
5786	:douta	=	16'h	10a3;
5787	:douta	=	16'h	31a8;
5788	:douta	=	16'h	5acd;
5789	:douta	=	16'h	6b4f;
5790	:douta	=	16'h	7414;
5791	:douta	=	16'h	7414;
5792	:douta	=	16'h	84f9;
5793	:douta	=	16'h	955b;
5794	:douta	=	16'h	74d9;
5795	:douta	=	16'h	6457;
5796	:douta	=	16'h	74f9;
5797	:douta	=	16'h	7d1a;
5798	:douta	=	16'h	853a;
5799	:douta	=	16'h	7d1a;
5800	:douta	=	16'h	6cb9;
5801	:douta	=	16'h	7d1a;
5802	:douta	=	16'h	6cb9;
5803	:douta	=	16'h	74d9;
5804	:douta	=	16'h	4bf7;
5805	:douta	=	16'h	6c79;
5806	:douta	=	16'h	6478;
5807	:douta	=	16'h	6c78;
5808	:douta	=	16'h	6437;
5809	:douta	=	16'h	7d1a;
5810	:douta	=	16'h	7cfa;
5811	:douta	=	16'h	74b9;
5812	:douta	=	16'h	5c16;
5813	:douta	=	16'h	6436;
5814	:douta	=	16'h	7499;
5815	:douta	=	16'h	7d1a;
5816	:douta	=	16'h	7cf9;
5817	:douta	=	16'h	7cf9;
5818	:douta	=	16'h	7cd9;
5819	:douta	=	16'h	6c57;
5820	:douta	=	16'h	6c78;
5821	:douta	=	16'h	6c78;
5822	:douta	=	16'h	6cb9;
5823	:douta	=	16'h	74da;
5824	:douta	=	16'h	855b;
5825	:douta	=	16'h	6478;
5826	:douta	=	16'h	7d3b;
5827	:douta	=	16'h	6cb9;
5828	:douta	=	16'h	6cb9;
5829	:douta	=	16'h	6478;
5830	:douta	=	16'h	855c;
5831	:douta	=	16'h	857b;
5832	:douta	=	16'h	74da;
5833	:douta	=	16'h	74da;
5834	:douta	=	16'h	6cb8;
5835	:douta	=	16'h	751a;
5836	:douta	=	16'h	74da;
5837	:douta	=	16'h	7d5b;
5838	:douta	=	16'h	857c;
5839	:douta	=	16'h	6436;
5840	:douta	=	16'h	5bf5;
5841	:douta	=	16'h	5351;
5842	:douta	=	16'h	42d0;
5843	:douta	=	16'h	42af;
5844	:douta	=	16'h	2989;
5845	:douta	=	16'h	0884;
5846	:douta	=	16'h	0062;
5847	:douta	=	16'h	08a4;
5848	:douta	=	16'h	10a4;
5849	:douta	=	16'h	10c5;
5850	:douta	=	16'h	08a4;
5851	:douta	=	16'h	10c4;
5852	:douta	=	16'h	0863;
5853	:douta	=	16'h	0064;
5854	:douta	=	16'h	32af;
5855	:douta	=	16'h	5b92;
5856	:douta	=	16'h	7cb5;
5857	:douta	=	16'h	8c75;
5858	:douta	=	16'h	8454;
5859	:douta	=	16'h	6bb2;
5860	:douta	=	16'h	7413;
5861	:douta	=	16'h	7c34;
5862	:douta	=	16'h	328e;
5863	:douta	=	16'h	3acf;
5864	:douta	=	16'h	3acf;
5865	:douta	=	16'h	7c54;
5866	:douta	=	16'h	7c94;
5867	:douta	=	16'h	6bf2;
5868	:douta	=	16'h	94b5;
5869	:douta	=	16'h	5b92;
5870	:douta	=	16'h	53b4;
5871	:douta	=	16'h	21ec;
5872	:douta	=	16'h	4b32;
5873	:douta	=	16'h	222e;
5874	:douta	=	16'h	6c35;
5875	:douta	=	16'h	3ad1;
5876	:douta	=	16'h	53b4;
5877	:douta	=	16'h	959b;
5878	:douta	=	16'h	957a;
5879	:douta	=	16'h	4375;
5880	:douta	=	16'h	4bb5;
5881	:douta	=	16'h	4b95;
5882	:douta	=	16'h	3b33;
5883	:douta	=	16'h	5bf5;
5884	:douta	=	16'h	5416;
5885	:douta	=	16'h	5c37;
5886	:douta	=	16'h	5bb3;
5887	:douta	=	16'h	8519;
5888	:douta	=	16'h	4374;
5889	:douta	=	16'h	224f;
5890	:douta	=	16'h	32b0;
5891	:douta	=	16'h	6416;
5892	:douta	=	16'h	6437;
5893	:douta	=	16'h	6c78;
5894	:douta	=	16'h	63d4;
5895	:douta	=	16'h	42cf;
5896	:douta	=	16'h	6436;
5897	:douta	=	16'h	5372;
5898	:douta	=	16'h	4b52;
5899	:douta	=	16'h	6371;
5900	:douta	=	16'h	94f6;
5901	:douta	=	16'h	8454;
5902	:douta	=	16'h	8cf7;
5903	:douta	=	16'h	8c74;
5904	:douta	=	16'h	a579;
5905	:douta	=	16'h	8495;
5906	:douta	=	16'h	84d8;
5907	:douta	=	16'h	a536;
5908	:douta	=	16'h	5b50;
5909	:douta	=	16'h	ce17;
5910	:douta	=	16'h	ad56;
5911	:douta	=	16'h	d658;
5912	:douta	=	16'h	ce79;
5913	:douta	=	16'h	9d15;
5914	:douta	=	16'h	bdf8;
5915	:douta	=	16'h	6c34;
5916	:douta	=	16'h	73d1;
5917	:douta	=	16'h	8433;
5918	:douta	=	16'h	ad36;
5919	:douta	=	16'h	7433;
5920	:douta	=	16'h	9d15;
5921	:douta	=	16'h	adb7;
5922	:douta	=	16'h	ce58;
5923	:douta	=	16'h	ef3a;
5924	:douta	=	16'h	a535;
5925	:douta	=	16'h	8c72;
5926	:douta	=	16'h	9d36;
5927	:douta	=	16'h	d678;
5928	:douta	=	16'h	d678;
5929	:douta	=	16'h	a514;
5930	:douta	=	16'h	e698;
5931	:douta	=	16'h	d698;
5932	:douta	=	16'h	ef3a;
5933	:douta	=	16'h	a515;
5934	:douta	=	16'h	a4b3;
5935	:douta	=	16'h	ce37;
5936	:douta	=	16'h	8411;
5937	:douta	=	16'h	a514;
5938	:douta	=	16'h	9c91;
5939	:douta	=	16'h	ef5a;
5940	:douta	=	16'h	b595;
5941	:douta	=	16'h	ce16;
5942	:douta	=	16'h	632d;
5943	:douta	=	16'h	83ae;
5944	:douta	=	16'h	a511;
5945	:douta	=	16'h	ad12;
5946	:douta	=	16'h	9470;
5947	:douta	=	16'h	e6b8;
5948	:douta	=	16'h	de77;
5949	:douta	=	16'h	632d;
5950	:douta	=	16'h	6b2c;
5951	:douta	=	16'h	4aad;
5952	:douta	=	16'h	d676;
5953	:douta	=	16'h	ce15;
5954	:douta	=	16'h	e6d7;
5955	:douta	=	16'h	c5d4;
5956	:douta	=	16'h	acf2;
5957	:douta	=	16'h	a512;
5958	:douta	=	16'h	532d;
5959	:douta	=	16'h	9450;
5960	:douta	=	16'h	7c51;
5961	:douta	=	16'h	94b2;
5962	:douta	=	16'h	9d55;
5963	:douta	=	16'h	8431;
5964	:douta	=	16'h	b5d7;
5965	:douta	=	16'h	6bf2;
5966	:douta	=	16'h	b5d7;
5967	:douta	=	16'h	5b50;
5968	:douta	=	16'h	7c74;
5969	:douta	=	16'h	428d;
5970	:douta	=	16'h	73f1;
5971	:douta	=	16'h	ad96;
5972	:douta	=	16'h	c638;
5973	:douta	=	16'h	9d76;
5974	:douta	=	16'h	9d36;
5975	:douta	=	16'h	c658;
5976	:douta	=	16'h	8476;
5977	:douta	=	16'h	d699;
5978	:douta	=	16'h	4353;
5979	:douta	=	16'h	6bd3;
5980	:douta	=	16'h	7433;
5981	:douta	=	16'h	7434;
5982	:douta	=	16'h	8cf6;
5983	:douta	=	16'h	6477;
5984	:douta	=	16'h	be39;
5985	:douta	=	16'h	8d5a;
5986	:douta	=	16'h	5bb2;
5987	:douta	=	16'h	5c15;
5988	:douta	=	16'h	4311;
5989	:douta	=	16'h	4b51;
5990	:douta	=	16'h	4332;
5991	:douta	=	16'h	4b73;
5992	:douta	=	16'h	6c98;
5993	:douta	=	16'h	6414;
5994	:douta	=	16'h	7c96;
5995	:douta	=	16'h	855a;
5996	:douta	=	16'h	7cd8;
5997	:douta	=	16'h	a5b9;
5998	:douta	=	16'h	6436;
5999	:douta	=	16'h	53d4;
6000	:douta	=	16'h	32b1;
6001	:douta	=	16'h	b5f8;
6002	:douta	=	16'h	a5b9;
6003	:douta	=	16'h	3aaf;
6004	:douta	=	16'h	4b31;
6005	:douta	=	16'h	6c76;
6006	:douta	=	16'h	a535;
6007	:douta	=	16'h	be59;
6008	:douta	=	16'h	8517;
6009	:douta	=	16'h	63f4;
6010	:douta	=	16'h	84d7;
6011	:douta	=	16'h	be3a;
6012	:douta	=	16'h	6bf4;
6013	:douta	=	16'h	b5b7;
6014	:douta	=	16'h	5371;
6015	:douta	=	16'h	4aad;
6016	:douta	=	16'h	3a4c;
6017	:douta	=	16'h	7c33;
6018	:douta	=	16'h	5392;
6019	:douta	=	16'h	7c96;
6020	:douta	=	16'h	9515;
6021	:douta	=	16'h	9473;
6022	:douta	=	16'h	9d56;
6023	:douta	=	16'h	3a4e;
6024	:douta	=	16'h	5bd3;
6025	:douta	=	16'h	21ed;
6026	:douta	=	16'h	b659;
6027	:douta	=	16'h	6c35;
6028	:douta	=	16'h	84f8;
6029	:douta	=	16'h	7496;
6030	:douta	=	16'h	8d37;
6031	:douta	=	16'h	1127;
6032	:douta	=	16'h	18e5;
6033	:douta	=	16'h	1906;
6034	:douta	=	16'h	2125;
6035	:douta	=	16'h	1905;
6036	:douta	=	16'h	1905;
6037	:douta	=	16'h	10c5;
6038	:douta	=	16'h	1083;
6039	:douta	=	16'h	39c8;
6040	:douta	=	16'h	422a;
6041	:douta	=	16'h	6b70;
6042	:douta	=	16'h	8434;
6043	:douta	=	16'h	7c55;
6044	:douta	=	16'h	7cd9;
6045	:douta	=	16'h	7cf9;
6046	:douta	=	16'h	853a;
6047	:douta	=	16'h	855a;
6048	:douta	=	16'h	7cd9;
6049	:douta	=	16'h	8d5b;
6050	:douta	=	16'h	9dbc;
6051	:douta	=	16'h	a61c;
6052	:douta	=	16'h	959b;
6053	:douta	=	16'h	7cda;
6054	:douta	=	16'h	74fa;
6055	:douta	=	16'h	74d9;
6056	:douta	=	16'h	74fa;
6057	:douta	=	16'h	74b9;
6058	:douta	=	16'h	6c57;
6059	:douta	=	16'h	6c98;
6060	:douta	=	16'h	855b;
6061	:douta	=	16'h	5c17;
6062	:douta	=	16'h	6479;
6063	:douta	=	16'h	6478;
6064	:douta	=	16'h	6478;
6065	:douta	=	16'h	7d3a;
6066	:douta	=	16'h	6457;
6067	:douta	=	16'h	6458;
6068	:douta	=	16'h	7d1a;
6069	:douta	=	16'h	7cfa;
6070	:douta	=	16'h	7499;
6071	:douta	=	16'h	6c98;
6072	:douta	=	16'h	74da;
6073	:douta	=	16'h	857b;
6074	:douta	=	16'h	7d3b;
6075	:douta	=	16'h	74d9;
6076	:douta	=	16'h	7d1a;
6077	:douta	=	16'h	855b;
6078	:douta	=	16'h	74d9;
6079	:douta	=	16'h	74d9;
6080	:douta	=	16'h	6c98;
6081	:douta	=	16'h	6cb9;
6082	:douta	=	16'h	74d9;
6083	:douta	=	16'h	8d9b;
6084	:douta	=	16'h	855b;
6085	:douta	=	16'h	74fa;
6086	:douta	=	16'h	751a;
6087	:douta	=	16'h	751a;
6088	:douta	=	16'h	7d1b;
6089	:douta	=	16'h	7d1b;
6090	:douta	=	16'h	6cb9;
6091	:douta	=	16'h	6498;
6092	:douta	=	16'h	6cb8;
6093	:douta	=	16'h	6478;
6094	:douta	=	16'h	6457;
6095	:douta	=	16'h	7d3b;
6096	:douta	=	16'h	751b;
6097	:douta	=	16'h	6cfa;
6098	:douta	=	16'h	755b;
6099	:douta	=	16'h	74fa;
6100	:douta	=	16'h	6c77;
6101	:douta	=	16'h	5331;
6102	:douta	=	16'h	42cf;
6103	:douta	=	16'h	29eb;
6104	:douta	=	16'h	2189;
6105	:douta	=	16'h	0863;
6106	:douta	=	16'h	08a4;
6107	:douta	=	16'h	10c5;
6108	:douta	=	16'h	10e5;
6109	:douta	=	16'h	10e5;
6110	:douta	=	16'h	08c4;
6111	:douta	=	16'h	0064;
6112	:douta	=	16'h	0907;
6113	:douta	=	16'h	63b2;
6114	:douta	=	16'h	6414;
6115	:douta	=	16'h	7c53;
6116	:douta	=	16'h	7c13;
6117	:douta	=	16'h	6bb2;
6118	:douta	=	16'h	9d16;
6119	:douta	=	16'h	8cb6;
6120	:douta	=	16'h	7c55;
6121	:douta	=	16'h	2a4d;
6122	:douta	=	16'h	1989;
6123	:douta	=	16'h	6bd3;
6124	:douta	=	16'h	42cf;
6125	:douta	=	16'h	ad77;
6126	:douta	=	16'h	3b12;
6127	:douta	=	16'h	5b72;
6128	:douta	=	16'h	3b33;
6129	:douta	=	16'h	4bb5;
6130	:douta	=	16'h	11cc;
6131	:douta	=	16'h	3ad0;
6132	:douta	=	16'h	4312;
6133	:douta	=	16'h	5bf5;
6134	:douta	=	16'h	7498;
6135	:douta	=	16'h	6c56;
6136	:douta	=	16'h	955a;
6137	:douta	=	16'h	53f6;
6138	:douta	=	16'h	53d5;
6139	:douta	=	16'h	53d5;
6140	:douta	=	16'h	3af2;
6141	:douta	=	16'h	2a2f;
6142	:douta	=	16'h	2a4e;
6143	:douta	=	16'h	53d4;
6144	:douta	=	16'h	5c37;
6145	:douta	=	16'h	53f6;
6146	:douta	=	16'h	42d1;
6147	:douta	=	16'h	6c77;
6148	:douta	=	16'h	3b33;
6149	:douta	=	16'h	3b12;
6150	:douta	=	16'h	6c36;
6151	:douta	=	16'h	7cb8;
6152	:douta	=	16'h	5b93;
6153	:douta	=	16'h	955a;
6154	:douta	=	16'h	953a;
6155	:douta	=	16'h	5310;
6156	:douta	=	16'h	6bd3;
6157	:douta	=	16'h	5b31;
6158	:douta	=	16'h	5b51;
6159	:douta	=	16'h	8454;
6160	:douta	=	16'h	94f6;
6161	:douta	=	16'h	a536;
6162	:douta	=	16'h	a5ba;
6163	:douta	=	16'h	8cb5;
6164	:douta	=	16'h	6391;
6165	:douta	=	16'h	73f1;
6166	:douta	=	16'h	6b90;
6167	:douta	=	16'h	8432;
6168	:douta	=	16'h	ad55;
6169	:douta	=	16'h	bdd7;
6170	:douta	=	16'h	e6da;
6171	:douta	=	16'h	add9;
6172	:douta	=	16'h	c5f9;
6173	:douta	=	16'h	bdd8;
6174	:douta	=	16'h	8494;
6175	:douta	=	16'h	a557;
6176	:douta	=	16'h	6392;
6177	:douta	=	16'h	8c94;
6178	:douta	=	16'h	94f5;
6179	:douta	=	16'h	94d3;
6180	:douta	=	16'h	d679;
6181	:douta	=	16'h	deb9;
6182	:douta	=	16'h	b5d8;
6183	:douta	=	16'h	d698;
6184	:douta	=	16'h	9d56;
6185	:douta	=	16'h	a4f3;
6186	:douta	=	16'h	8472;
6187	:douta	=	16'h	b595;
6188	:douta	=	16'h	d698;
6189	:douta	=	16'h	bd94;
6190	:douta	=	16'h	e6f9;
6191	:douta	=	16'h	de99;
6192	:douta	=	16'h	73f1;
6193	:douta	=	16'h	7c12;
6194	:douta	=	16'h	326c;
6195	:douta	=	16'h	bd94;
6196	:douta	=	16'h	bdb4;
6197	:douta	=	16'h	e719;
6198	:douta	=	16'h	cdd4;
6199	:douta	=	16'h	de77;
6200	:douta	=	16'h	5b0d;
6201	:douta	=	16'h	8410;
6202	:douta	=	16'h	52cd;
6203	:douta	=	16'h	c5d4;
6204	:douta	=	16'h	d657;
6205	:douta	=	16'h	9470;
6206	:douta	=	16'h	d616;
6207	:douta	=	16'h	632c;
6208	:douta	=	16'h	d697;
6209	:douta	=	16'h	ad54;
6210	:douta	=	16'h	8c4f;
6211	:douta	=	16'h	a512;
6212	:douta	=	16'h	a4f1;
6213	:douta	=	16'h	ce15;
6214	:douta	=	16'h	8431;
6215	:douta	=	16'h	c5d4;
6216	:douta	=	16'h	7c30;
6217	:douta	=	16'h	9cf3;
6218	:douta	=	16'h	530f;
6219	:douta	=	16'h	7b8e;
6220	:douta	=	16'h	9d34;
6221	:douta	=	16'h	8c73;
6222	:douta	=	16'h	e71a;
6223	:douta	=	16'h	73f2;
6224	:douta	=	16'h	9d16;
6225	:douta	=	16'h	4b0f;
6226	:douta	=	16'h	5b51;
6227	:douta	=	16'h	9d76;
6228	:douta	=	16'h	42ee;
6229	:douta	=	16'h	6bf2;
6230	:douta	=	16'h	7433;
6231	:douta	=	16'h	4b30;
6232	:douta	=	16'h	8cd6;
6233	:douta	=	16'h	be18;
6234	:douta	=	16'h	5bf5;
6235	:douta	=	16'h	94f6;
6236	:douta	=	16'h	a598;
6237	:douta	=	16'h	6c13;
6238	:douta	=	16'h	3aaf;
6239	:douta	=	16'h	5373;
6240	:douta	=	16'h	9517;
6241	:douta	=	16'h	6cd8;
6242	:douta	=	16'h	9579;
6243	:douta	=	16'h	6478;
6244	:douta	=	16'h	8496;
6245	:douta	=	16'h	6436;
6246	:douta	=	16'h	7c76;
6247	:douta	=	16'h	3312;
6248	:douta	=	16'h	4b94;
6249	:douta	=	16'h	42f1;
6250	:douta	=	16'h	63d5;
6251	:douta	=	16'h	3af1;
6252	:douta	=	16'h	95bb;
6253	:douta	=	16'h	9599;
6254	:douta	=	16'h	7497;
6255	:douta	=	16'h	7498;
6256	:douta	=	16'h	4b94;
6257	:douta	=	16'h	9d57;
6258	:douta	=	16'h	6c55;
6259	:douta	=	16'h	5b2f;
6260	:douta	=	16'h	220d;
6261	:douta	=	16'h	6c14;
6262	:douta	=	16'h	5351;
6263	:douta	=	16'h	5372;
6264	:douta	=	16'h	63b3;
6265	:douta	=	16'h	6414;
6266	:douta	=	16'h	6c14;
6267	:douta	=	16'h	7c96;
6268	:douta	=	16'h	5351;
6269	:douta	=	16'h	9557;
6270	:douta	=	16'h	7455;
6271	:douta	=	16'h	9d36;
6272	:douta	=	16'h	6bd3;
6273	:douta	=	16'h	9538;
6274	:douta	=	16'h	428f;
6275	:douta	=	16'h	428e;
6276	:douta	=	16'h	424b;
6277	:douta	=	16'h	add8;
6278	:douta	=	16'h	7cb5;
6279	:douta	=	16'h	84b6;
6280	:douta	=	16'h	84d7;
6281	:douta	=	16'h	4ad0;
6282	:douta	=	16'h	5bb3;
6283	:douta	=	16'h	21ec;
6284	:douta	=	16'h	7c54;
6285	:douta	=	16'h	5330;
6286	:douta	=	16'h	322b;
6287	:douta	=	16'h	18c4;
6288	:douta	=	16'h	2126;
6289	:douta	=	16'h	2126;
6290	:douta	=	16'h	2125;
6291	:douta	=	16'h	10e5;
6292	:douta	=	16'h	1083;
6293	:douta	=	16'h	2105;
6294	:douta	=	16'h	522a;
6295	:douta	=	16'h	5b0e;
6296	:douta	=	16'h	7c74;
6297	:douta	=	16'h	7434;
6298	:douta	=	16'h	7c98;
6299	:douta	=	16'h	851a;
6300	:douta	=	16'h	853a;
6301	:douta	=	16'h	851a;
6302	:douta	=	16'h	8519;
6303	:douta	=	16'h	8d5b;
6304	:douta	=	16'h	8519;
6305	:douta	=	16'h	7d3a;
6306	:douta	=	16'h	853b;
6307	:douta	=	16'h	959b;
6308	:douta	=	16'h	a5fc;
6309	:douta	=	16'h	95bb;
6310	:douta	=	16'h	853a;
6311	:douta	=	16'h	8d5b;
6312	:douta	=	16'h	74d9;
6313	:douta	=	16'h	74d9;
6314	:douta	=	16'h	6478;
6315	:douta	=	16'h	5c16;
6316	:douta	=	16'h	7cfa;
6317	:douta	=	16'h	74da;
6318	:douta	=	16'h	74da;
6319	:douta	=	16'h	6cba;
6320	:douta	=	16'h	74da;
6321	:douta	=	16'h	5c38;
6322	:douta	=	16'h	74f9;
6323	:douta	=	16'h	7cf9;
6324	:douta	=	16'h	6cb9;
6325	:douta	=	16'h	7cd9;
6326	:douta	=	16'h	74d9;
6327	:douta	=	16'h	6c99;
6328	:douta	=	16'h	6cb9;
6329	:douta	=	16'h	74d9;
6330	:douta	=	16'h	855b;
6331	:douta	=	16'h	7d5a;
6332	:douta	=	16'h	6cb9;
6333	:douta	=	16'h	74f9;
6334	:douta	=	16'h	857b;
6335	:douta	=	16'h	95bc;
6336	:douta	=	16'h	6437;
6337	:douta	=	16'h	6c98;
6338	:douta	=	16'h	74f9;
6339	:douta	=	16'h	7d3a;
6340	:douta	=	16'h	859b;
6341	:douta	=	16'h	857b;
6342	:douta	=	16'h	74fa;
6343	:douta	=	16'h	74fa;
6344	:douta	=	16'h	7d1a;
6345	:douta	=	16'h	857b;
6346	:douta	=	16'h	855b;
6347	:douta	=	16'h	74d9;
6348	:douta	=	16'h	6cb9;
6349	:douta	=	16'h	855b;
6350	:douta	=	16'h	7d1a;
6351	:douta	=	16'h	5c37;
6352	:douta	=	16'h	7d5b;
6353	:douta	=	16'h	7d3b;
6354	:douta	=	16'h	7d3b;
6355	:douta	=	16'h	7d5c;
6356	:douta	=	16'h	753b;
6357	:douta	=	16'h	74d9;
6358	:douta	=	16'h	6c37;
6359	:douta	=	16'h	4310;
6360	:douta	=	16'h	3a8e;
6361	:douta	=	16'h	31ca;
6362	:douta	=	16'h	10e4;
6363	:douta	=	16'h	0063;
6364	:douta	=	16'h	10e5;
6365	:douta	=	16'h	10e5;
6366	:douta	=	16'h	08c5;
6367	:douta	=	16'h	10c5;
6368	:douta	=	16'h	0884;
6369	:douta	=	16'h	29ca;
6370	:douta	=	16'h	42ef;
6371	:douta	=	16'h	7434;
6372	:douta	=	16'h	8473;
6373	:douta	=	16'h	7c33;
6374	:douta	=	16'h	9d35;
6375	:douta	=	16'h	ad77;
6376	:douta	=	16'h	7c53;
6377	:douta	=	16'h	5b50;
6378	:douta	=	16'h	7412;
6379	:douta	=	16'h	2a4e;
6380	:douta	=	16'h	2a4e;
6381	:douta	=	16'h	7433;
6382	:douta	=	16'h	4b11;
6383	:douta	=	16'h	8cb6;
6384	:douta	=	16'h	5bb4;
6385	:douta	=	16'h	4332;
6386	:douta	=	16'h	32b0;
6387	:douta	=	16'h	4332;
6388	:douta	=	16'h	2a6f;
6389	:douta	=	16'h	11cd;
6390	:douta	=	16'h	1a2f;
6391	:douta	=	16'h	851a;
6392	:douta	=	16'h	7497;
6393	:douta	=	16'h	9d7a;
6394	:douta	=	16'h	6c57;
6395	:douta	=	16'h	6436;
6396	:douta	=	16'h	7498;
6397	:douta	=	16'h	32d1;
6398	:douta	=	16'h	19cd;
6399	:douta	=	16'h	4b73;
6400	:douta	=	16'h	2ab1;
6401	:douta	=	16'h	224f;
6402	:douta	=	16'h	2a6f;
6403	:douta	=	16'h	6437;
6404	:douta	=	16'h	6416;
6405	:douta	=	16'h	5c37;
6406	:douta	=	16'h	7cb8;
6407	:douta	=	16'h	6415;
6408	:douta	=	16'h	5352;
6409	:douta	=	16'h	63d4;
6410	:douta	=	16'h	5bd5;
6411	:douta	=	16'h	7413;
6412	:douta	=	16'h	9d17;
6413	:douta	=	16'h	94b6;
6414	:douta	=	16'h	8cd6;
6415	:douta	=	16'h	8475;
6416	:douta	=	16'h	bdf9;
6417	:douta	=	16'h	7c96;
6418	:douta	=	16'h	6c35;
6419	:douta	=	16'h	8c74;
6420	:douta	=	16'h	9493;
6421	:douta	=	16'h	b5b7;
6422	:douta	=	16'h	bdf8;
6423	:douta	=	16'h	ad57;
6424	:douta	=	16'h	deb9;
6425	:douta	=	16'h	a598;
6426	:douta	=	16'h	9452;
6427	:douta	=	16'h	7c54;
6428	:douta	=	16'h	8c53;
6429	:douta	=	16'h	7c53;
6430	:douta	=	16'h	8c73;
6431	:douta	=	16'h	c638;
6432	:douta	=	16'h	c618;
6433	:douta	=	16'h	d678;
6434	:douta	=	16'h	8c73;
6435	:douta	=	16'h	94d4;
6436	:douta	=	16'h	4b0e;
6437	:douta	=	16'h	5b2f;
6438	:douta	=	16'h	c638;
6439	:douta	=	16'h	bdd6;
6440	:douta	=	16'h	ff9b;
6441	:douta	=	16'h	b5b6;
6442	:douta	=	16'h	b597;
6443	:douta	=	16'h	e698;
6444	:douta	=	16'h	de77;
6445	:douta	=	16'h	b5d7;
6446	:douta	=	16'h	a4b2;
6447	:douta	=	16'h	ce37;
6448	:douta	=	16'h	b573;
6449	:douta	=	16'h	b575;
6450	:douta	=	16'h	9c70;
6451	:douta	=	16'h	ef5a;
6452	:douta	=	16'h	8c50;
6453	:douta	=	16'h	bd74;
6454	:douta	=	16'h	3a2b;
6455	:douta	=	16'h	9430;
6456	:douta	=	16'h	ad32;
6457	:douta	=	16'h	c5f5;
6458	:douta	=	16'h	cdd4;
6459	:douta	=	16'h	d656;
6460	:douta	=	16'h	e6b8;
6461	:douta	=	16'h	9cd1;
6462	:douta	=	16'h	9c90;
6463	:douta	=	16'h	52cc;
6464	:douta	=	16'h	ce35;
6465	:douta	=	16'h	ad53;
6466	:douta	=	16'h	f719;
6467	:douta	=	16'h	ef59;
6468	:douta	=	16'h	bd33;
6469	:douta	=	16'h	6bce;
6470	:douta	=	16'h	4aac;
6471	:douta	=	16'h	c636;
6472	:douta	=	16'h	638e;
6473	:douta	=	16'h	bdf5;
6474	:douta	=	16'h	73d1;
6475	:douta	=	16'h	b534;
6476	:douta	=	16'h	7412;
6477	:douta	=	16'h	52f0;
6478	:douta	=	16'h	adb6;
6479	:douta	=	16'h	3a4c;
6480	:douta	=	16'h	a555;
6481	:douta	=	16'h	29eb;
6482	:douta	=	16'h	8451;
6483	:douta	=	16'h	9d76;
6484	:douta	=	16'h	adb6;
6485	:douta	=	16'h	8cd4;
6486	:douta	=	16'h	ef5c;
6487	:douta	=	16'h	9db8;
6488	:douta	=	16'h	8494;
6489	:douta	=	16'h	8495;
6490	:douta	=	16'h	5bb2;
6491	:douta	=	16'h	5b70;
6492	:douta	=	16'h	8c95;
6493	:douta	=	16'h	7c52;
6494	:douta	=	16'h	7497;
6495	:douta	=	16'h	4bb4;
6496	:douta	=	16'h	9ddb;
6497	:douta	=	16'h	3b34;
6498	:douta	=	16'h	5b91;
6499	:douta	=	16'h	42d0;
6500	:douta	=	16'h	5373;
6501	:douta	=	16'h	5373;
6502	:douta	=	16'h	5bf4;
6503	:douta	=	16'h	53b5;
6504	:douta	=	16'h	74d8;
6505	:douta	=	16'h	8518;
6506	:douta	=	16'h	857b;
6507	:douta	=	16'h	5416;
6508	:douta	=	16'h	9539;
6509	:douta	=	16'h	9db9;
6510	:douta	=	16'h	84d8;
6511	:douta	=	16'h	2a70;
6512	:douta	=	16'h	4b12;
6513	:douta	=	16'h	8d17;
6514	:douta	=	16'h	5bd4;
6515	:douta	=	16'h	7c95;
6516	:douta	=	16'h	6416;
6517	:douta	=	16'h	7c96;
6518	:douta	=	16'h	adda;
6519	:douta	=	16'h	8cf7;
6520	:douta	=	16'h	5352;
6521	:douta	=	16'h	426d;
6522	:douta	=	16'h	8412;
6523	:douta	=	16'h	3aaf;
6524	:douta	=	16'h	4ace;
6525	:douta	=	16'h	530f;
6526	:douta	=	16'h	7475;
6527	:douta	=	16'h	5b92;
6528	:douta	=	16'h	7453;
6529	:douta	=	16'h	add8;
6530	:douta	=	16'h	8497;
6531	:douta	=	16'h	ad34;
6532	:douta	=	16'h	c638;
6533	:douta	=	16'h	7bd0;
6534	:douta	=	16'h	8cf6;
6535	:douta	=	16'h	3a8d;
6536	:douta	=	16'h	324e;
6537	:douta	=	16'h	8453;
6538	:douta	=	16'h	7455;
6539	:douta	=	16'h	7c75;
6540	:douta	=	16'h	2126;
6541	:douta	=	16'h	2146;
6542	:douta	=	16'h	2126;
6543	:douta	=	16'h	2126;
6544	:douta	=	16'h	1926;
6545	:douta	=	16'h	1084;
6546	:douta	=	16'h	520a;
6547	:douta	=	16'h	62ab;
6548	:douta	=	16'h	634e;
6549	:douta	=	16'h	73d2;
6550	:douta	=	16'h	955a;
6551	:douta	=	16'h	8d5b;
6552	:douta	=	16'h	8d1a;
6553	:douta	=	16'h	7d19;
6554	:douta	=	16'h	7cd8;
6555	:douta	=	16'h	853a;
6556	:douta	=	16'h	851a;
6557	:douta	=	16'h	7cd9;
6558	:douta	=	16'h	8d7b;
6559	:douta	=	16'h	8d5b;
6560	:douta	=	16'h	8d5b;
6561	:douta	=	16'h	853a;
6562	:douta	=	16'h	853b;
6563	:douta	=	16'h	853a;
6564	:douta	=	16'h	855a;
6565	:douta	=	16'h	855a;
6566	:douta	=	16'h	7cf9;
6567	:douta	=	16'h	8d3a;
6568	:douta	=	16'h	853a;
6569	:douta	=	16'h	7d1a;
6570	:douta	=	16'h	7d3a;
6571	:douta	=	16'h	7d3a;
6572	:douta	=	16'h	7cfa;
6573	:douta	=	16'h	5bf6;
6574	:douta	=	16'h	6437;
6575	:douta	=	16'h	74b9;
6576	:douta	=	16'h	6c98;
6577	:douta	=	16'h	857b;
6578	:douta	=	16'h	5c37;
6579	:douta	=	16'h	6478;
6580	:douta	=	16'h	751a;
6581	:douta	=	16'h	7cfa;
6582	:douta	=	16'h	7498;
6583	:douta	=	16'h	74d9;
6584	:douta	=	16'h	7d1a;
6585	:douta	=	16'h	7d1b;
6586	:douta	=	16'h	7d3b;
6587	:douta	=	16'h	7d1a;
6588	:douta	=	16'h	6cba;
6589	:douta	=	16'h	855b;
6590	:douta	=	16'h	7d3a;
6591	:douta	=	16'h	7cfa;
6592	:douta	=	16'h	7d1a;
6593	:douta	=	16'h	7cf9;
6594	:douta	=	16'h	6c57;
6595	:douta	=	16'h	6c98;
6596	:douta	=	16'h	6cb9;
6597	:douta	=	16'h	6c99;
6598	:douta	=	16'h	7d3a;
6599	:douta	=	16'h	7d7b;
6600	:douta	=	16'h	6cb9;
6601	:douta	=	16'h	6cb8;
6602	:douta	=	16'h	857b;
6603	:douta	=	16'h	74d9;
6604	:douta	=	16'h	7d1a;
6605	:douta	=	16'h	7d3a;
6606	:douta	=	16'h	6478;
6607	:douta	=	16'h	7d3b;
6608	:douta	=	16'h	7d5b;
6609	:douta	=	16'h	751b;
6610	:douta	=	16'h	6478;
6611	:douta	=	16'h	6cfa;
6612	:douta	=	16'h	7d5b;
6613	:douta	=	16'h	7d3b;
6614	:douta	=	16'h	7d5c;
6615	:douta	=	16'h	6cb9;
6616	:douta	=	16'h	6cd9;
6617	:douta	=	16'h	6cb8;
6618	:douta	=	16'h	5372;
6619	:douta	=	16'h	42af;
6620	:douta	=	16'h	29ca;
6621	:douta	=	16'h	2147;
6622	:douta	=	16'h	08a4;
6623	:douta	=	16'h	10e6;
6624	:douta	=	16'h	10e5;
6625	:douta	=	16'h	1106;
6626	:douta	=	16'h	10e6;
6627	:douta	=	16'h	0085;
6628	:douta	=	16'h	9517;
6629	:douta	=	16'h	8cb6;
6630	:douta	=	16'h	6bf3;
6631	:douta	=	16'h	2a6f;
6632	:douta	=	16'h	326d;
6633	:douta	=	16'h	8452;
6634	:douta	=	16'h	94f5;
6635	:douta	=	16'h	73f3;
6636	:douta	=	16'h	326d;
6637	:douta	=	16'h	21ec;
6638	:douta	=	16'h	19ab;
6639	:douta	=	16'h	32b0;
6640	:douta	=	16'h	84d7;
6641	:douta	=	16'h	8d39;
6642	:douta	=	16'h	84b7;
6643	:douta	=	16'h	7cd8;
6644	:douta	=	16'h	9d9a;
6645	:douta	=	16'h	5416;
6646	:douta	=	16'h	4b74;
6647	:douta	=	16'h	32d2;
6648	:douta	=	16'h	3b13;
6649	:douta	=	16'h	32d2;
6650	:douta	=	16'h	3b32;
6651	:douta	=	16'h	7cb8;
6652	:douta	=	16'h	7497;
6653	:douta	=	16'h	8d7b;
6654	:douta	=	16'h	751a;
6655	:douta	=	16'h	7c97;
6656	:douta	=	16'h	3b34;
6657	:douta	=	16'h	5c57;
6658	:douta	=	16'h	3af1;
6659	:douta	=	16'h	6457;
6660	:douta	=	16'h	4b94;
6661	:douta	=	16'h	53b5;
6662	:douta	=	16'h	6c36;
6663	:douta	=	16'h	74b8;
6664	:douta	=	16'h	6c15;
6665	:douta	=	16'h	8d18;
6666	:douta	=	16'h	953a;
6667	:douta	=	16'h	6bd3;
6668	:douta	=	16'h	5330;
6669	:douta	=	16'h	6392;
6670	:douta	=	16'h	7c34;
6671	:douta	=	16'h	8475;
6672	:douta	=	16'h	ce39;
6673	:douta	=	16'h	c63a;
6674	:douta	=	16'h	add9;
6675	:douta	=	16'h	7433;
6676	:douta	=	16'h	73d1;
6677	:douta	=	16'h	63b1;
6678	:douta	=	16'h	73f2;
6679	:douta	=	16'h	9cf5;
6680	:douta	=	16'h	eefa;
6681	:douta	=	16'h	c639;
6682	:douta	=	16'h	bd76;
6683	:douta	=	16'h	d69a;
6684	:douta	=	16'h	9cd5;
6685	:douta	=	16'h	b5d8;
6686	:douta	=	16'h	6bf3;
6687	:douta	=	16'h	8cb4;
6688	:douta	=	16'h	94d5;
6689	:douta	=	16'h	de99;
6690	:douta	=	16'h	d679;
6691	:douta	=	16'h	deb8;
6692	:douta	=	16'h	4aae;
6693	:douta	=	16'h	73f1;
6694	:douta	=	16'h	9d15;
6695	:douta	=	16'h	8c52;
6696	:douta	=	16'h	94d4;
6697	:douta	=	16'h	b5b5;
6698	:douta	=	16'h	b554;
6699	:douta	=	16'h	ce36;
6700	:douta	=	16'h	fffc;
6701	:douta	=	16'h	de98;
6702	:douta	=	16'h	bdb5;
6703	:douta	=	16'h	de78;
6704	:douta	=	16'h	a514;
6705	:douta	=	16'h	636f;
6706	:douta	=	16'h	9450;
6707	:douta	=	16'h	de97;
6708	:douta	=	16'h	b552;
6709	:douta	=	16'h	f77a;
6710	:douta	=	16'h	9410;
6711	:douta	=	16'h	cdf5;
6712	:douta	=	16'h	5b6f;
6713	:douta	=	16'h	31a8;
6714	:douta	=	16'h	63af;
6715	:douta	=	16'h	ef18;
6716	:douta	=	16'h	e6d8;
6717	:douta	=	16'h	d655;
6718	:douta	=	16'h	c5d4;
6719	:douta	=	16'h	8c0e;
6720	:douta	=	16'h	bdd4;
6721	:douta	=	16'h	8c4f;
6722	:douta	=	16'h	ad31;
6723	:douta	=	16'h	be15;
6724	:douta	=	16'h	bd93;
6725	:douta	=	16'h	bd93;
6726	:douta	=	16'h	634d;
6727	:douta	=	16'h	c615;
6728	:douta	=	16'h	328c;
6729	:douta	=	16'h	c616;
6730	:douta	=	16'h	4a8d;
6731	:douta	=	16'h	acd3;
6732	:douta	=	16'h	94b4;
6733	:douta	=	16'h	94b4;
6734	:douta	=	16'h	be59;
6735	:douta	=	16'h	52ef;
6736	:douta	=	16'h	7c11;
6737	:douta	=	16'h	29ca;
6738	:douta	=	16'h	6b90;
6739	:douta	=	16'h	5b4e;
6740	:douta	=	16'h	4a8c;
6741	:douta	=	16'h	7410;
6742	:douta	=	16'h	9d14;
6743	:douta	=	16'h	9515;
6744	:douta	=	16'h	4b2f;
6745	:douta	=	16'h	7474;
6746	:douta	=	16'h	7496;
6747	:douta	=	16'h	63b1;
6748	:douta	=	16'h	8cb5;
6749	:douta	=	16'h	5371;
6750	:douta	=	16'h	328e;
6751	:douta	=	16'h	4b73;
6752	:douta	=	16'h	74d8;
6753	:douta	=	16'h	4b94;
6754	:douta	=	16'h	84f7;
6755	:douta	=	16'h	53d4;
6756	:douta	=	16'h	6c15;
6757	:douta	=	16'h	7435;
6758	:douta	=	16'h	6c56;
6759	:douta	=	16'h	3b11;
6760	:douta	=	16'h	4b52;
6761	:douta	=	16'h	5c15;
6762	:douta	=	16'h	5c16;
6763	:douta	=	16'h	3af1;
6764	:douta	=	16'h	8d39;
6765	:douta	=	16'h	a63d;
6766	:douta	=	16'h	8d38;
6767	:douta	=	16'h	32b1;
6768	:douta	=	16'h	326f;
6769	:douta	=	16'h	5c14;
6770	:douta	=	16'h	52f0;
6771	:douta	=	16'h	4b52;
6772	:douta	=	16'h	7497;
6773	:douta	=	16'h	84d7;
6774	:douta	=	16'h	84d6;
6775	:douta	=	16'h	7496;
6776	:douta	=	16'h	7476;
6777	:douta	=	16'h	6c14;
6778	:douta	=	16'h	ad96;
6779	:douta	=	16'h	7c96;
6780	:douta	=	16'h	8495;
6781	:douta	=	16'h	322c;
6782	:douta	=	16'h	52ef;
6783	:douta	=	16'h	73d1;
6784	:douta	=	16'h	63b2;
6785	:douta	=	16'h	3aaf;
6786	:douta	=	16'h	94f5;
6787	:douta	=	16'h	9d36;
6788	:douta	=	16'h	8cf5;
6789	:douta	=	16'h	be19;
6790	:douta	=	16'h	7c96;
6791	:douta	=	16'h	8cb7;
6792	:douta	=	16'h	5b93;
6793	:douta	=	16'h	8cf7;
6794	:douta	=	16'h	31ea;
6795	:douta	=	16'h	1926;
6796	:douta	=	16'h	2146;
6797	:douta	=	16'h	2126;
6798	:douta	=	16'h	2146;
6799	:douta	=	16'h	10c4;
6800	:douta	=	16'h	1063;
6801	:douta	=	16'h	524a;
6802	:douta	=	16'h	7b8f;
6803	:douta	=	16'h	6b70;
6804	:douta	=	16'h	84b7;
6805	:douta	=	16'h	7c98;
6806	:douta	=	16'h	853a;
6807	:douta	=	16'h	74b9;
6808	:douta	=	16'h	8d1a;
6809	:douta	=	16'h	8d5b;
6810	:douta	=	16'h	853a;
6811	:douta	=	16'h	8519;
6812	:douta	=	16'h	8d3a;
6813	:douta	=	16'h	7cf9;
6814	:douta	=	16'h	8519;
6815	:douta	=	16'h	8519;
6816	:douta	=	16'h	853b;
6817	:douta	=	16'h	8d7b;
6818	:douta	=	16'h	8d5b;
6819	:douta	=	16'h	851a;
6820	:douta	=	16'h	851a;
6821	:douta	=	16'h	853a;
6822	:douta	=	16'h	7c77;
6823	:douta	=	16'h	7c97;
6824	:douta	=	16'h	851a;
6825	:douta	=	16'h	7cf9;
6826	:douta	=	16'h	74b9;
6827	:douta	=	16'h	7d1a;
6828	:douta	=	16'h	8d7b;
6829	:douta	=	16'h	74fa;
6830	:douta	=	16'h	74ba;
6831	:douta	=	16'h	74fa;
6832	:douta	=	16'h	6cb9;
6833	:douta	=	16'h	7d1b;
6834	:douta	=	16'h	7d3a;
6835	:douta	=	16'h	6478;
6836	:douta	=	16'h	751a;
6837	:douta	=	16'h	857b;
6838	:douta	=	16'h	74da;
6839	:douta	=	16'h	74fa;
6840	:douta	=	16'h	7d1b;
6841	:douta	=	16'h	74d9;
6842	:douta	=	16'h	7d3a;
6843	:douta	=	16'h	7d3a;
6844	:douta	=	16'h	7d3a;
6845	:douta	=	16'h	74ba;
6846	:douta	=	16'h	751a;
6847	:douta	=	16'h	8d9c;
6848	:douta	=	16'h	7d1a;
6849	:douta	=	16'h	74b8;
6850	:douta	=	16'h	74b9;
6851	:douta	=	16'h	7d1a;
6852	:douta	=	16'h	74b9;
6853	:douta	=	16'h	6c99;
6854	:douta	=	16'h	6cb8;
6855	:douta	=	16'h	6478;
6856	:douta	=	16'h	7d1b;
6857	:douta	=	16'h	7d1a;
6858	:douta	=	16'h	85bc;
6859	:douta	=	16'h	7d1a;
6860	:douta	=	16'h	6cb9;
6861	:douta	=	16'h	95dc;
6862	:douta	=	16'h	8dbc;
6863	:douta	=	16'h	6cd9;
6864	:douta	=	16'h	6cd9;
6865	:douta	=	16'h	859c;
6866	:douta	=	16'h	6cd9;
6867	:douta	=	16'h	6cda;
6868	:douta	=	16'h	753b;
6869	:douta	=	16'h	6cda;
6870	:douta	=	16'h	6cba;
6871	:douta	=	16'h	7d7c;
6872	:douta	=	16'h	74fa;
6873	:douta	=	16'h	6cba;
6874	:douta	=	16'h	74d9;
6875	:douta	=	16'h	6c16;
6876	:douta	=	16'h	42cf;
6877	:douta	=	16'h	320b;
6878	:douta	=	16'h	2168;
6879	:douta	=	16'h	0884;
6880	:douta	=	16'h	10c5;
6881	:douta	=	16'h	10e5;
6882	:douta	=	16'h	10e6;
6883	:douta	=	16'h	10c4;
6884	:douta	=	16'h	1169;
6885	:douta	=	16'h	4b50;
6886	:douta	=	16'h	a557;
6887	:douta	=	16'h	6bd3;
6888	:douta	=	16'h	6bb1;
6889	:douta	=	16'h	322c;
6890	:douta	=	16'h	4b0f;
6891	:douta	=	16'h	b5d8;
6892	:douta	=	16'h	63b2;
6893	:douta	=	16'h	73f2;
6894	:douta	=	16'h	222f;
6895	:douta	=	16'h	3af1;
6896	:douta	=	16'h	2a6e;
6897	:douta	=	16'h	4b31;
6898	:douta	=	16'h	5392;
6899	:douta	=	16'h	7498;
6900	:douta	=	16'h	7cd9;
6901	:douta	=	16'h	74b8;
6902	:douta	=	16'h	9559;
6903	:douta	=	16'h	8cf8;
6904	:douta	=	16'h	6478;
6905	:douta	=	16'h	3ad1;
6906	:douta	=	16'h	4332;
6907	:douta	=	16'h	4b95;
6908	:douta	=	16'h	32b0;
6909	:douta	=	16'h	5c17;
6910	:douta	=	16'h	6478;
6911	:douta	=	16'h	a5bc;
6912	:douta	=	16'h	224f;
6913	:douta	=	16'h	116c;
6914	:douta	=	16'h	32b0;
6915	:douta	=	16'h	6415;
6916	:douta	=	16'h	6415;
6917	:douta	=	16'h	53b5;
6918	:douta	=	16'h	5bf5;
6919	:douta	=	16'h	6c57;
6920	:douta	=	16'h	4b11;
6921	:douta	=	16'h	4311;
6922	:douta	=	16'h	4b73;
6923	:douta	=	16'h	6bd4;
6924	:douta	=	16'h	9cb6;
6925	:douta	=	16'h	9517;
6926	:douta	=	16'h	8cb5;
6927	:douta	=	16'h	6bf4;
6928	:douta	=	16'h	ce39;
6929	:douta	=	16'h	add9;
6930	:douta	=	16'h	8474;
6931	:douta	=	16'h	5b92;
6932	:douta	=	16'h	a536;
6933	:douta	=	16'h	9cf5;
6934	:douta	=	16'h	d659;
6935	:douta	=	16'h	ad97;
6936	:douta	=	16'h	bd97;
6937	:douta	=	16'h	94f5;
6938	:douta	=	16'h	ad76;
6939	:douta	=	16'h	b5b7;
6940	:douta	=	16'h	8cb5;
6941	:douta	=	16'h	d678;
6942	:douta	=	16'h	94d5;
6943	:douta	=	16'h	ffdb;
6944	:douta	=	16'h	b5b7;
6945	:douta	=	16'h	e6d9;
6946	:douta	=	16'h	8473;
6947	:douta	=	16'h	a534;
6948	:douta	=	16'h	8c73;
6949	:douta	=	16'h	ce16;
6950	:douta	=	16'h	b5d6;
6951	:douta	=	16'h	ff7b;
6952	:douta	=	16'h	ffbc;
6953	:douta	=	16'h	634f;
6954	:douta	=	16'h	c5b4;
6955	:douta	=	16'h	4acd;
6956	:douta	=	16'h	83ef;
6957	:douta	=	16'h	8471;
6958	:douta	=	16'h	9c92;
6959	:douta	=	16'h	de98;
6960	:douta	=	16'h	ce16;
6961	:douta	=	16'h	94b2;
6962	:douta	=	16'h	8bce;
6963	:douta	=	16'h	ce57;
6964	:douta	=	16'h	634e;
6965	:douta	=	16'h	94b0;
6966	:douta	=	16'h	428a;
6967	:douta	=	16'h	bd74;
6968	:douta	=	16'h	946f;
6969	:douta	=	16'h	f71a;
6970	:douta	=	16'h	a4b1;
6971	:douta	=	16'h	a4d0;
6972	:douta	=	16'h	bd72;
6973	:douta	=	16'h	4a28;
6974	:douta	=	16'h	6b8c;
6975	:douta	=	16'h	5b0c;
6976	:douta	=	16'h	b593;
6977	:douta	=	16'h	9470;
6978	:douta	=	16'h	fffb;
6979	:douta	=	16'h	840f;
6980	:douta	=	16'h	d615;
6981	:douta	=	16'h	7c10;
6982	:douta	=	16'h	630c;
6983	:douta	=	16'h	94b2;
6984	:douta	=	16'h	634d;
6985	:douta	=	16'h	c636;
6986	:douta	=	16'h	5b0e;
6987	:douta	=	16'h	de77;
6988	:douta	=	16'h	5b50;
6989	:douta	=	16'h	7bf1;
6990	:douta	=	16'h	5b90;
6991	:douta	=	16'h	5aaa;
6992	:douta	=	16'h	a4f3;
6993	:douta	=	16'h	6b2d;
6994	:douta	=	16'h	bd94;
6995	:douta	=	16'h	3a2a;
6996	:douta	=	16'h	7c11;
6997	:douta	=	16'h	a512;
6998	:douta	=	16'h	63b0;
6999	:douta	=	16'h	324d;
7000	:douta	=	16'h	4b71;
7001	:douta	=	16'h	32b0;
7002	:douta	=	16'h	0044;
7003	:douta	=	16'h	5bb3;
7004	:douta	=	16'h	3b11;
7005	:douta	=	16'h	7496;
7006	:douta	=	16'h	5393;
7007	:douta	=	16'h	5372;
7008	:douta	=	16'h	6414;
7009	:douta	=	16'h	3ad0;
7010	:douta	=	16'h	42f0;
7011	:douta	=	16'h	4311;
7012	:douta	=	16'h	5351;
7013	:douta	=	16'h	74b7;
7014	:douta	=	16'h	7519;
7015	:douta	=	16'h	4bd6;
7016	:douta	=	16'h	957a;
7017	:douta	=	16'h	5c37;
7018	:douta	=	16'h	859d;
7019	:douta	=	16'h	5395;
7020	:douta	=	16'h	4aaf;
7021	:douta	=	16'h	1949;
7022	:douta	=	16'h	3ad1;
7023	:douta	=	16'h	53d5;
7024	:douta	=	16'h	53b4;
7025	:douta	=	16'h	7cb6;
7026	:douta	=	16'h	7cb6;
7027	:douta	=	16'h	53f5;
7028	:douta	=	16'h	5b73;
7029	:douta	=	16'h	7433;
7030	:douta	=	16'h	6456;
7031	:douta	=	16'h	42b0;
7032	:douta	=	16'h	2a4e;
7033	:douta	=	16'h	2a0c;
7034	:douta	=	16'h	5b91;
7035	:douta	=	16'h	4b11;
7036	:douta	=	16'h	6bf2;
7037	:douta	=	16'h	5b91;
7038	:douta	=	16'h	a598;
7039	:douta	=	16'h	a578;
7040	:douta	=	16'h	9d77;
7041	:douta	=	16'h	a5d9;
7042	:douta	=	16'h	6392;
7043	:douta	=	16'h	324e;
7044	:douta	=	16'h	5b50;
7045	:douta	=	16'h	42ae;
7046	:douta	=	16'h	5b71;
7047	:douta	=	16'h	5b71;
7048	:douta	=	16'h	3a4b;
7049	:douta	=	16'h	2146;
7050	:douta	=	16'h	2966;
7051	:douta	=	16'h	2966;
7052	:douta	=	16'h	2146;
7053	:douta	=	16'h	18a4;
7054	:douta	=	16'h	49e8;
7055	:douta	=	16'h	7b6e;
7056	:douta	=	16'h	8cb5;
7057	:douta	=	16'h	8cf8;
7058	:douta	=	16'h	7498;
7059	:douta	=	16'h	8519;
7060	:douta	=	16'h	953a;
7061	:douta	=	16'h	8d19;
7062	:douta	=	16'h	7d19;
7063	:douta	=	16'h	851a;
7064	:douta	=	16'h	8d5b;
7065	:douta	=	16'h	8d3a;
7066	:douta	=	16'h	851a;
7067	:douta	=	16'h	851a;
7068	:douta	=	16'h	8d7b;
7069	:douta	=	16'h	8d3a;
7070	:douta	=	16'h	8d5b;
7071	:douta	=	16'h	851a;
7072	:douta	=	16'h	853a;
7073	:douta	=	16'h	7cd9;
7074	:douta	=	16'h	8519;
7075	:douta	=	16'h	8d5b;
7076	:douta	=	16'h	853a;
7077	:douta	=	16'h	7cd8;
7078	:douta	=	16'h	855a;
7079	:douta	=	16'h	8d7b;
7080	:douta	=	16'h	8519;
7081	:douta	=	16'h	851a;
7082	:douta	=	16'h	959b;
7083	:douta	=	16'h	8d7b;
7084	:douta	=	16'h	853a;
7085	:douta	=	16'h	7cf9;
7086	:douta	=	16'h	853a;
7087	:douta	=	16'h	6cb9;
7088	:douta	=	16'h	6458;
7089	:douta	=	16'h	5c17;
7090	:douta	=	16'h	6438;
7091	:douta	=	16'h	6c99;
7092	:douta	=	16'h	6478;
7093	:douta	=	16'h	6478;
7094	:douta	=	16'h	6c99;
7095	:douta	=	16'h	7d3b;
7096	:douta	=	16'h	6478;
7097	:douta	=	16'h	6478;
7098	:douta	=	16'h	7d1b;
7099	:douta	=	16'h	7d3a;
7100	:douta	=	16'h	8dbc;
7101	:douta	=	16'h	859d;
7102	:douta	=	16'h	95dd;
7103	:douta	=	16'h	7d3a;
7104	:douta	=	16'h	7d1a;
7105	:douta	=	16'h	8dbc;
7106	:douta	=	16'h	855b;
7107	:douta	=	16'h	855a;
7108	:douta	=	16'h	7d1a;
7109	:douta	=	16'h	855b;
7110	:douta	=	16'h	6cd9;
7111	:douta	=	16'h	6c99;
7112	:douta	=	16'h	8d9b;
7113	:douta	=	16'h	855a;
7114	:douta	=	16'h	6478;
7115	:douta	=	16'h	7d1a;
7116	:douta	=	16'h	74da;
7117	:douta	=	16'h	751a;
7118	:douta	=	16'h	7d3a;
7119	:douta	=	16'h	7d1a;
7120	:douta	=	16'h	7d1a;
7121	:douta	=	16'h	6457;
7122	:douta	=	16'h	6478;
7123	:douta	=	16'h	751a;
7124	:douta	=	16'h	753b;
7125	:douta	=	16'h	74d9;
7126	:douta	=	16'h	6478;
7127	:douta	=	16'h	74d9;
7128	:douta	=	16'h	74f9;
7129	:douta	=	16'h	755c;
7130	:douta	=	16'h	74fb;
7131	:douta	=	16'h	751a;
7132	:douta	=	16'h	6cda;
7133	:douta	=	16'h	74da;
7134	:douta	=	16'h	5353;
7135	:douta	=	16'h	29aa;
7136	:douta	=	16'h	2168;
7137	:douta	=	16'h	10e5;
7138	:douta	=	16'h	08c5;
7139	:douta	=	16'h	1107;
7140	:douta	=	16'h	1127;
7141	:douta	=	16'h	1106;
7142	:douta	=	16'h	00c6;
7143	:douta	=	16'h	42ee;
7144	:douta	=	16'h	a516;
7145	:douta	=	16'h	73f2;
7146	:douta	=	16'h	73f4;
7147	:douta	=	16'h	19ab;
7148	:douta	=	16'h	42d0;
7149	:douta	=	16'h	326e;
7150	:douta	=	16'h	b63b;
7151	:douta	=	16'h	9d79;
7152	:douta	=	16'h	73f4;
7153	:douta	=	16'h	9d37;
7154	:douta	=	16'h	6416;
7155	:douta	=	16'h	5c38;
7156	:douta	=	16'h	4374;
7157	:douta	=	16'h	3b54;
7158	:douta	=	16'h	2ad2;
7159	:douta	=	16'h	6c97;
7160	:douta	=	16'h	7c76;
7161	:douta	=	16'h	adba;
7162	:douta	=	16'h	6cb9;
7163	:douta	=	16'h	6c57;
7164	:douta	=	16'h	32f2;
7165	:douta	=	16'h	2a4f;
7166	:douta	=	16'h	2a8f;
7167	:douta	=	16'h	3b12;
7168	:douta	=	16'h	3b33;
7169	:douta	=	16'h	4b94;
7170	:douta	=	16'h	2a90;
7171	:douta	=	16'h	6436;
7172	:douta	=	16'h	5bd4;
7173	:douta	=	16'h	5bd5;
7174	:douta	=	16'h	5b94;
7175	:douta	=	16'h	7d19;
7176	:douta	=	16'h	5b92;
7177	:douta	=	16'h	7c76;
7178	:douta	=	16'h	8d19;
7179	:douta	=	16'h	5b93;
7180	:douta	=	16'h	5330;
7181	:douta	=	16'h	5b71;
7182	:douta	=	16'h	6c14;
7183	:douta	=	16'h	6bd3;
7184	:douta	=	16'h	bdd7;
7185	:douta	=	16'h	ef1c;
7186	:douta	=	16'h	a577;
7187	:douta	=	16'h	84b6;
7188	:douta	=	16'h	6bb1;
7189	:douta	=	16'h	73f3;
7190	:douta	=	16'h	7c32;
7191	:douta	=	16'h	7412;
7192	:douta	=	16'h	e6b9;
7193	:douta	=	16'h	c639;
7194	:douta	=	16'h	b596;
7195	:douta	=	16'h	ce59;
7196	:douta	=	16'h	6bd2;
7197	:douta	=	16'h	7c53;
7198	:douta	=	16'h	6bf3;
7199	:douta	=	16'h	b596;
7200	:douta	=	16'h	b556;
7201	:douta	=	16'h	e6f9;
7202	:douta	=	16'h	b576;
7203	:douta	=	16'h	b5b6;
7204	:douta	=	16'h	52ef;
7205	:douta	=	16'h	530e;
7206	:douta	=	16'h	b5f8;
7207	:douta	=	16'h	c5d6;
7208	:douta	=	16'h	ffbb;
7209	:douta	=	16'h	bd73;
7210	:douta	=	16'h	ef19;
7211	:douta	=	16'h	b575;
7212	:douta	=	16'h	a4b3;
7213	:douta	=	16'h	bdd6;
7214	:douta	=	16'h	62ee;
7215	:douta	=	16'h	cdd6;
7216	:douta	=	16'h	a4f3;
7217	:douta	=	16'h	a491;
7218	:douta	=	16'h	e696;
7219	:douta	=	16'h	d676;
7220	:douta	=	16'h	7bed;
7221	:douta	=	16'h	ef18;
7222	:douta	=	16'h	528b;
7223	:douta	=	16'h	8c0f;
7224	:douta	=	16'h	840f;
7225	:douta	=	16'h	9cb1;
7226	:douta	=	16'h	ad31;
7227	:douta	=	16'h	eef8;
7228	:douta	=	16'h	e6f8;
7229	:douta	=	16'h	e676;
7230	:douta	=	16'h	c615;
7231	:douta	=	16'h	41c8;
7232	:douta	=	16'h	b593;
7233	:douta	=	16'h	52eb;
7234	:douta	=	16'h	e6d7;
7235	:douta	=	16'h	ad10;
7236	:douta	=	16'h	ef18;
7237	:douta	=	16'h	94b0;
7238	:douta	=	16'h	734c;
7239	:douta	=	16'h	8cd3;
7240	:douta	=	16'h	2a0a;
7241	:douta	=	16'h	b594;
7242	:douta	=	16'h	4aad;
7243	:douta	=	16'h	bd95;
7244	:douta	=	16'h	73d1;
7245	:douta	=	16'h	b554;
7246	:douta	=	16'h	6bf1;
7247	:douta	=	16'h	7bcf;
7248	:douta	=	16'h	8410;
7249	:douta	=	16'h	31c9;
7250	:douta	=	16'h	7bcf;
7251	:douta	=	16'h	4a8b;
7252	:douta	=	16'h	29a7;
7253	:douta	=	16'h	52aa;
7254	:douta	=	16'h	3a8d;
7255	:douta	=	16'h	31ea;
7256	:douta	=	16'h	3acf;
7257	:douta	=	16'h	42f0;
7258	:douta	=	16'h	29aa;
7259	:douta	=	16'h	00c6;
7260	:douta	=	16'h	1968;
7261	:douta	=	16'h	4b31;
7262	:douta	=	16'h	2a2d;
7263	:douta	=	16'h	5373;
7264	:douta	=	16'h	6415;
7265	:douta	=	16'h	5394;
7266	:douta	=	16'h	5352;
7267	:douta	=	16'h	222d;
7268	:douta	=	16'h	5b71;
7269	:douta	=	16'h	6bd3;
7270	:douta	=	16'h	5c15;
7271	:douta	=	16'h	4b73;
7272	:douta	=	16'h	63f4;
7273	:douta	=	16'h	53d5;
7274	:douta	=	16'h	4bf6;
7275	:douta	=	16'h	3b13;
7276	:douta	=	16'h	8d59;
7277	:douta	=	16'h	5bd3;
7278	:douta	=	16'h	4b74;
7279	:douta	=	16'h	3af2;
7280	:douta	=	16'h	32d1;
7281	:douta	=	16'h	6c14;
7282	:douta	=	16'h	5bb4;
7283	:douta	=	16'h	2a4e;
7284	:douta	=	16'h	8d7a;
7285	:douta	=	16'h	9517;
7286	:douta	=	16'h	7cd8;
7287	:douta	=	16'h	63d3;
7288	:douta	=	16'h	5372;
7289	:douta	=	16'h	6330;
7290	:douta	=	16'h	7c55;
7291	:douta	=	16'h	7413;
7292	:douta	=	16'h	6b91;
7293	:douta	=	16'h	5b92;
7294	:douta	=	16'h	7453;
7295	:douta	=	16'h	5b91;
7296	:douta	=	16'h	9d77;
7297	:douta	=	16'h	9579;
7298	:douta	=	16'h	8cf5;
7299	:douta	=	16'h	4312;
7300	:douta	=	16'h	4310;
7301	:douta	=	16'h	7454;
7302	:douta	=	16'h	4b10;
7303	:douta	=	16'h	5350;
7304	:douta	=	16'h	2105;
7305	:douta	=	16'h	2966;
7306	:douta	=	16'h	2967;
7307	:douta	=	16'h	2145;
7308	:douta	=	16'h	10a4;
7309	:douta	=	16'h	6aab;
7310	:douta	=	16'h	83af;
7311	:douta	=	16'h	73d1;
7312	:douta	=	16'h	7c96;
7313	:douta	=	16'h	7cd8;
7314	:douta	=	16'h	7498;
7315	:douta	=	16'h	7457;
7316	:douta	=	16'h	8d3a;
7317	:douta	=	16'h	9d9b;
7318	:douta	=	16'h	851a;
7319	:douta	=	16'h	8519;
7320	:douta	=	16'h	7cf9;
7321	:douta	=	16'h	9d9b;
7322	:douta	=	16'h	959c;
7323	:douta	=	16'h	7cf9;
7324	:douta	=	16'h	853a;
7325	:douta	=	16'h	855a;
7326	:douta	=	16'h	8d7b;
7327	:douta	=	16'h	959b;
7328	:douta	=	16'h	8d5b;
7329	:douta	=	16'h	8d3a;
7330	:douta	=	16'h	7cf9;
7331	:douta	=	16'h	8d5a;
7332	:douta	=	16'h	851a;
7333	:douta	=	16'h	7c98;
7334	:douta	=	16'h	95bc;
7335	:douta	=	16'h	8d7b;
7336	:douta	=	16'h	851a;
7337	:douta	=	16'h	8d5b;
7338	:douta	=	16'h	8d7b;
7339	:douta	=	16'h	8d5a;
7340	:douta	=	16'h	95bc;
7341	:douta	=	16'h	853a;
7342	:douta	=	16'h	7cf9;
7343	:douta	=	16'h	7d3b;
7344	:douta	=	16'h	7cd9;
7345	:douta	=	16'h	6c79;
7346	:douta	=	16'h	6498;
7347	:douta	=	16'h	859c;
7348	:douta	=	16'h	6cba;
7349	:douta	=	16'h	5c38;
7350	:douta	=	16'h	4b75;
7351	:douta	=	16'h	7d7c;
7352	:douta	=	16'h	9e5f;
7353	:douta	=	16'h	5c58;
7354	:douta	=	16'h	6499;
7355	:douta	=	16'h	74d9;
7356	:douta	=	16'h	74fa;
7357	:douta	=	16'h	855b;
7358	:douta	=	16'h	95bc;
7359	:douta	=	16'h	961d;
7360	:douta	=	16'h	7d3b;
7361	:douta	=	16'h	7d5b;
7362	:douta	=	16'h	857b;
7363	:douta	=	16'h	857b;
7364	:douta	=	16'h	8d9b;
7365	:douta	=	16'h	7d1a;
7366	:douta	=	16'h	8d9b;
7367	:douta	=	16'h	855b;
7368	:douta	=	16'h	74f9;
7369	:douta	=	16'h	85bc;
7370	:douta	=	16'h	74d9;
7371	:douta	=	16'h	7cfa;
7372	:douta	=	16'h	7d1a;
7373	:douta	=	16'h	6c98;
7374	:douta	=	16'h	6c98;
7375	:douta	=	16'h	6498;
7376	:douta	=	16'h	7d1a;
7377	:douta	=	16'h	7d3a;
7378	:douta	=	16'h	74d9;
7379	:douta	=	16'h	74d9;
7380	:douta	=	16'h	6498;
7381	:douta	=	16'h	857b;
7382	:douta	=	16'h	6c98;
7383	:douta	=	16'h	6c98;
7384	:douta	=	16'h	6cb9;
7385	:douta	=	16'h	74da;
7386	:douta	=	16'h	753b;
7387	:douta	=	16'h	751a;
7388	:douta	=	16'h	6cfa;
7389	:douta	=	16'h	6cda;
7390	:douta	=	16'h	74fa;
7391	:douta	=	16'h	5332;
7392	:douta	=	16'h	324d;
7393	:douta	=	16'h	2168;
7394	:douta	=	16'h	2168;
7395	:douta	=	16'h	08c5;
7396	:douta	=	16'h	1106;
7397	:douta	=	16'h	1126;
7398	:douta	=	16'h	10e7;
7399	:douta	=	16'h	08e6;
7400	:douta	=	16'h	4310;
7401	:douta	=	16'h	be19;
7402	:douta	=	16'h	94b6;
7403	:douta	=	16'h	5351;
7404	:douta	=	16'h	5372;
7405	:douta	=	16'h	4b10;
7406	:douta	=	16'h	42f1;
7407	:douta	=	16'h	4b11;
7408	:douta	=	16'h	9d16;
7409	:douta	=	16'h	9d38;
7410	:douta	=	16'h	955a;
7411	:douta	=	16'h	6c98;
7412	:douta	=	16'h	74b8;
7413	:douta	=	16'h	4b75;
7414	:douta	=	16'h	53d5;
7415	:douta	=	16'h	2291;
7416	:douta	=	16'h	7cb7;
7417	:douta	=	16'h	8cd7;
7418	:douta	=	16'h	84d8;
7419	:douta	=	16'h	a59a;
7420	:douta	=	16'h	5c16;
7421	:douta	=	16'h	8d5a;
7422	:douta	=	16'h	6477;
7423	:douta	=	16'h	53d4;
7424	:douta	=	16'h	222e;
7425	:douta	=	16'h	32d2;
7426	:douta	=	16'h	2ab1;
7427	:douta	=	16'h	6c37;
7428	:douta	=	16'h	74b8;
7429	:douta	=	16'h	6c36;
7430	:douta	=	16'h	74b8;
7431	:douta	=	16'h	5bb4;
7432	:douta	=	16'h	42f0;
7433	:douta	=	16'h	5b73;
7434	:douta	=	16'h	6415;
7435	:douta	=	16'h	7435;
7436	:douta	=	16'h	94d6;
7437	:douta	=	16'h	9517;
7438	:douta	=	16'h	9d37;
7439	:douta	=	16'h	7434;
7440	:douta	=	16'h	9cf5;
7441	:douta	=	16'h	7413;
7442	:douta	=	16'h	7c75;
7443	:douta	=	16'h	5b92;
7444	:douta	=	16'h	ad56;
7445	:douta	=	16'h	d679;
7446	:douta	=	16'h	bdd7;
7447	:douta	=	16'h	bdf8;
7448	:douta	=	16'h	9cd5;
7449	:douta	=	16'h	c5f7;
7450	:douta	=	16'h	a556;
7451	:douta	=	16'h	a515;
7452	:douta	=	16'h	9d15;
7453	:douta	=	16'h	e6f9;
7454	:douta	=	16'h	ce58;
7455	:douta	=	16'h	c658;
7456	:douta	=	16'h	5350;
7457	:douta	=	16'h	c5f7;
7458	:douta	=	16'h	8473;
7459	:douta	=	16'h	8c51;
7460	:douta	=	16'h	c5f7;
7461	:douta	=	16'h	de98;
7462	:douta	=	16'h	ad96;
7463	:douta	=	16'h	f71a;
7464	:douta	=	16'h	c638;
7465	:douta	=	16'h	8452;
7466	:douta	=	16'h	73d0;
7467	:douta	=	16'h	8430;
7468	:douta	=	16'h	deb8;
7469	:douta	=	16'h	d6b8;
7470	:douta	=	16'h	d636;
7471	:douta	=	16'h	f73a;
7472	:douta	=	16'h	ce16;
7473	:douta	=	16'h	638f;
7474	:douta	=	16'h	2969;
7475	:douta	=	16'h	9512;
7476	:douta	=	16'h	424c;
7477	:douta	=	16'h	ad73;
7478	:douta	=	16'h	acd0;
7479	:douta	=	16'h	eeb7;
7480	:douta	=	16'h	840d;
7481	:douta	=	16'h	b4b0;
7482	:douta	=	16'h	94b0;
7483	:douta	=	16'h	bd72;
7484	:douta	=	16'h	8cb0;
7485	:douta	=	16'h	a46e;
7486	:douta	=	16'h	94b1;
7487	:douta	=	16'h	6b8d;
7488	:douta	=	16'h	bdf5;
7489	:douta	=	16'h	ad11;
7490	:douta	=	16'h	d695;
7491	:douta	=	16'h	634d;
7492	:douta	=	16'h	d655;
7493	:douta	=	16'h	52aa;
7494	:douta	=	16'h	62cb;
7495	:douta	=	16'h	94b2;
7496	:douta	=	16'h	736e;
7497	:douta	=	16'h	b5b4;
7498	:douta	=	16'h	a4b1;
7499	:douta	=	16'h	e6d7;
7500	:douta	=	16'h	4a8b;
7501	:douta	=	16'h	738f;
7502	:douta	=	16'h	426b;
7503	:douta	=	16'h	9c91;
7504	:douta	=	16'h	ad73;
7505	:douta	=	16'h	8c2e;
7506	:douta	=	16'h	ce57;
7507	:douta	=	16'h	18e4;
7508	:douta	=	16'h	8c71;
7509	:douta	=	16'h	4a8c;
7510	:douta	=	16'h	5b50;
7511	:douta	=	16'h	6bf2;
7512	:douta	=	16'h	39c9;
7513	:douta	=	16'h	0841;
7514	:douta	=	16'h	2146;
7515	:douta	=	16'h	3a4d;
7516	:douta	=	16'h	1107;
7517	:douta	=	16'h	29ec;
7518	:douta	=	16'h	328e;
7519	:douta	=	16'h	5bd3;
7520	:douta	=	16'h	328f;
7521	:douta	=	16'h	42af;
7522	:douta	=	16'h	1a0d;
7523	:douta	=	16'h	2a2d;
7524	:douta	=	16'h	4310;
7525	:douta	=	16'h	84d7;
7526	:douta	=	16'h	6477;
7527	:douta	=	16'h	7c56;
7528	:douta	=	16'h	9559;
7529	:douta	=	16'h	5395;
7530	:douta	=	16'h	2a91;
7531	:douta	=	16'h	4333;
7532	:douta	=	16'h	6c56;
7533	:douta	=	16'h	4b53;
7534	:douta	=	16'h	64b8;
7535	:douta	=	16'h	6456;
7536	:douta	=	16'h	9d58;
7537	:douta	=	16'h	6415;
7538	:douta	=	16'h	63d4;
7539	:douta	=	16'h	4352;
7540	:douta	=	16'h	5b30;
7541	:douta	=	16'h	8cd7;
7542	:douta	=	16'h	29ec;
7543	:douta	=	16'h	53b4;
7544	:douta	=	16'h	4312;
7545	:douta	=	16'h	7454;
7546	:douta	=	16'h	6414;
7547	:douta	=	16'h	8495;
7548	:douta	=	16'h	7476;
7549	:douta	=	16'h	4b11;
7550	:douta	=	16'h	a597;
7551	:douta	=	16'h	84b7;
7552	:douta	=	16'h	7475;
7553	:douta	=	16'h	42ef;
7554	:douta	=	16'h	3a4c;
7555	:douta	=	16'h	4af0;
7556	:douta	=	16'h	73f3;
7557	:douta	=	16'h	5b91;
7558	:douta	=	16'h	3a2a;
7559	:douta	=	16'h	3167;
7560	:douta	=	16'h	29a6;
7561	:douta	=	16'h	1946;
7562	:douta	=	16'h	3925;
7563	:douta	=	16'h	72aa;
7564	:douta	=	16'h	9431;
7565	:douta	=	16'h	7c96;
7566	:douta	=	16'h	84f8;
7567	:douta	=	16'h	7477;
7568	:douta	=	16'h	7497;
7569	:douta	=	16'h	7497;
7570	:douta	=	16'h	84f9;
7571	:douta	=	16'h	84f9;
7572	:douta	=	16'h	6c15;
7573	:douta	=	16'h	6415;
7574	:douta	=	16'h	63f5;
7575	:douta	=	16'h	957b;
7576	:douta	=	16'h	adfd;
7577	:douta	=	16'h	853b;
7578	:douta	=	16'h	853a;
7579	:douta	=	16'h	8d3a;
7580	:douta	=	16'h	853a;
7581	:douta	=	16'h	8d7b;
7582	:douta	=	16'h	8d3a;
7583	:douta	=	16'h	8d3a;
7584	:douta	=	16'h	8d5a;
7585	:douta	=	16'h	84f9;
7586	:douta	=	16'h	84f9;
7587	:douta	=	16'h	8d3a;
7588	:douta	=	16'h	84f9;
7589	:douta	=	16'h	853a;
7590	:douta	=	16'h	957b;
7591	:douta	=	16'h	8d7b;
7592	:douta	=	16'h	8d5b;
7593	:douta	=	16'h	957b;
7594	:douta	=	16'h	8d5b;
7595	:douta	=	16'h	853a;
7596	:douta	=	16'h	959b;
7597	:douta	=	16'h	855a;
7598	:douta	=	16'h	853a;
7599	:douta	=	16'h	959b;
7600	:douta	=	16'h	8d5a;
7601	:douta	=	16'h	957b;
7602	:douta	=	16'h	8d9c;
7603	:douta	=	16'h	6cb9;
7604	:douta	=	16'h	6cba;
7605	:douta	=	16'h	751a;
7606	:douta	=	16'h	7d7c;
7607	:douta	=	16'h	53f6;
7608	:douta	=	16'h	32d2;
7609	:douta	=	16'h	7d1b;
7610	:douta	=	16'h	7d5b;
7611	:douta	=	16'h	859c;
7612	:douta	=	16'h	751a;
7613	:douta	=	16'h	7d1a;
7614	:douta	=	16'h	74fa;
7615	:douta	=	16'h	5c37;
7616	:douta	=	16'h	7d3a;
7617	:douta	=	16'h	855b;
7618	:douta	=	16'h	74da;
7619	:douta	=	16'h	7d3a;
7620	:douta	=	16'h	855b;
7621	:douta	=	16'h	855b;
7622	:douta	=	16'h	857b;
7623	:douta	=	16'h	7d3a;
7624	:douta	=	16'h	857b;
7625	:douta	=	16'h	7d3a;
7626	:douta	=	16'h	859b;
7627	:douta	=	16'h	7d1a;
7628	:douta	=	16'h	74d9;
7629	:douta	=	16'h	74d9;
7630	:douta	=	16'h	74d9;
7631	:douta	=	16'h	7d1a;
7632	:douta	=	16'h	6cb9;
7633	:douta	=	16'h	853b;
7634	:douta	=	16'h	855b;
7635	:douta	=	16'h	74da;
7636	:douta	=	16'h	857c;
7637	:douta	=	16'h	6cb9;
7638	:douta	=	16'h	6cb9;
7639	:douta	=	16'h	7d5c;
7640	:douta	=	16'h	751a;
7641	:douta	=	16'h	6c98;
7642	:douta	=	16'h	6cda;
7643	:douta	=	16'h	7d5c;
7644	:douta	=	16'h	6cba;
7645	:douta	=	16'h	6499;
7646	:douta	=	16'h	751a;
7647	:douta	=	16'h	74fa;
7648	:douta	=	16'h	751b;
7649	:douta	=	16'h	6436;
7650	:douta	=	16'h	42af;
7651	:douta	=	16'h	29ca;
7652	:douta	=	16'h	1906;
7653	:douta	=	16'h	08e5;
7654	:douta	=	16'h	1947;
7655	:douta	=	16'h	1927;
7656	:douta	=	16'h	1927;
7657	:douta	=	16'h	2a4e;
7658	:douta	=	16'h	5392;
7659	:douta	=	16'h	4b51;
7660	:douta	=	16'h	63f3;
7661	:douta	=	16'h	84d6;
7662	:douta	=	16'h	8cb5;
7663	:douta	=	16'h	a578;
7664	:douta	=	16'h	5394;
7665	:douta	=	16'h	5bf5;
7666	:douta	=	16'h	2a50;
7667	:douta	=	16'h	2ab0;
7668	:douta	=	16'h	4b73;
7669	:douta	=	16'h	b63b;
7670	:douta	=	16'h	8d7a;
7671	:douta	=	16'h	9579;
7672	:douta	=	16'h	6c78;
7673	:douta	=	16'h	6478;
7674	:douta	=	16'h	2ab1;
7675	:douta	=	16'h	5395;
7676	:douta	=	16'h	4b73;
7677	:douta	=	16'h	6c77;
7678	:douta	=	16'h	b65c;
7679	:douta	=	16'h	6458;
7680	:douta	=	16'h	2a6f;
7681	:douta	=	16'h	2a70;
7682	:douta	=	16'h	19ad;
7683	:douta	=	16'h	42d1;
7684	:douta	=	16'h	32b0;
7685	:douta	=	16'h	32b0;
7686	:douta	=	16'h	5c15;
7687	:douta	=	16'h	63d4;
7688	:douta	=	16'h	63f4;
7689	:douta	=	16'h	6bf5;
7690	:douta	=	16'h	7c96;
7691	:douta	=	16'h	5bb3;
7692	:douta	=	16'h	6b91;
7693	:douta	=	16'h	7c34;
7694	:douta	=	16'h	9517;
7695	:douta	=	16'h	7c74;
7696	:douta	=	16'h	ce38;
7697	:douta	=	16'h	d6bb;
7698	:douta	=	16'h	8474;
7699	:douta	=	16'h	2a70;
7700	:douta	=	16'h	8454;
7701	:douta	=	16'h	8451;
7702	:douta	=	16'h	ad75;
7703	:douta	=	16'h	ad56;
7704	:douta	=	16'h	ce38;
7705	:douta	=	16'h	d638;
7706	:douta	=	16'h	b597;
7707	:douta	=	16'h	8c93;
7708	:douta	=	16'h	63d3;
7709	:douta	=	16'h	ad55;
7710	:douta	=	16'h	bdb6;
7711	:douta	=	16'h	ad95;
7712	:douta	=	16'h	94b4;
7713	:douta	=	16'h	ef3a;
7714	:douta	=	16'h	6bb2;
7715	:douta	=	16'h	94b2;
7716	:douta	=	16'h	8411;
7717	:douta	=	16'h	b595;
7718	:douta	=	16'h	ded8;
7719	:douta	=	16'h	d637;
7720	:douta	=	16'h	ffdb;
7721	:douta	=	16'h	8451;
7722	:douta	=	16'h	9cd3;
7723	:douta	=	16'h	ce36;
7724	:douta	=	16'h	b575;
7725	:douta	=	16'h	b5d6;
7726	:douta	=	16'h	7bd0;
7727	:douta	=	16'h	ce16;
7728	:douta	=	16'h	b533;
7729	:douta	=	16'h	a513;
7730	:douta	=	16'h	9430;
7731	:douta	=	16'h	ad53;
7732	:douta	=	16'h	632d;
7733	:douta	=	16'h	a4f1;
7734	:douta	=	16'h	3a2a;
7735	:douta	=	16'h	8c2e;
7736	:douta	=	16'h	944e;
7737	:douta	=	16'h	c593;
7738	:douta	=	16'h	734b;
7739	:douta	=	16'h	ffba;
7740	:douta	=	16'h	d698;
7741	:douta	=	16'h	cd73;
7742	:douta	=	16'h	b5f4;
7743	:douta	=	16'h	62ec;
7744	:douta	=	16'h	5b4c;
7745	:douta	=	16'h	52ca;
7746	:douta	=	16'h	7c2f;
7747	:douta	=	16'h	4a8a;
7748	:douta	=	16'h	740f;
7749	:douta	=	16'h	5aaa;
7750	:douta	=	16'h	4a28;
7751	:douta	=	16'h	6bf0;
7752	:douta	=	16'h	426b;
7753	:douta	=	16'h	a573;
7754	:douta	=	16'h	7bcf;
7755	:douta	=	16'h	ce76;
7756	:douta	=	16'h	8c30;
7757	:douta	=	16'h	c5d5;
7758	:douta	=	16'h	634e;
7759	:douta	=	16'h	840f;
7760	:douta	=	16'h	73cf;
7761	:douta	=	16'h	528a;
7762	:douta	=	16'h	8c4f;
7763	:douta	=	16'h	2945;
7764	:douta	=	16'h	63d1;
7765	:douta	=	16'h	5b50;
7766	:douta	=	16'h	4aef;
7767	:douta	=	16'h	63d2;
7768	:douta	=	16'h	0881;
7769	:douta	=	16'h	0841;
7770	:douta	=	16'h	0840;
7771	:douta	=	16'h	2147;
7772	:douta	=	16'h	320b;
7773	:douta	=	16'h	29ab;
7774	:douta	=	16'h	3a8f;
7775	:douta	=	16'h	2a4d;
7776	:douta	=	16'h	3ab0;
7777	:douta	=	16'h	5392;
7778	:douta	=	16'h	328f;
7779	:douta	=	16'h	5371;
7780	:douta	=	16'h	2a4e;
7781	:douta	=	16'h	63f4;
7782	:douta	=	16'h	32b0;
7783	:douta	=	16'h	63f4;
7784	:douta	=	16'h	8d38;
7785	:douta	=	16'h	6cb8;
7786	:douta	=	16'h	3b34;
7787	:douta	=	16'h	5bd4;
7788	:douta	=	16'h	7497;
7789	:douta	=	16'h	6c77;
7790	:douta	=	16'h	3b11;
7791	:douta	=	16'h	5352;
7792	:douta	=	16'h	84d6;
7793	:douta	=	16'h	6415;
7794	:douta	=	16'h	7c96;
7795	:douta	=	16'h	6436;
7796	:douta	=	16'h	9d16;
7797	:douta	=	16'h	a61c;
7798	:douta	=	16'h	5b93;
7799	:douta	=	16'h	5bd4;
7800	:douta	=	16'h	4b31;
7801	:douta	=	16'h	5393;
7802	:douta	=	16'h	324e;
7803	:douta	=	16'h	42ef;
7804	:douta	=	16'h	21ec;
7805	:douta	=	16'h	5372;
7806	:douta	=	16'h	8cd5;
7807	:douta	=	16'h	6bf4;
7808	:douta	=	16'h	8d59;
7809	:douta	=	16'h	5bd4;
7810	:douta	=	16'h	8433;
7811	:douta	=	16'h	7433;
7812	:douta	=	16'h	6c13;
7813	:douta	=	16'h	3187;
7814	:douta	=	16'h	2945;
7815	:douta	=	16'h	31a7;
7816	:douta	=	16'h	10e5;
7817	:douta	=	16'h	2905;
7818	:douta	=	16'h	8b8d;
7819	:douta	=	16'h	9452;
7820	:douta	=	16'h	7c76;
7821	:douta	=	16'h	7cd7;
7822	:douta	=	16'h	84d8;
7823	:douta	=	16'h	7c98;
7824	:douta	=	16'h	7497;
7825	:douta	=	16'h	7cb8;
7826	:douta	=	16'h	7c98;
7827	:douta	=	16'h	7477;
7828	:douta	=	16'h	8d5a;
7829	:douta	=	16'h	84f9;
7830	:douta	=	16'h	63f5;
7831	:douta	=	16'h	63f6;
7832	:douta	=	16'h	7cd9;
7833	:douta	=	16'h	a61d;
7834	:douta	=	16'h	9dbc;
7835	:douta	=	16'h	959c;
7836	:douta	=	16'h	853a;
7837	:douta	=	16'h	851a;
7838	:douta	=	16'h	8d5a;
7839	:douta	=	16'h	8d5a;
7840	:douta	=	16'h	8519;
7841	:douta	=	16'h	7cd9;
7842	:douta	=	16'h	7cf9;
7843	:douta	=	16'h	8d7b;
7844	:douta	=	16'h	853a;
7845	:douta	=	16'h	851a;
7846	:douta	=	16'h	8d5b;
7847	:douta	=	16'h	8d9b;
7848	:douta	=	16'h	851a;
7849	:douta	=	16'h	8d5a;
7850	:douta	=	16'h	95bc;
7851	:douta	=	16'h	95bc;
7852	:douta	=	16'h	957b;
7853	:douta	=	16'h	8d5b;
7854	:douta	=	16'h	8d5b;
7855	:douta	=	16'h	8d5b;
7856	:douta	=	16'h	8d5b;
7857	:douta	=	16'h	8d7b;
7858	:douta	=	16'h	8d7b;
7859	:douta	=	16'h	8d9b;
7860	:douta	=	16'h	6cba;
7861	:douta	=	16'h	6499;
7862	:douta	=	16'h	6478;
7863	:douta	=	16'h	8dbd;
7864	:douta	=	16'h	859c;
7865	:douta	=	16'h	5c38;
7866	:douta	=	16'h	6cba;
7867	:douta	=	16'h	74fa;
7868	:douta	=	16'h	7d5b;
7869	:douta	=	16'h	7d3a;
7870	:douta	=	16'h	7d1a;
7871	:douta	=	16'h	74f9;
7872	:douta	=	16'h	6cb9;
7873	:douta	=	16'h	857b;
7874	:douta	=	16'h	8d9c;
7875	:douta	=	16'h	6cb9;
7876	:douta	=	16'h	6c99;
7877	:douta	=	16'h	859b;
7878	:douta	=	16'h	7d5b;
7879	:douta	=	16'h	74d9;
7880	:douta	=	16'h	855b;
7881	:douta	=	16'h	7d5b;
7882	:douta	=	16'h	8d9b;
7883	:douta	=	16'h	74d9;
7884	:douta	=	16'h	855b;
7885	:douta	=	16'h	8d9b;
7886	:douta	=	16'h	7d3a;
7887	:douta	=	16'h	7d1a;
7888	:douta	=	16'h	74fa;
7889	:douta	=	16'h	74fa;
7890	:douta	=	16'h	857b;
7891	:douta	=	16'h	857b;
7892	:douta	=	16'h	6cb9;
7893	:douta	=	16'h	7d5b;
7894	:douta	=	16'h	753a;
7895	:douta	=	16'h	857b;
7896	:douta	=	16'h	7d3b;
7897	:douta	=	16'h	7d5b;
7898	:douta	=	16'h	6c78;
7899	:douta	=	16'h	6cd9;
7900	:douta	=	16'h	6cb9;
7901	:douta	=	16'h	6cb9;
7902	:douta	=	16'h	6cb9;
7903	:douta	=	16'h	74fa;
7904	:douta	=	16'h	753b;
7905	:douta	=	16'h	74fa;
7906	:douta	=	16'h	6cba;
7907	:douta	=	16'h	3a4c;
7908	:douta	=	16'h	2168;
7909	:douta	=	16'h	2188;
7910	:douta	=	16'h	1106;
7911	:douta	=	16'h	1127;
7912	:douta	=	16'h	1127;
7913	:douta	=	16'h	218a;
7914	:douta	=	16'h	7456;
7915	:douta	=	16'h	4332;
7916	:douta	=	16'h	5393;
7917	:douta	=	16'h	4b10;
7918	:douta	=	16'h	9d16;
7919	:douta	=	16'h	b5da;
7920	:douta	=	16'h	9539;
7921	:douta	=	16'h	ae1c;
7922	:douta	=	16'h	4b53;
7923	:douta	=	16'h	2a90;
7924	:douta	=	16'h	222f;
7925	:douta	=	16'h	32d1;
7926	:douta	=	16'h	2ab0;
7927	:douta	=	16'h	7497;
7928	:douta	=	16'h	959b;
7929	:douta	=	16'h	957a;
7930	:douta	=	16'h	4b75;
7931	:douta	=	16'h	5bd4;
7932	:douta	=	16'h	3b12;
7933	:douta	=	16'h	6c77;
7934	:douta	=	16'h	53d4;
7935	:douta	=	16'h	4b94;
7936	:douta	=	16'h	32f2;
7937	:douta	=	16'h	5416;
7938	:douta	=	16'h	53d5;
7939	:douta	=	16'h	7457;
7940	:douta	=	16'h	6477;
7941	:douta	=	16'h	6416;
7942	:douta	=	16'h	4373;
7943	:douta	=	16'h	5373;
7944	:douta	=	16'h	198b;
7945	:douta	=	16'h	5372;
7946	:douta	=	16'h	6c14;
7947	:douta	=	16'h	7455;
7948	:douta	=	16'h	94d6;
7949	:douta	=	16'h	a599;
7950	:douta	=	16'h	8454;
7951	:douta	=	16'h	73f3;
7952	:douta	=	16'h	8473;
7953	:douta	=	16'h	8494;
7954	:douta	=	16'h	7c12;
7955	:douta	=	16'h	9d56;
7956	:douta	=	16'h	bdd8;
7957	:douta	=	16'h	b597;
7958	:douta	=	16'h	8c94;
7959	:douta	=	16'h	a557;
7960	:douta	=	16'h	9cb5;
7961	:douta	=	16'h	ce58;
7962	:douta	=	16'h	9d15;
7963	:douta	=	16'h	c5f7;
7964	:douta	=	16'h	a556;
7965	:douta	=	16'h	ce17;
7966	:douta	=	16'h	9cd4;
7967	:douta	=	16'h	b575;
7968	:douta	=	16'h	8cb3;
7969	:douta	=	16'h	a4d4;
7970	:douta	=	16'h	ad55;
7971	:douta	=	16'h	bdb5;
7972	:douta	=	16'h	de98;
7973	:douta	=	16'h	ce57;
7974	:douta	=	16'h	8474;
7975	:douta	=	16'h	de98;
7976	:douta	=	16'h	8c72;
7977	:douta	=	16'h	b532;
7978	:douta	=	16'h	a514;
7979	:douta	=	16'h	73f0;
7980	:douta	=	16'h	ce15;
7981	:douta	=	16'h	de98;
7982	:douta	=	16'h	cdf5;
7983	:douta	=	16'h	ef19;
7984	:douta	=	16'h	acd1;
7985	:douta	=	16'h	426a;
7986	:douta	=	16'h	5acb;
7987	:douta	=	16'h	d655;
7988	:douta	=	16'h	acf1;
7989	:douta	=	16'h	e6d7;
7990	:douta	=	16'h	ac8f;
7991	:douta	=	16'h	ff38;
7992	:douta	=	16'h	5289;
7993	:douta	=	16'h	6aca;
7994	:douta	=	16'h	8410;
7995	:douta	=	16'h	b510;
7996	:douta	=	16'h	ad92;
7997	:douta	=	16'h	946f;
7998	:douta	=	16'h	7bcd;
7999	:douta	=	16'h	62cb;
8000	:douta	=	16'h	10e4;
8001	:douta	=	16'h	2127;
8002	:douta	=	16'h	1926;
8003	:douta	=	16'h	18e5;
8004	:douta	=	16'h	1905;
8005	:douta	=	16'h	0043;
8006	:douta	=	16'h	736d;
8007	:douta	=	16'h	73ae;
8008	:douta	=	16'h	9c91;
8009	:douta	=	16'h	7410;
8010	:douta	=	16'h	c5b5;
8011	:douta	=	16'h	ad32;
8012	:douta	=	16'h	31ea;
8013	:douta	=	16'h	8c50;
8014	:douta	=	16'h	4a8c;
8015	:douta	=	16'h	9cb0;
8016	:douta	=	16'h	8470;
8017	:douta	=	16'h	de97;
8018	:douta	=	16'h	a574;
8019	:douta	=	16'h	5b4e;
8020	:douta	=	16'h	3a6e;
8021	:douta	=	16'h	63d3;
8022	:douta	=	16'h	4aae;
8023	:douta	=	16'h	4a4b;
8024	:douta	=	16'h	0840;
8025	:douta	=	16'h	18a2;
8026	:douta	=	16'h	1083;
8027	:douta	=	16'h	1082;
8028	:douta	=	16'h	0860;
8029	:douta	=	16'h	1882;
8030	:douta	=	16'h	2967;
8031	:douta	=	16'h	3aaf;
8032	:douta	=	16'h	0108;
8033	:douta	=	16'h	0907;
8034	:douta	=	16'h	2a2c;
8035	:douta	=	16'h	5393;
8036	:douta	=	16'h	322d;
8037	:douta	=	16'h	6477;
8038	:douta	=	16'h	3b73;
8039	:douta	=	16'h	6c56;
8040	:douta	=	16'h	5393;
8041	:douta	=	16'h	5b93;
8042	:douta	=	16'h	42f1;
8043	:douta	=	16'h	4b53;
8044	:douta	=	16'h	6436;
8045	:douta	=	16'h	63f5;
8046	:douta	=	16'h	5c37;
8047	:douta	=	16'h	6bf2;
8048	:douta	=	16'h	9dba;
8049	:douta	=	16'h	4acf;
8050	:douta	=	16'h	6c35;
8051	:douta	=	16'h	5352;
8052	:douta	=	16'h	6bf5;
8053	:douta	=	16'h	42f1;
8054	:douta	=	16'h	4b94;
8055	:douta	=	16'h	32b1;
8056	:douta	=	16'h	7c56;
8057	:douta	=	16'h	6c56;
8058	:douta	=	16'h	6c15;
8059	:douta	=	16'h	63d3;
8060	:douta	=	16'h	6414;
8061	:douta	=	16'h	9d57;
8062	:douta	=	16'h	63d3;
8063	:douta	=	16'h	a599;
8064	:douta	=	16'h	42ef;
8065	:douta	=	16'h	7413;
8066	:douta	=	16'h	42ae;
8067	:douta	=	16'h	4aad;
8068	:douta	=	16'h	3147;
8069	:douta	=	16'h	31c7;
8070	:douta	=	16'h	2988;
8071	:douta	=	16'h	41a6;
8072	:douta	=	16'h	9bee;
8073	:douta	=	16'h	8c52;
8074	:douta	=	16'h	7477;
8075	:douta	=	16'h	84f8;
8076	:douta	=	16'h	7cb7;
8077	:douta	=	16'h	84f8;
8078	:douta	=	16'h	84f8;
8079	:douta	=	16'h	7c97;
8080	:douta	=	16'h	7c97;
8081	:douta	=	16'h	8d39;
8082	:douta	=	16'h	7cb8;
8083	:douta	=	16'h	84f9;
8084	:douta	=	16'h	84d8;
8085	:douta	=	16'h	7cb8;
8086	:douta	=	16'h	6c36;
8087	:douta	=	16'h	84f9;
8088	:douta	=	16'h	7cd8;
8089	:douta	=	16'h	5373;
8090	:douta	=	16'h	4b12;
8091	:douta	=	16'h	8d7b;
8092	:douta	=	16'h	957b;
8093	:douta	=	16'h	959b;
8094	:douta	=	16'h	9dbc;
8095	:douta	=	16'h	8d5a;
8096	:douta	=	16'h	851a;
8097	:douta	=	16'h	7477;
8098	:douta	=	16'h	6c36;
8099	:douta	=	16'h	84d9;
8100	:douta	=	16'h	84d9;
8101	:douta	=	16'h	959b;
8102	:douta	=	16'h	8d3a;
8103	:douta	=	16'h	8d5b;
8104	:douta	=	16'h	851a;
8105	:douta	=	16'h	853a;
8106	:douta	=	16'h	851a;
8107	:douta	=	16'h	74b8;
8108	:douta	=	16'h	8d5a;
8109	:douta	=	16'h	8d7b;
8110	:douta	=	16'h	959b;
8111	:douta	=	16'h	957b;
8112	:douta	=	16'h	957b;
8113	:douta	=	16'h	8d7b;
8114	:douta	=	16'h	959c;
8115	:douta	=	16'h	95bc;
8116	:douta	=	16'h	95bc;
8117	:douta	=	16'h	959c;
8118	:douta	=	16'h	6c98;
8119	:douta	=	16'h	74da;
8120	:douta	=	16'h	6c99;
8121	:douta	=	16'h	5c58;
8122	:douta	=	16'h	6cb9;
8123	:douta	=	16'h	859c;
8124	:douta	=	16'h	4b75;
8125	:douta	=	16'h	4b76;
8126	:douta	=	16'h	857c;
8127	:douta	=	16'h	8dbc;
8128	:douta	=	16'h	7d3b;
8129	:douta	=	16'h	74da;
8130	:douta	=	16'h	74d9;
8131	:douta	=	16'h	855b;
8132	:douta	=	16'h	9e3e;
8133	:douta	=	16'h	7d3a;
8134	:douta	=	16'h	6cb9;
8135	:douta	=	16'h	859c;
8136	:douta	=	16'h	855b;
8137	:douta	=	16'h	855b;
8138	:douta	=	16'h	7d5b;
8139	:douta	=	16'h	7d3b;
8140	:douta	=	16'h	7d5b;
8141	:douta	=	16'h	5c17;
8142	:douta	=	16'h	6478;
8143	:douta	=	16'h	8d9b;
8144	:douta	=	16'h	7d3a;
8145	:douta	=	16'h	7d3a;
8146	:douta	=	16'h	855b;
8147	:douta	=	16'h	7d3a;
8148	:douta	=	16'h	7d3b;
8149	:douta	=	16'h	7d3b;
8150	:douta	=	16'h	7d5b;
8151	:douta	=	16'h	753a;
8152	:douta	=	16'h	8dbc;
8153	:douta	=	16'h	8d9b;
8154	:douta	=	16'h	7d7b;
8155	:douta	=	16'h	7d7c;
8156	:douta	=	16'h	6cba;
8157	:douta	=	16'h	6458;
8158	:douta	=	16'h	7d3a;
8159	:douta	=	16'h	74fa;
8160	:douta	=	16'h	74da;
8161	:douta	=	16'h	6d1a;
8162	:douta	=	16'h	755b;
8163	:douta	=	16'h	753b;
8164	:douta	=	16'h	74b8;
8165	:douta	=	16'h	42cf;
8166	:douta	=	16'h	21a8;
8167	:douta	=	16'h	21a8;
8168	:douta	=	16'h	1107;
8169	:douta	=	16'h	1927;
8170	:douta	=	16'h	1107;
8171	:douta	=	16'h	32af;
8172	:douta	=	16'h	8518;
8173	:douta	=	16'h	8c94;
8174	:douta	=	16'h	7455;
8175	:douta	=	16'h	63f5;
8176	:douta	=	16'h	1a0e;
8177	:douta	=	16'h	3ab0;
8178	:douta	=	16'h	5373;
8179	:douta	=	16'h	addb;
8180	:douta	=	16'h	adfc;
8181	:douta	=	16'h	63d4;
8182	:douta	=	16'h	957a;
8183	:douta	=	16'h	2a90;
8184	:douta	=	16'h	2a70;
8185	:douta	=	16'h	4395;
8186	:douta	=	16'h	5bb3;
8187	:douta	=	16'h	8518;
8188	:douta	=	16'h	be3b;
8189	:douta	=	16'h	9dbb;
8190	:douta	=	16'h	6416;
8191	:douta	=	16'h	8d5a;
8192	:douta	=	16'h	2a4f;
8193	:douta	=	16'h	2250;
8194	:douta	=	16'h	1a0e;
8195	:douta	=	16'h	5374;
8196	:douta	=	16'h	74b9;
8197	:douta	=	16'h	6c77;
8198	:douta	=	16'h	6437;
8199	:douta	=	16'h	4b53;
8200	:douta	=	16'h	3a8e;
8201	:douta	=	16'h	5352;
8202	:douta	=	16'h	2a2e;
8203	:douta	=	16'h	42f2;
8204	:douta	=	16'h	8475;
8205	:douta	=	16'h	6350;
8206	:douta	=	16'h	ad97;
8207	:douta	=	16'h	8cb5;
8208	:douta	=	16'h	9453;
8209	:douta	=	16'h	ce39;
8210	:douta	=	16'h	8c75;
8211	:douta	=	16'h	63f4;
8212	:douta	=	16'h	9d15;
8213	:douta	=	16'h	94b4;
8214	:douta	=	16'h	ad36;
8215	:douta	=	16'h	bdf8;
8216	:douta	=	16'h	bdb7;
8217	:douta	=	16'h	ce38;
8218	:douta	=	16'h	6bf3;
8219	:douta	=	16'h	8412;
8220	:douta	=	16'h	5bb1;
8221	:douta	=	16'h	b596;
8222	:douta	=	16'h	c5f7;
8223	:douta	=	16'h	de98;
8224	:douta	=	16'h	bdb6;
8225	:douta	=	16'h	c617;
8226	:douta	=	16'h	7c33;
8227	:douta	=	16'h	94d4;
8228	:douta	=	16'h	8432;
8229	:douta	=	16'h	d657;
8230	:douta	=	16'h	de98;
8231	:douta	=	16'h	e6d9;
8232	:douta	=	16'h	bdb5;
8233	:douta	=	16'h	e6d8;
8234	:douta	=	16'h	b595;
8235	:douta	=	16'h	94d3;
8236	:douta	=	16'h	ad13;
8237	:douta	=	16'h	8cb3;
8238	:douta	=	16'h	d655;
8239	:douta	=	16'h	d677;
8240	:douta	=	16'h	de55;
8241	:douta	=	16'h	a4b0;
8242	:douta	=	16'h	9430;
8243	:douta	=	16'h	bdd3;
8244	:douta	=	16'h	52ac;
8245	:douta	=	16'h	bdd4;
8246	:douta	=	16'h	9c8e;
8247	:douta	=	16'h	b551;
8248	:douta	=	16'h	8bcc;
8249	:douta	=	16'h	cdf4;
8250	:douta	=	16'h	6b4c;
8251	:douta	=	16'h	f779;
8252	:douta	=	16'h	9d12;
8253	:douta	=	16'h	5a8a;
8254	:douta	=	16'h	41c7;
8255	:douta	=	16'h	2967;
8256	:douta	=	16'h	2967;
8257	:douta	=	16'h	2126;
8258	:douta	=	16'h	2126;
8259	:douta	=	16'h	1926;
8260	:douta	=	16'h	1925;
8261	:douta	=	16'h	10e5;
8262	:douta	=	16'h	0042;
8263	:douta	=	16'h	3a4b;
8264	:douta	=	16'h	738e;
8265	:douta	=	16'h	9cd2;
8266	:douta	=	16'h	9450;
8267	:douta	=	16'h	ad53;
8268	:douta	=	16'h	9430;
8269	:douta	=	16'h	bd74;
8270	:douta	=	16'h	42ac;
8271	:douta	=	16'h	83ee;
8272	:douta	=	16'h	5b2c;
8273	:douta	=	16'h	83ee;
8274	:douta	=	16'h	9cf2;
8275	:douta	=	16'h	63f3;
8276	:douta	=	16'h	29eb;
8277	:douta	=	16'h	5b71;
8278	:douta	=	16'h	5bb1;
8279	:douta	=	16'h	5350;
8280	:douta	=	16'h	4a8b;
8281	:douta	=	16'h	18a2;
8282	:douta	=	16'h	1883;
8283	:douta	=	16'h	18a2;
8284	:douta	=	16'h	18a3;
8285	:douta	=	16'h	1020;
8286	:douta	=	16'h	0800;
8287	:douta	=	16'h	320b;
8288	:douta	=	16'h	21ea;
8289	:douta	=	16'h	08e6;
8290	:douta	=	16'h	21aa;
8291	:douta	=	16'h	3af0;
8292	:douta	=	16'h	4bb3;
8293	:douta	=	16'h	2a8f;
8294	:douta	=	16'h	19ac;
8295	:douta	=	16'h	6435;
8296	:douta	=	16'h	4b93;
8297	:douta	=	16'h	5c16;
8298	:douta	=	16'h	7476;
8299	:douta	=	16'h	8559;
8300	:douta	=	16'h	5373;
8301	:douta	=	16'h	5c15;
8302	:douta	=	16'h	2a6f;
8303	:douta	=	16'h	84d6;
8304	:douta	=	16'h	7d19;
8305	:douta	=	16'h	84d6;
8306	:douta	=	16'h	6477;
8307	:douta	=	16'h	74b7;
8308	:douta	=	16'h	9d9a;
8309	:douta	=	16'h	5bf5;
8310	:douta	=	16'h	5394;
8311	:douta	=	16'h	3b12;
8312	:douta	=	16'h	8475;
8313	:douta	=	16'h	4b52;
8314	:douta	=	16'h	5311;
8315	:douta	=	16'h	3aaf;
8316	:douta	=	16'h	6c35;
8317	:douta	=	16'h	7c96;
8318	:douta	=	16'h	6bf4;
8319	:douta	=	16'h	a5b9;
8320	:douta	=	16'h	4b31;
8321	:douta	=	16'h	5b71;
8322	:douta	=	16'h	428d;
8323	:douta	=	16'h	3168;
8324	:douta	=	16'h	39a8;
8325	:douta	=	16'h	2147;
8326	:douta	=	16'h	20e5;
8327	:douta	=	16'h	a40e;
8328	:douta	=	16'h	6bb3;
8329	:douta	=	16'h	7c54;
8330	:douta	=	16'h	8518;
8331	:douta	=	16'h	7c97;
8332	:douta	=	16'h	7456;
8333	:douta	=	16'h	6c35;
8334	:douta	=	16'h	7c97;
8335	:douta	=	16'h	8d18;
8336	:douta	=	16'h	84f8;
8337	:douta	=	16'h	7c76;
8338	:douta	=	16'h	8519;
8339	:douta	=	16'h	7cb7;
8340	:douta	=	16'h	84f8;
8341	:douta	=	16'h	84f9;
8342	:douta	=	16'h	7c97;
8343	:douta	=	16'h	8519;
8344	:douta	=	16'h	74b8;
8345	:douta	=	16'h	8d1a;
8346	:douta	=	16'h	7477;
8347	:douta	=	16'h	4b74;
8348	:douta	=	16'h	84f9;
8349	:douta	=	16'h	851a;
8350	:douta	=	16'h	851a;
8351	:douta	=	16'h	957b;
8352	:douta	=	16'h	8519;
8353	:douta	=	16'h	7cb9;
8354	:douta	=	16'h	7497;
8355	:douta	=	16'h	8d5a;
8356	:douta	=	16'h	7cb8;
8357	:douta	=	16'h	851a;
8358	:douta	=	16'h	95bc;
8359	:douta	=	16'h	9dbc;
8360	:douta	=	16'h	957b;
8361	:douta	=	16'h	8d5a;
8362	:douta	=	16'h	8d5b;
8363	:douta	=	16'h	8d3a;
8364	:douta	=	16'h	8d5a;
8365	:douta	=	16'h	8d5b;
8366	:douta	=	16'h	8d5b;
8367	:douta	=	16'h	95bc;
8368	:douta	=	16'h	95bc;
8369	:douta	=	16'h	959b;
8370	:douta	=	16'h	853a;
8371	:douta	=	16'h	8d7b;
8372	:douta	=	16'h	9dbc;
8373	:douta	=	16'h	9dbc;
8374	:douta	=	16'h	95bc;
8375	:douta	=	16'h	6cb9;
8376	:douta	=	16'h	6c58;
8377	:douta	=	16'h	5395;
8378	:douta	=	16'h	4353;
8379	:douta	=	16'h	6498;
8380	:douta	=	16'h	753b;
8381	:douta	=	16'h	5c38;
8382	:douta	=	16'h	53f7;
8383	:douta	=	16'h	74da;
8384	:douta	=	16'h	857c;
8385	:douta	=	16'h	6cda;
8386	:douta	=	16'h	7d3b;
8387	:douta	=	16'h	74da;
8388	:douta	=	16'h	74fa;
8389	:douta	=	16'h	95bc;
8390	:douta	=	16'h	7d3b;
8391	:douta	=	16'h	74da;
8392	:douta	=	16'h	74d9;
8393	:douta	=	16'h	74da;
8394	:douta	=	16'h	859c;
8395	:douta	=	16'h	857b;
8396	:douta	=	16'h	7d5b;
8397	:douta	=	16'h	6478;
8398	:douta	=	16'h	74fa;
8399	:douta	=	16'h	74d9;
8400	:douta	=	16'h	8d9b;
8401	:douta	=	16'h	8d9b;
8402	:douta	=	16'h	6cd9;
8403	:douta	=	16'h	7d3b;
8404	:douta	=	16'h	74da;
8405	:douta	=	16'h	6cba;
8406	:douta	=	16'h	753a;
8407	:douta	=	16'h	7d3b;
8408	:douta	=	16'h	857b;
8409	:douta	=	16'h	7d1a;
8410	:douta	=	16'h	8dbc;
8411	:douta	=	16'h	95dc;
8412	:douta	=	16'h	855b;
8413	:douta	=	16'h	7d1a;
8414	:douta	=	16'h	6c99;
8415	:douta	=	16'h	857c;
8416	:douta	=	16'h	753b;
8417	:douta	=	16'h	6c99;
8418	:douta	=	16'h	6cda;
8419	:douta	=	16'h	753b;
8420	:douta	=	16'h	74b9;
8421	:douta	=	16'h	7cd8;
8422	:douta	=	16'h	29e9;
8423	:douta	=	16'h	2147;
8424	:douta	=	16'h	1968;
8425	:douta	=	16'h	1148;
8426	:douta	=	16'h	1148;
8427	:douta	=	16'h	08c6;
8428	:douta	=	16'h	21eb;
8429	:douta	=	16'h	7454;
8430	:douta	=	16'h	84d7;
8431	:douta	=	16'h	8539;
8432	:douta	=	16'h	63f5;
8433	:douta	=	16'h	7435;
8434	:douta	=	16'h	222f;
8435	:douta	=	16'h	53d4;
8436	:douta	=	16'h	5bf5;
8437	:douta	=	16'h	b63b;
8438	:douta	=	16'h	955a;
8439	:douta	=	16'h	84d7;
8440	:douta	=	16'h	5c16;
8441	:douta	=	16'h	4353;
8442	:douta	=	16'h	2ab1;
8443	:douta	=	16'h	3b32;
8444	:douta	=	16'h	a5da;
8445	:douta	=	16'h	6416;
8446	:douta	=	16'h	8d39;
8447	:douta	=	16'h	7cf9;
8448	:douta	=	16'h	2ab1;
8449	:douta	=	16'h	53f6;
8450	:douta	=	16'h	6498;
8451	:douta	=	16'h	5374;
8452	:douta	=	16'h	6cb8;
8453	:douta	=	16'h	5bb4;
8454	:douta	=	16'h	5394;
8455	:douta	=	16'h	6436;
8456	:douta	=	16'h	5332;
8457	:douta	=	16'h	5b93;
8458	:douta	=	16'h	9559;
8459	:douta	=	16'h	7c76;
8460	:douta	=	16'h	7414;
8461	:douta	=	16'h	c5f9;
8462	:douta	=	16'h	8c95;
8463	:douta	=	16'h	7c74;
8464	:douta	=	16'h	73f2;
8465	:douta	=	16'h	6bd2;
8466	:douta	=	16'h	9d15;
8467	:douta	=	16'h	73f3;
8468	:douta	=	16'h	ad97;
8469	:douta	=	16'h	a4d4;
8470	:douta	=	16'h	ad35;
8471	:douta	=	16'h	a4f5;
8472	:douta	=	16'h	52ce;
8473	:douta	=	16'h	b596;
8474	:douta	=	16'h	9cd4;
8475	:douta	=	16'h	bdb6;
8476	:douta	=	16'h	b575;
8477	:douta	=	16'h	eef9;
8478	:douta	=	16'h	b5b6;
8479	:douta	=	16'h	a4d3;
8480	:douta	=	16'h	8473;
8481	:douta	=	16'h	a4d3;
8482	:douta	=	16'h	ad75;
8483	:douta	=	16'h	de98;
8484	:douta	=	16'h	9cd4;
8485	:douta	=	16'h	cdf6;
8486	:douta	=	16'h	bdd6;
8487	:douta	=	16'h	d637;
8488	:douta	=	16'h	b575;
8489	:douta	=	16'h	a4d2;
8490	:douta	=	16'h	7bce;
8491	:douta	=	16'h	c5d4;
8492	:douta	=	16'h	e719;
8493	:douta	=	16'h	9cd1;
8494	:douta	=	16'h	e6b7;
8495	:douta	=	16'h	d696;
8496	:douta	=	16'h	9c71;
8497	:douta	=	16'h	634d;
8498	:douta	=	16'h	bd93;
8499	:douta	=	16'h	b593;
8500	:douta	=	16'h	bd92;
8501	:douta	=	16'h	bdd3;
8502	:douta	=	16'h	bd32;
8503	:douta	=	16'h	eeb7;
8504	:douta	=	16'h	31a6;
8505	:douta	=	16'h	7b4b;
8506	:douta	=	16'h	6b4d;
8507	:douta	=	16'h	6b0b;
8508	:douta	=	16'h	6aeb;
8509	:douta	=	16'h	5289;
8510	:douta	=	16'h	5a89;
8511	:douta	=	16'h	4a29;
8512	:douta	=	16'h	3a08;
8513	:douta	=	16'h	18e5;
8514	:douta	=	16'h	2146;
8515	:douta	=	16'h	2146;
8516	:douta	=	16'h	18e5;
8517	:douta	=	16'h	10e4;
8518	:douta	=	16'h	18e5;
8519	:douta	=	16'h	1043;
8520	:douta	=	16'h	bd11;
8521	:douta	=	16'h	5b0e;
8522	:douta	=	16'h	e695;
8523	:douta	=	16'h	a513;
8524	:douta	=	16'h	31c9;
8525	:douta	=	16'h	9450;
8526	:douta	=	16'h	2986;
8527	:douta	=	16'h	bdf5;
8528	:douta	=	16'h	428a;
8529	:douta	=	16'h	8c50;
8530	:douta	=	16'h	42cd;
8531	:douta	=	16'h	4b10;
8532	:douta	=	16'h	5b91;
8533	:douta	=	16'h	428d;
8534	:douta	=	16'h	328d;
8535	:douta	=	16'h	52ee;
8536	:douta	=	16'h	63d2;
8537	:douta	=	16'h	3b11;
8538	:douta	=	16'h	8c51;
8539	:douta	=	16'h	0000;
8540	:douta	=	16'h	1081;
8541	:douta	=	16'h	18e3;
8542	:douta	=	16'h	20e3;
8543	:douta	=	16'h	10c2;
8544	:douta	=	16'h	1082;
8545	:douta	=	16'h	29a8;
8546	:douta	=	16'h	3a2b;
8547	:douta	=	16'h	1127;
8548	:douta	=	16'h	32d0;
8549	:douta	=	16'h	32f0;
8550	:douta	=	16'h	4b72;
8551	:douta	=	16'h	53b4;
8552	:douta	=	16'h	5393;
8553	:douta	=	16'h	19cc;
8554	:douta	=	16'h	5bd4;
8555	:douta	=	16'h	53b4;
8556	:douta	=	16'h	4311;
8557	:douta	=	16'h	42f1;
8558	:douta	=	16'h	6c56;
8559	:douta	=	16'h	7d19;
8560	:douta	=	16'h	4332;
8561	:douta	=	16'h	5c14;
8562	:douta	=	16'h	32af;
8563	:douta	=	16'h	426d;
8564	:douta	=	16'h	3b32;
8565	:douta	=	16'h	4b53;
8566	:douta	=	16'h	3b33;
8567	:douta	=	16'h	4b53;
8568	:douta	=	16'h	8d7a;
8569	:douta	=	16'h	7c97;
8570	:douta	=	16'h	8d38;
8571	:douta	=	16'h	4b31;
8572	:douta	=	16'h	4af0;
8573	:douta	=	16'h	6c34;
8574	:douta	=	16'h	7c75;
8575	:douta	=	16'h	3a8f;
8576	:douta	=	16'h	63d3;
8577	:douta	=	16'h	4aac;
8578	:douta	=	16'h	39c7;
8579	:douta	=	16'h	29a8;
8580	:douta	=	16'h	1926;
8581	:douta	=	16'h	ac0e;
8582	:douta	=	16'h	838d;
8583	:douta	=	16'h	94f7;
8584	:douta	=	16'h	7c76;
8585	:douta	=	16'h	8d19;
8586	:douta	=	16'h	63f4;
8587	:douta	=	16'h	6c15;
8588	:douta	=	16'h	7c76;
8589	:douta	=	16'h	84b7;
8590	:douta	=	16'h	63d3;
8591	:douta	=	16'h	6c15;
8592	:douta	=	16'h	7477;
8593	:douta	=	16'h	8d39;
8594	:douta	=	16'h	8d19;
8595	:douta	=	16'h	957a;
8596	:douta	=	16'h	8d39;
8597	:douta	=	16'h	8d5a;
8598	:douta	=	16'h	8d5a;
8599	:douta	=	16'h	7cd8;
8600	:douta	=	16'h	8519;
8601	:douta	=	16'h	8d3a;
8602	:douta	=	16'h	8d5a;
8603	:douta	=	16'h	84d8;
8604	:douta	=	16'h	8519;
8605	:douta	=	16'h	7477;
8606	:douta	=	16'h	8d3a;
8607	:douta	=	16'h	957b;
8608	:douta	=	16'h	95bc;
8609	:douta	=	16'h	853a;
8610	:douta	=	16'h	8d3a;
8611	:douta	=	16'h	7cb8;
8612	:douta	=	16'h	6c36;
8613	:douta	=	16'h	8d5b;
8614	:douta	=	16'h	853a;
8615	:douta	=	16'h	851a;
8616	:douta	=	16'h	853a;
8617	:douta	=	16'h	855a;
8618	:douta	=	16'h	851a;
8619	:douta	=	16'h	853a;
8620	:douta	=	16'h	959c;
8621	:douta	=	16'h	8d5a;
8622	:douta	=	16'h	853a;
8623	:douta	=	16'h	8d7b;
8624	:douta	=	16'h	8d5a;
8625	:douta	=	16'h	8d5a;
8626	:douta	=	16'h	8d5a;
8627	:douta	=	16'h	8d7b;
8628	:douta	=	16'h	8d7b;
8629	:douta	=	16'h	8d3a;
8630	:douta	=	16'h	8d5a;
8631	:douta	=	16'h	8d9b;
8632	:douta	=	16'h	95bc;
8633	:douta	=	16'h	8d9b;
8634	:douta	=	16'h	8d5b;
8635	:douta	=	16'h	6cb9;
8636	:douta	=	16'h	4354;
8637	:douta	=	16'h	5c37;
8638	:douta	=	16'h	751b;
8639	:douta	=	16'h	6c99;
8640	:douta	=	16'h	6cb9;
8641	:douta	=	16'h	7d7c;
8642	:douta	=	16'h	751a;
8643	:douta	=	16'h	753b;
8644	:douta	=	16'h	859d;
8645	:douta	=	16'h	6cb9;
8646	:douta	=	16'h	6cd9;
8647	:douta	=	16'h	855a;
8648	:douta	=	16'h	9dfd;
8649	:douta	=	16'h	8d9c;
8650	:douta	=	16'h	6c99;
8651	:douta	=	16'h	751a;
8652	:douta	=	16'h	859c;
8653	:douta	=	16'h	859c;
8654	:douta	=	16'h	6cda;
8655	:douta	=	16'h	7d1b;
8656	:douta	=	16'h	74fa;
8657	:douta	=	16'h	74d9;
8658	:douta	=	16'h	8dbc;
8659	:douta	=	16'h	859c;
8660	:douta	=	16'h	751a;
8661	:douta	=	16'h	859c;
8662	:douta	=	16'h	859c;
8663	:douta	=	16'h	6cda;
8664	:douta	=	16'h	6cba;
8665	:douta	=	16'h	751a;
8666	:douta	=	16'h	7d1a;
8667	:douta	=	16'h	6cb9;
8668	:douta	=	16'h	859b;
8669	:douta	=	16'h	8d9b;
8670	:douta	=	16'h	857b;
8671	:douta	=	16'h	5bd6;
8672	:douta	=	16'h	5bd5;
8673	:douta	=	16'h	7d7c;
8674	:douta	=	16'h	857b;
8675	:douta	=	16'h	6cb9;
8676	:douta	=	16'h	6cfa;
8677	:douta	=	16'h	6d1a;
8678	:douta	=	16'h	74ba;
8679	:douta	=	16'h	857b;
8680	:douta	=	16'h	31a9;
8681	:douta	=	16'h	21a9;
8682	:douta	=	16'h	1127;
8683	:douta	=	16'h	1948;
8684	:douta	=	16'h	1968;
8685	:douta	=	16'h	2a2d;
8686	:douta	=	16'h	6438;
8687	:douta	=	16'h	220e;
8688	:douta	=	16'h	4b73;
8689	:douta	=	16'h	5393;
8690	:douta	=	16'h	9dda;
8691	:douta	=	16'h	6c36;
8692	:douta	=	16'h	8cd7;
8693	:douta	=	16'h	3b34;
8694	:douta	=	16'h	19ee;
8695	:douta	=	16'h	53d5;
8696	:douta	=	16'h	4b11;
8697	:douta	=	16'h	7c96;
8698	:douta	=	16'h	b61a;
8699	:douta	=	16'h	cefe;
8700	:douta	=	16'h	63f5;
8701	:douta	=	16'h	5c16;
8702	:douta	=	16'h	3333;
8703	:douta	=	16'h	4b95;
8704	:douta	=	16'h	32d1;
8705	:douta	=	16'h	3af2;
8706	:douta	=	16'h	32f2;
8707	:douta	=	16'h	4b73;
8708	:douta	=	16'h	8d9b;
8709	:douta	=	16'h	853a;
8710	:douta	=	16'h	74b8;
8711	:douta	=	16'h	6436;
8712	:douta	=	16'h	5352;
8713	:douta	=	16'h	5332;
8714	:douta	=	16'h	7456;
8715	:douta	=	16'h	6c36;
8716	:douta	=	16'h	6bf4;
8717	:douta	=	16'h	bdb8;
8718	:douta	=	16'h	9d16;
8719	:douta	=	16'h	9cf6;
8720	:douta	=	16'h	8c74;
8721	:douta	=	16'h	b596;
8722	:douta	=	16'h	8cb5;
8723	:douta	=	16'h	6bd2;
8724	:douta	=	16'h	6bd2;
8725	:douta	=	16'h	ad14;
8726	:douta	=	16'h	c5f8;
8727	:douta	=	16'h	d699;
8728	:douta	=	16'h	9453;
8729	:douta	=	16'h	ce38;
8730	:douta	=	16'h	6372;
8731	:douta	=	16'h	83f1;
8732	:douta	=	16'h	7c52;
8733	:douta	=	16'h	ad34;
8734	:douta	=	16'h	d677;
8735	:douta	=	16'h	eed9;
8736	:douta	=	16'h	a514;
8737	:douta	=	16'h	a4f4;
8738	:douta	=	16'h	7413;
8739	:douta	=	16'h	8c52;
8740	:douta	=	16'h	7c11;
8741	:douta	=	16'h	9cb2;
8742	:douta	=	16'h	e6b8;
8743	:douta	=	16'h	e6d8;
8744	:douta	=	16'h	9cf3;
8745	:douta	=	16'h	e6d8;
8746	:douta	=	16'h	b573;
8747	:douta	=	16'h	73b0;
8748	:douta	=	16'h	a553;
8749	:douta	=	16'h	528b;
8750	:douta	=	16'h	e6b6;
8751	:douta	=	16'h	e719;
8752	:douta	=	16'h	d616;
8753	:douta	=	16'h	7b8c;
8754	:douta	=	16'h	942f;
8755	:douta	=	16'h	8c4f;
8756	:douta	=	16'h	62eb;
8757	:douta	=	16'h	a510;
8758	:douta	=	16'h	8c2e;
8759	:douta	=	16'h	deb7;
8760	:douta	=	16'h	8bec;
8761	:douta	=	16'h	e697;
8762	:douta	=	16'h	732b;
8763	:douta	=	16'h	6b2a;
8764	:douta	=	16'h	62aa;
8765	:douta	=	16'h	5aaa;
8766	:douta	=	16'h	5249;
8767	:douta	=	16'h	2987;
8768	:douta	=	16'h	3a09;
8769	:douta	=	16'h	2967;
8770	:douta	=	16'h	1906;
8771	:douta	=	16'h	1926;
8772	:douta	=	16'h	1905;
8773	:douta	=	16'h	10a5;
8774	:douta	=	16'h	10e4;
8775	:douta	=	16'h	0042;
8776	:douta	=	16'h	736d;
8777	:douta	=	16'h	6b8f;
8778	:douta	=	16'h	e717;
8779	:douta	=	16'h	73f0;
8780	:douta	=	16'h	b512;
8781	:douta	=	16'h	b573;
8782	:douta	=	16'h	52aa;
8783	:douta	=	16'h	5b2c;
8784	:douta	=	16'h	18e4;
8785	:douta	=	16'h	8453;
8786	:douta	=	16'h	324d;
8787	:douta	=	16'h	5bd3;
8788	:douta	=	16'h	328d;
8789	:douta	=	16'h	4aad;
8790	:douta	=	16'h	5351;
8791	:douta	=	16'h	5b6f;
8792	:douta	=	16'h	4b30;
8793	:douta	=	16'h	11ab;
8794	:douta	=	16'h	a5b7;
8795	:douta	=	16'h	39e9;
8796	:douta	=	16'h	2945;
8797	:douta	=	16'h	18e2;
8798	:douta	=	16'h	20e3;
8799	:douta	=	16'h	18e3;
8800	:douta	=	16'h	1082;
8801	:douta	=	16'h	0820;
8802	:douta	=	16'h	3a2a;
8803	:douta	=	16'h	4aef;
8804	:douta	=	16'h	19ec;
8805	:douta	=	16'h	00e6;
8806	:douta	=	16'h	19ab;
8807	:douta	=	16'h	4bb5;
8808	:douta	=	16'h	5394;
8809	:douta	=	16'h	2ad1;
8810	:douta	=	16'h	7c97;
8811	:douta	=	16'h	4b72;
8812	:douta	=	16'h	3aaf;
8813	:douta	=	16'h	116a;
8814	:douta	=	16'h	3aaf;
8815	:douta	=	16'h	6477;
8816	:douta	=	16'h	53d5;
8817	:douta	=	16'h	53f5;
8818	:douta	=	16'h	53b4;
8819	:douta	=	16'h	9d38;
8820	:douta	=	16'h	4333;
8821	:douta	=	16'h	4b52;
8822	:douta	=	16'h	3270;
8823	:douta	=	16'h	63f4;
8824	:douta	=	16'h	53d4;
8825	:douta	=	16'h	7476;
8826	:douta	=	16'h	6c76;
8827	:douta	=	16'h	6c36;
8828	:douta	=	16'h	63f4;
8829	:douta	=	16'h	6c55;
8830	:douta	=	16'h	9579;
8831	:douta	=	16'h	63f5;
8832	:douta	=	16'h	4a8c;
8833	:douta	=	16'h	39a6;
8834	:douta	=	16'h	4209;
8835	:douta	=	16'h	2127;
8836	:douta	=	16'h	934b;
8837	:douta	=	16'h	634d;
8838	:douta	=	16'h	73f3;
8839	:douta	=	16'h	7496;
8840	:douta	=	16'h	955a;
8841	:douta	=	16'h	7c97;
8842	:douta	=	16'h	9d9a;
8843	:douta	=	16'h	84d7;
8844	:douta	=	16'h	7476;
8845	:douta	=	16'h	7c96;
8846	:douta	=	16'h	84d7;
8847	:douta	=	16'h	6c15;
8848	:douta	=	16'h	6c15;
8849	:douta	=	16'h	7cb7;
8850	:douta	=	16'h	7c97;
8851	:douta	=	16'h	84d8;
8852	:douta	=	16'h	8d59;
8853	:douta	=	16'h	8d39;
8854	:douta	=	16'h	7cf8;
8855	:douta	=	16'h	7cb8;
8856	:douta	=	16'h	84f9;
8857	:douta	=	16'h	8d7a;
8858	:douta	=	16'h	8d3a;
8859	:douta	=	16'h	7cb8;
8860	:douta	=	16'h	957a;
8861	:douta	=	16'h	959b;
8862	:douta	=	16'h	8d5a;
8863	:douta	=	16'h	8d39;
8864	:douta	=	16'h	7d19;
8865	:douta	=	16'h	8d3b;
8866	:douta	=	16'h	8d9b;
8867	:douta	=	16'h	853a;
8868	:douta	=	16'h	84f9;
8869	:douta	=	16'h	8d3a;
8870	:douta	=	16'h	7cf9;
8871	:douta	=	16'h	8d5b;
8872	:douta	=	16'h	959c;
8873	:douta	=	16'h	959b;
8874	:douta	=	16'h	7cf9;
8875	:douta	=	16'h	7cf9;
8876	:douta	=	16'h	8d5b;
8877	:douta	=	16'h	8d9b;
8878	:douta	=	16'h	8d5b;
8879	:douta	=	16'h	8519;
8880	:douta	=	16'h	853a;
8881	:douta	=	16'h	959b;
8882	:douta	=	16'h	8d5b;
8883	:douta	=	16'h	853a;
8884	:douta	=	16'h	8d5a;
8885	:douta	=	16'h	7477;
8886	:douta	=	16'h	8539;
8887	:douta	=	16'h	8d7b;
8888	:douta	=	16'h	8d7b;
8889	:douta	=	16'h	853a;
8890	:douta	=	16'h	8d7b;
8891	:douta	=	16'h	959c;
8892	:douta	=	16'h	74b9;
8893	:douta	=	16'h	6458;
8894	:douta	=	16'h	53d6;
8895	:douta	=	16'h	5c58;
8896	:douta	=	16'h	6478;
8897	:douta	=	16'h	6cd9;
8898	:douta	=	16'h	7d5b;
8899	:douta	=	16'h	6478;
8900	:douta	=	16'h	753b;
8901	:douta	=	16'h	7d3b;
8902	:douta	=	16'h	7d3b;
8903	:douta	=	16'h	74da;
8904	:douta	=	16'h	857b;
8905	:douta	=	16'h	95fd;
8906	:douta	=	16'h	8dbc;
8907	:douta	=	16'h	6c99;
8908	:douta	=	16'h	6cfa;
8909	:douta	=	16'h	8dbd;
8910	:douta	=	16'h	8dbc;
8911	:douta	=	16'h	751a;
8912	:douta	=	16'h	7d1a;
8913	:douta	=	16'h	6cb9;
8914	:douta	=	16'h	74fa;
8915	:douta	=	16'h	7d3b;
8916	:douta	=	16'h	859c;
8917	:douta	=	16'h	751b;
8918	:douta	=	16'h	7d7b;
8919	:douta	=	16'h	7d5b;
8920	:douta	=	16'h	751a;
8921	:douta	=	16'h	6cda;
8922	:douta	=	16'h	7d3b;
8923	:douta	=	16'h	8dbc;
8924	:douta	=	16'h	7d1a;
8925	:douta	=	16'h	7d1a;
8926	:douta	=	16'h	8dbc;
8927	:douta	=	16'h	857b;
8928	:douta	=	16'h	6c78;
8929	:douta	=	16'h	5bf6;
8930	:douta	=	16'h	74d9;
8931	:douta	=	16'h	859c;
8932	:douta	=	16'h	74da;
8933	:douta	=	16'h	6498;
8934	:douta	=	16'h	753a;
8935	:douta	=	16'h	6cd9;
8936	:douta	=	16'h	7c98;
8937	:douta	=	16'h	2988;
8938	:douta	=	16'h	29ca;
8939	:douta	=	16'h	1927;
8940	:douta	=	16'h	1948;
8941	:douta	=	16'h	08a5;
8942	:douta	=	16'h	5c37;
8943	:douta	=	16'h	5bf5;
8944	:douta	=	16'h	5394;
8945	:douta	=	16'h	4b33;
8946	:douta	=	16'h	1a4f;
8947	:douta	=	16'h	a579;
8948	:douta	=	16'h	c69d;
8949	:douta	=	16'h	851a;
8950	:douta	=	16'h	6457;
8951	:douta	=	16'h	4bb5;
8952	:douta	=	16'h	5393;
8953	:douta	=	16'h	3af2;
8954	:douta	=	16'h	84f7;
8955	:douta	=	16'h	9559;
8956	:douta	=	16'h	adb9;
8957	:douta	=	16'h	7cb8;
8958	:douta	=	16'h	6416;
8959	:douta	=	16'h	7cda;
8960	:douta	=	16'h	32f2;
8961	:douta	=	16'h	4375;
8962	:douta	=	16'h	74d9;
8963	:douta	=	16'h	4312;
8964	:douta	=	16'h	74b9;
8965	:douta	=	16'h	6c78;
8966	:douta	=	16'h	3af1;
8967	:douta	=	16'h	2a70;
8968	:douta	=	16'h	5b93;
8969	:douta	=	16'h	5b73;
8970	:douta	=	16'h	7414;
8971	:douta	=	16'h	6bd4;
8972	:douta	=	16'h	8475;
8973	:douta	=	16'h	7c33;
8974	:douta	=	16'h	8cd5;
8975	:douta	=	16'h	6bd2;
8976	:douta	=	16'h	6b71;
8977	:douta	=	16'h	6350;
8978	:douta	=	16'h	c5f8;
8979	:douta	=	16'h	8c94;
8980	:douta	=	16'h	ad56;
8981	:douta	=	16'h	9cd4;
8982	:douta	=	16'h	c5f7;
8983	:douta	=	16'h	8453;
8984	:douta	=	16'h	8453;
8985	:douta	=	16'h	ad55;
8986	:douta	=	16'h	b555;
8987	:douta	=	16'h	d657;
8988	:douta	=	16'h	94b5;
8989	:douta	=	16'h	deb9;
8990	:douta	=	16'h	8cb5;
8991	:douta	=	16'h	a4d2;
8992	:douta	=	16'h	ad75;
8993	:douta	=	16'h	9cd3;
8994	:douta	=	16'h	bdb4;
8995	:douta	=	16'h	f738;
8996	:douta	=	16'h	a4f2;
8997	:douta	=	16'h	c5d5;
8998	:douta	=	16'h	f719;
8999	:douta	=	16'h	c5b5;
9000	:douta	=	16'h	ce37;
9001	:douta	=	16'h	cdf5;
9002	:douta	=	16'h	ce14;
9003	:douta	=	16'h	de76;
9004	:douta	=	16'h	ce76;
9005	:douta	=	16'h	a48f;
9006	:douta	=	16'h	e6f9;
9007	:douta	=	16'h	ce16;
9008	:douta	=	16'h	9c91;
9009	:douta	=	16'h	6b4d;
9010	:douta	=	16'h	b531;
9011	:douta	=	16'h	b551;
9012	:douta	=	16'h	ad10;
9013	:douta	=	16'h	c5d3;
9014	:douta	=	16'h	d5f4;
9015	:douta	=	16'h	de96;
9016	:douta	=	16'h	5269;
9017	:douta	=	16'h	7b4b;
9018	:douta	=	16'h	732b;
9019	:douta	=	16'h	62ca;
9020	:douta	=	16'h	62a9;
9021	:douta	=	16'h	31a7;
9022	:douta	=	16'h	41e7;
9023	:douta	=	16'h	2167;
9024	:douta	=	16'h	2987;
9025	:douta	=	16'h	31e9;
9026	:douta	=	16'h	2968;
9027	:douta	=	16'h	2988;
9028	:douta	=	16'h	29a9;
9029	:douta	=	16'h	10e4;
9030	:douta	=	16'h	10c4;
9031	:douta	=	16'h	0084;
9032	:douta	=	16'h	39c7;
9033	:douta	=	16'h	4aac;
9034	:douta	=	16'h	9cf1;
9035	:douta	=	16'h	530c;
9036	:douta	=	16'h	6b4c;
9037	:douta	=	16'h	840f;
9038	:douta	=	16'h	b552;
9039	:douta	=	16'h	7bce;
9040	:douta	=	16'h	634d;
9041	:douta	=	16'h	6c34;
9042	:douta	=	16'h	8d58;
9043	:douta	=	16'h	4b31;
9044	:douta	=	16'h	1148;
9045	:douta	=	16'h	29c9;
9046	:douta	=	16'h	3209;
9047	:douta	=	16'h	9472;
9048	:douta	=	16'h	84f7;
9049	:douta	=	16'h	4331;
9050	:douta	=	16'h	53b3;
9051	:douta	=	16'h	4b0f;
9052	:douta	=	16'h	5bb2;
9053	:douta	=	16'h	3a0c;
9054	:douta	=	16'h	31c7;
9055	:douta	=	16'h	1061;
9056	:douta	=	16'h	20e3;
9057	:douta	=	16'h	18e4;
9058	:douta	=	16'h	18e3;
9059	:douta	=	16'h	1061;
9060	:douta	=	16'h	1967;
9061	:douta	=	16'h	5bb4;
9062	:douta	=	16'h	3b11;
9063	:douta	=	16'h	00e7;
9064	:douta	=	16'h	220c;
9065	:douta	=	16'h	32d1;
9066	:douta	=	16'h	3b11;
9067	:douta	=	16'h	3b31;
9068	:douta	=	16'h	53b4;
9069	:douta	=	16'h	4b73;
9070	:douta	=	16'h	6c33;
9071	:douta	=	16'h	29ec;
9072	:douta	=	16'h	5351;
9073	:douta	=	16'h	216a;
9074	:douta	=	16'h	322c;
9075	:douta	=	16'h	4b31;
9076	:douta	=	16'h	5c15;
9077	:douta	=	16'h	6477;
9078	:douta	=	16'h	53d5;
9079	:douta	=	16'h	74b8;
9080	:douta	=	16'h	6cb8;
9081	:douta	=	16'h	74f9;
9082	:douta	=	16'h	53d5;
9083	:douta	=	16'h	6bd2;
9084	:douta	=	16'h	7c96;
9085	:douta	=	16'h	21cc;
9086	:douta	=	16'h	4b10;
9087	:douta	=	16'h	52f0;
9088	:douta	=	16'h	4208;
9089	:douta	=	16'h	4229;
9090	:douta	=	16'h	5a29;
9091	:douta	=	16'h	836c;
9092	:douta	=	16'h	528d;
9093	:douta	=	16'h	84d8;
9094	:douta	=	16'h	7476;
9095	:douta	=	16'h	9d9a;
9096	:douta	=	16'h	7c97;
9097	:douta	=	16'h	7435;
9098	:douta	=	16'h	7cb7;
9099	:douta	=	16'h	9519;
9100	:douta	=	16'h	7cb7;
9101	:douta	=	16'h	84f8;
9102	:douta	=	16'h	8d18;
9103	:douta	=	16'h	7456;
9104	:douta	=	16'h	7456;
9105	:douta	=	16'h	8d18;
9106	:douta	=	16'h	7cb8;
9107	:douta	=	16'h	84d8;
9108	:douta	=	16'h	7c98;
9109	:douta	=	16'h	7cb8;
9110	:douta	=	16'h	7cd8;
9111	:douta	=	16'h	84f9;
9112	:douta	=	16'h	7497;
9113	:douta	=	16'h	6c56;
9114	:douta	=	16'h	6c56;
9115	:douta	=	16'h	8d3a;
9116	:douta	=	16'h	7cd8;
9117	:douta	=	16'h	7cd8;
9118	:douta	=	16'h	7cd8;
9119	:douta	=	16'h	8519;
9120	:douta	=	16'h	855a;
9121	:douta	=	16'h	8519;
9122	:douta	=	16'h	7c98;
9123	:douta	=	16'h	7cb9;
9124	:douta	=	16'h	8d5a;
9125	:douta	=	16'h	853a;
9126	:douta	=	16'h	851a;
9127	:douta	=	16'h	8d7b;
9128	:douta	=	16'h	8d7b;
9129	:douta	=	16'h	853a;
9130	:douta	=	16'h	853a;
9131	:douta	=	16'h	853a;
9132	:douta	=	16'h	8d5a;
9133	:douta	=	16'h	8d9b;
9134	:douta	=	16'h	8d7b;
9135	:douta	=	16'h	959c;
9136	:douta	=	16'h	9ddc;
9137	:douta	=	16'h	853a;
9138	:douta	=	16'h	8d5a;
9139	:douta	=	16'h	8d7a;
9140	:douta	=	16'h	95bb;
9141	:douta	=	16'h	959b;
9142	:douta	=	16'h	8d5a;
9143	:douta	=	16'h	8519;
9144	:douta	=	16'h	8d3a;
9145	:douta	=	16'h	8d5a;
9146	:douta	=	16'h	959c;
9147	:douta	=	16'h	851a;
9148	:douta	=	16'h	959c;
9149	:douta	=	16'h	959c;
9150	:douta	=	16'h	95bc;
9151	:douta	=	16'h	853a;
9152	:douta	=	16'h	6458;
9153	:douta	=	16'h	6458;
9154	:douta	=	16'h	6c98;
9155	:douta	=	16'h	74fa;
9156	:douta	=	16'h	6478;
9157	:douta	=	16'h	64b9;
9158	:douta	=	16'h	7d5c;
9159	:douta	=	16'h	7d7b;
9160	:douta	=	16'h	857c;
9161	:douta	=	16'h	8dfd;
9162	:douta	=	16'h	7d5b;
9163	:douta	=	16'h	8dbd;
9164	:douta	=	16'h	8d9c;
9165	:douta	=	16'h	7d5b;
9166	:douta	=	16'h	6cba;
9167	:douta	=	16'h	95bc;
9168	:douta	=	16'h	857c;
9169	:douta	=	16'h	7d3b;
9170	:douta	=	16'h	857c;
9171	:douta	=	16'h	7d3a;
9172	:douta	=	16'h	7d3b;
9173	:douta	=	16'h	857c;
9174	:douta	=	16'h	855b;
9175	:douta	=	16'h	74fa;
9176	:douta	=	16'h	753b;
9177	:douta	=	16'h	8d9b;
9178	:douta	=	16'h	751a;
9179	:douta	=	16'h	6499;
9180	:douta	=	16'h	751a;
9181	:douta	=	16'h	7d5a;
9182	:douta	=	16'h	8dbc;
9183	:douta	=	16'h	74d9;
9184	:douta	=	16'h	74fa;
9185	:douta	=	16'h	7d3a;
9186	:douta	=	16'h	74d9;
9187	:douta	=	16'h	5c16;
9188	:douta	=	16'h	753a;
9189	:douta	=	16'h	7d7b;
9190	:douta	=	16'h	74b9;
9191	:douta	=	16'h	6cb9;
9192	:douta	=	16'h	6cfa;
9193	:douta	=	16'h	7cfa;
9194	:douta	=	16'h	5b53;
9195	:douta	=	16'h	29a8;
9196	:douta	=	16'h	2188;
9197	:douta	=	16'h	1968;
9198	:douta	=	16'h	1148;
9199	:douta	=	16'h	53d4;
9200	:douta	=	16'h	9538;
9201	:douta	=	16'h	b61b;
9202	:douta	=	16'h	84f8;
9203	:douta	=	16'h	5c16;
9204	:douta	=	16'h	32b0;
9205	:douta	=	16'h	220d;
9206	:douta	=	16'h	3ad1;
9207	:douta	=	16'h	5392;
9208	:douta	=	16'h	8d17;
9209	:douta	=	16'h	be3b;
9210	:douta	=	16'h	53b4;
9211	:douta	=	16'h	7456;
9212	:douta	=	16'h	3b12;
9213	:douta	=	16'h	6c77;
9214	:douta	=	16'h	74d8;
9215	:douta	=	16'h	84d7;
9216	:douta	=	16'h	2ad0;
9217	:douta	=	16'h	2ab1;
9218	:douta	=	16'h	4333;
9219	:douta	=	16'h	53f5;
9220	:douta	=	16'h	7d3b;
9221	:douta	=	16'h	7d3a;
9222	:douta	=	16'h	6477;
9223	:douta	=	16'h	74da;
9224	:douta	=	16'h	5352;
9225	:douta	=	16'h	4b11;
9226	:douta	=	16'h	5353;
9227	:douta	=	16'h	4b31;
9228	:douta	=	16'h	5331;
9229	:douta	=	16'h	a557;
9230	:douta	=	16'h	ad77;
9231	:douta	=	16'h	9d17;
9232	:douta	=	16'h	8c74;
9233	:douta	=	16'h	8c33;
9234	:douta	=	16'h	7433;
9235	:douta	=	16'h	6bd2;
9236	:douta	=	16'h	8cb5;
9237	:douta	=	16'h	9451;
9238	:douta	=	16'h	bd96;
9239	:douta	=	16'h	e6fa;
9240	:douta	=	16'h	8c74;
9241	:douta	=	16'h	b596;
9242	:douta	=	16'h	b575;
9243	:douta	=	16'h	c5d6;
9244	:douta	=	16'h	73f2;
9245	:douta	=	16'h	e698;
9246	:douta	=	16'h	ce16;
9247	:douta	=	16'h	de97;
9248	:douta	=	16'h	de98;
9249	:douta	=	16'h	6b70;
9250	:douta	=	16'h	8c31;
9251	:douta	=	16'h	c5b5;
9252	:douta	=	16'h	8c51;
9253	:douta	=	16'h	ad33;
9254	:douta	=	16'h	deb8;
9255	:douta	=	16'h	e6b8;
9256	:douta	=	16'h	d637;
9257	:douta	=	16'h	ef18;
9258	:douta	=	16'h	c5f4;
9259	:douta	=	16'h	e6f8;
9260	:douta	=	16'h	a4d0;
9261	:douta	=	16'h	840f;
9262	:douta	=	16'h	ce14;
9263	:douta	=	16'h	ce35;
9264	:douta	=	16'h	eeb7;
9265	:douta	=	16'h	4a49;
9266	:douta	=	16'h	bd12;
9267	:douta	=	16'h	94af;
9268	:douta	=	16'h	946f;
9269	:douta	=	16'h	94af;
9270	:douta	=	16'h	cd93;
9271	:douta	=	16'h	f759;
9272	:douta	=	16'h	732b;
9273	:douta	=	16'h	7b4c;
9274	:douta	=	16'h	732a;
9275	:douta	=	16'h	62ca;
9276	:douta	=	16'h	5a68;
9277	:douta	=	16'h	5249;
9278	:douta	=	16'h	4208;
9279	:douta	=	16'h	1926;
9280	:douta	=	16'h	18e5;
9281	:douta	=	16'h	1925;
9282	:douta	=	16'h	10e4;
9283	:douta	=	16'h	1905;
9284	:douta	=	16'h	2968;
9285	:douta	=	16'h	10e5;
9286	:douta	=	16'h	10e5;
9287	:douta	=	16'h	1105;
9288	:douta	=	16'h	0883;
9289	:douta	=	16'h	7bcf;
9290	:douta	=	16'h	bdf5;
9291	:douta	=	16'h	322a;
9292	:douta	=	16'h	83ad;
9293	:douta	=	16'h	ad73;
9294	:douta	=	16'h	5aaa;
9295	:douta	=	16'h	6baf;
9296	:douta	=	16'h	7c53;
9297	:douta	=	16'h	532f;
9298	:douta	=	16'h	74b5;
9299	:douta	=	16'h	5b4e;
9300	:douta	=	16'h	21a9;
9301	:douta	=	16'h	428c;
9302	:douta	=	16'h	10a5;
9303	:douta	=	16'h	8c30;
9304	:douta	=	16'h	7cb6;
9305	:douta	=	16'h	4b51;
9306	:douta	=	16'h	4310;
9307	:douta	=	16'h	52ee;
9308	:douta	=	16'h	5330;
9309	:douta	=	16'h	4aef;
9310	:douta	=	16'h	94f5;
9311	:douta	=	16'h	1926;
9312	:douta	=	16'h	18a2;
9313	:douta	=	16'h	18e3;
9314	:douta	=	16'h	1082;
9315	:douta	=	16'h	10a2;
9316	:douta	=	16'h	0000;
9317	:douta	=	16'h	29c9;
9318	:douta	=	16'h	4b11;
9319	:douta	=	16'h	2a0d;
9320	:douta	=	16'h	1149;
9321	:douta	=	16'h	19cc;
9322	:douta	=	16'h	4bb5;
9323	:douta	=	16'h	53d5;
9324	:douta	=	16'h	2a4e;
9325	:douta	=	16'h	2a8f;
9326	:douta	=	16'h	63d4;
9327	:douta	=	16'h	5392;
9328	:douta	=	16'h	5bd4;
9329	:douta	=	16'h	53b4;
9330	:douta	=	16'h	5b91;
9331	:douta	=	16'h	4b72;
9332	:douta	=	16'h	4332;
9333	:douta	=	16'h	1a2e;
9334	:douta	=	16'h	53d5;
9335	:douta	=	16'h	6436;
9336	:douta	=	16'h	5c57;
9337	:douta	=	16'h	6477;
9338	:douta	=	16'h	5c16;
9339	:douta	=	16'h	9579;
9340	:douta	=	16'h	8dbc;
9341	:douta	=	16'h	4aae;
9342	:douta	=	16'h	63b2;
9343	:douta	=	16'h	4a09;
9344	:douta	=	16'h	4229;
9345	:douta	=	16'h	2968;
9346	:douta	=	16'h	c4cf;
9347	:douta	=	16'h	5a6c;
9348	:douta	=	16'h	8454;
9349	:douta	=	16'h	84d7;
9350	:douta	=	16'h	6bd4;
9351	:douta	=	16'h	adfb;
9352	:douta	=	16'h	9559;
9353	:douta	=	16'h	8d18;
9354	:douta	=	16'h	63f4;
9355	:douta	=	16'h	7c96;
9356	:douta	=	16'h	957a;
9357	:douta	=	16'h	63f5;
9358	:douta	=	16'h	6c15;
9359	:douta	=	16'h	9559;
9360	:douta	=	16'h	8d18;
9361	:douta	=	16'h	7456;
9362	:douta	=	16'h	8d39;
9363	:douta	=	16'h	8d19;
9364	:douta	=	16'h	84d8;
9365	:douta	=	16'h	7497;
9366	:douta	=	16'h	6c57;
9367	:douta	=	16'h	84f9;
9368	:douta	=	16'h	957a;
9369	:douta	=	16'h	8d39;
9370	:douta	=	16'h	84f9;
9371	:douta	=	16'h	5bd5;
9372	:douta	=	16'h	957a;
9373	:douta	=	16'h	957a;
9374	:douta	=	16'h	84f8;
9375	:douta	=	16'h	8d5a;
9376	:douta	=	16'h	853a;
9377	:douta	=	16'h	8d7b;
9378	:douta	=	16'h	8d5a;
9379	:douta	=	16'h	7498;
9380	:douta	=	16'h	7498;
9381	:douta	=	16'h	959b;
9382	:douta	=	16'h	853a;
9383	:douta	=	16'h	7cf9;
9384	:douta	=	16'h	959c;
9385	:douta	=	16'h	857b;
9386	:douta	=	16'h	8d7b;
9387	:douta	=	16'h	853a;
9388	:douta	=	16'h	8d7b;
9389	:douta	=	16'h	8d5a;
9390	:douta	=	16'h	855a;
9391	:douta	=	16'h	8d5b;
9392	:douta	=	16'h	8d7b;
9393	:douta	=	16'h	8d7b;
9394	:douta	=	16'h	959b;
9395	:douta	=	16'h	853a;
9396	:douta	=	16'h	957b;
9397	:douta	=	16'h	8d7b;
9398	:douta	=	16'h	a5dc;
9399	:douta	=	16'h	851a;
9400	:douta	=	16'h	851a;
9401	:douta	=	16'h	851a;
9402	:douta	=	16'h	853a;
9403	:douta	=	16'h	8d7b;
9404	:douta	=	16'h	8d5a;
9405	:douta	=	16'h	8d7b;
9406	:douta	=	16'h	95bc;
9407	:douta	=	16'h	95bc;
9408	:douta	=	16'h	8d9b;
9409	:douta	=	16'h	6c98;
9410	:douta	=	16'h	5bf6;
9411	:douta	=	16'h	751a;
9412	:douta	=	16'h	7d5b;
9413	:douta	=	16'h	6c99;
9414	:douta	=	16'h	6cfa;
9415	:douta	=	16'h	7d3b;
9416	:douta	=	16'h	6cba;
9417	:douta	=	16'h	753b;
9418	:douta	=	16'h	7d5c;
9419	:douta	=	16'h	859c;
9420	:douta	=	16'h	7d7b;
9421	:douta	=	16'h	95dc;
9422	:douta	=	16'h	8d9c;
9423	:douta	=	16'h	74fb;
9424	:douta	=	16'h	857b;
9425	:douta	=	16'h	857b;
9426	:douta	=	16'h	8d9c;
9427	:douta	=	16'h	7d3b;
9428	:douta	=	16'h	7d3b;
9429	:douta	=	16'h	7d1a;
9430	:douta	=	16'h	857b;
9431	:douta	=	16'h	7d3b;
9432	:douta	=	16'h	6cb9;
9433	:douta	=	16'h	7d3b;
9434	:douta	=	16'h	85bc;
9435	:douta	=	16'h	857b;
9436	:douta	=	16'h	6cda;
9437	:douta	=	16'h	64b9;
9438	:douta	=	16'h	8dbc;
9439	:douta	=	16'h	7d3a;
9440	:douta	=	16'h	7499;
9441	:douta	=	16'h	7d1a;
9442	:douta	=	16'h	855b;
9443	:douta	=	16'h	6437;
9444	:douta	=	16'h	6478;
9445	:douta	=	16'h	6cb9;
9446	:douta	=	16'h	8dbc;
9447	:douta	=	16'h	7d3b;
9448	:douta	=	16'h	7d1a;
9449	:douta	=	16'h	6499;
9450	:douta	=	16'h	74fa;
9451	:douta	=	16'h	31ea;
9452	:douta	=	16'h	31a8;
9453	:douta	=	16'h	1908;
9454	:douta	=	16'h	1967;
9455	:douta	=	16'h	1968;
9456	:douta	=	16'h	5c16;
9457	:douta	=	16'h	5c15;
9458	:douta	=	16'h	a5ba;
9459	:douta	=	16'h	7497;
9460	:douta	=	16'h	7cb8;
9461	:douta	=	16'h	3b32;
9462	:douta	=	16'h	5351;
9463	:douta	=	16'h	1a0e;
9464	:douta	=	16'h	7cb7;
9465	:douta	=	16'h	957a;
9466	:douta	=	16'h	84b7;
9467	:douta	=	16'h	b63b;
9468	:douta	=	16'h	6c55;
9469	:douta	=	16'h	6456;
9470	:douta	=	16'h	1a50;
9471	:douta	=	16'h	8d39;
9472	:douta	=	16'h	3b53;
9473	:douta	=	16'h	4bf6;
9474	:douta	=	16'h	4bf6;
9475	:douta	=	16'h	5416;
9476	:douta	=	16'h	42f1;
9477	:douta	=	16'h	5c16;
9478	:douta	=	16'h	5373;
9479	:douta	=	16'h	32b1;
9480	:douta	=	16'h	6c15;
9481	:douta	=	16'h	6c14;
9482	:douta	=	16'h	7c55;
9483	:douta	=	16'h	8d18;
9484	:douta	=	16'h	8d18;
9485	:douta	=	16'h	5b30;
9486	:douta	=	16'h	6bd2;
9487	:douta	=	16'h	7c53;
9488	:douta	=	16'h	6350;
9489	:douta	=	16'h	8c53;
9490	:douta	=	16'h	9d16;
9491	:douta	=	16'h	b5f9;
9492	:douta	=	16'h	94d5;
9493	:douta	=	16'h	ce17;
9494	:douta	=	16'h	a556;
9495	:douta	=	16'h	9494;
9496	:douta	=	16'h	5b50;
9497	:douta	=	16'h	94b3;
9498	:douta	=	16'h	9cd3;
9499	:douta	=	16'h	c5f6;
9500	:douta	=	16'h	c637;
9501	:douta	=	16'h	a4f4;
9502	:douta	=	16'h	c5b5;
9503	:douta	=	16'h	bdb6;
9504	:douta	=	16'h	ad74;
9505	:douta	=	16'h	b533;
9506	:douta	=	16'h	d637;
9507	:douta	=	16'h	de77;
9508	:douta	=	16'h	9471;
9509	:douta	=	16'h	c5f5;
9510	:douta	=	16'h	d5f7;
9511	:douta	=	16'h	bdb5;
9512	:douta	=	16'h	bd95;
9513	:douta	=	16'h	ad11;
9514	:douta	=	16'h	d655;
9515	:douta	=	16'h	ad11;
9516	:douta	=	16'h	bd53;
9517	:douta	=	16'h	b531;
9518	:douta	=	16'h	de97;
9519	:douta	=	16'h	eef9;
9520	:douta	=	16'h	7bac;
9521	:douta	=	16'h	630c;
9522	:douta	=	16'h	732b;
9523	:douta	=	16'h	c5f4;
9524	:douta	=	16'h	b531;
9525	:douta	=	16'h	b532;
9526	:douta	=	16'h	c5f3;
9527	:douta	=	16'h	83ed;
9528	:douta	=	16'h	838c;
9529	:douta	=	16'h	7b4b;
9530	:douta	=	16'h	6b0a;
9531	:douta	=	16'h	62ca;
9532	:douta	=	16'h	732b;
9533	:douta	=	16'h	4a27;
9534	:douta	=	16'h	1945;
9535	:douta	=	16'h	10a4;
9536	:douta	=	16'h	0883;
9537	:douta	=	16'h	18e5;
9538	:douta	=	16'h	1906;
9539	:douta	=	16'h	1105;
9540	:douta	=	16'h	2146;
9541	:douta	=	16'h	2167;
9542	:douta	=	16'h	1905;
9543	:douta	=	16'h	10e5;
9544	:douta	=	16'h	10c4;
9545	:douta	=	16'h	62aa;
9546	:douta	=	16'h	6bee;
9547	:douta	=	16'h	4a4a;
9548	:douta	=	16'h	8c4f;
9549	:douta	=	16'h	9cf2;
9550	:douta	=	16'h	630c;
9551	:douta	=	16'h	63b2;
9552	:douta	=	16'h	6bf2;
9553	:douta	=	16'h	532f;
9554	:douta	=	16'h	3a4c;
9555	:douta	=	16'h	8c72;
9556	:douta	=	16'h	632d;
9557	:douta	=	16'h	7c30;
9558	:douta	=	16'h	29a8;
9559	:douta	=	16'h	840f;
9560	:douta	=	16'h	2989;
9561	:douta	=	16'h	52ac;
9562	:douta	=	16'h	3a6d;
9563	:douta	=	16'h	63b1;
9564	:douta	=	16'h	5b70;
9565	:douta	=	16'h	42ce;
9566	:douta	=	16'h	532f;
9567	:douta	=	16'h	63d1;
9568	:douta	=	16'h	42cf;
9569	:douta	=	16'h	3a6b;
9570	:douta	=	16'h	0820;
9571	:douta	=	16'h	1082;
9572	:douta	=	16'h	10a3;
9573	:douta	=	16'h	0040;
9574	:douta	=	16'h	0000;
9575	:douta	=	16'h	1925;
9576	:douta	=	16'h	4b0e;
9577	:douta	=	16'h	19ab;
9578	:douta	=	16'h	32af;
9579	:douta	=	16'h	328f;
9580	:douta	=	16'h	53f6;
9581	:douta	=	16'h	53f5;
9582	:douta	=	16'h	5393;
9583	:douta	=	16'h	324e;
9584	:douta	=	16'h	42f1;
9585	:douta	=	16'h	21ec;
9586	:douta	=	16'h	3acf;
9587	:douta	=	16'h	32af;
9588	:douta	=	16'h	4bd5;
9589	:douta	=	16'h	4374;
9590	:douta	=	16'h	63f4;
9591	:douta	=	16'h	853a;
9592	:douta	=	16'h	6c98;
9593	:douta	=	16'h	224f;
9594	:douta	=	16'h	42f1;
9595	:douta	=	16'h	6415;
9596	:douta	=	16'h	5393;
9597	:douta	=	16'h	5b93;
9598	:douta	=	16'h	5249;
9599	:douta	=	16'h	3a4a;
9600	:douta	=	16'h	a3ed;
9601	:douta	=	16'h	a44f;
9602	:douta	=	16'h	632f;
9603	:douta	=	16'h	7cb7;
9604	:douta	=	16'h	7c76;
9605	:douta	=	16'h	959a;
9606	:douta	=	16'h	959a;
9607	:douta	=	16'h	5b93;
9608	:douta	=	16'h	7cb8;
9609	:douta	=	16'h	8d5a;
9610	:douta	=	16'h	957b;
9611	:douta	=	16'h	957b;
9612	:douta	=	16'h	8d39;
9613	:douta	=	16'h	7c96;
9614	:douta	=	16'h	7c97;
9615	:douta	=	16'h	84b8;
9616	:douta	=	16'h	7477;
9617	:douta	=	16'h	9559;
9618	:douta	=	16'h	7476;
9619	:douta	=	16'h	6c56;
9620	:douta	=	16'h	7456;
9621	:douta	=	16'h	7c97;
9622	:douta	=	16'h	8d39;
9623	:douta	=	16'h	8519;
9624	:douta	=	16'h	7497;
9625	:douta	=	16'h	7cb8;
9626	:douta	=	16'h	84d8;
9627	:douta	=	16'h	8d7a;
9628	:douta	=	16'h	7c98;
9629	:douta	=	16'h	7c98;
9630	:douta	=	16'h	8519;
9631	:douta	=	16'h	6c56;
9632	:douta	=	16'h	7457;
9633	:douta	=	16'h	6c36;
9634	:douta	=	16'h	853a;
9635	:douta	=	16'h	7cd9;
9636	:douta	=	16'h	7cd9;
9637	:douta	=	16'h	8d7b;
9638	:douta	=	16'h	8d5a;
9639	:douta	=	16'h	959b;
9640	:douta	=	16'h	8d7b;
9641	:douta	=	16'h	8d5a;
9642	:douta	=	16'h	6416;
9643	:douta	=	16'h	7498;
9644	:douta	=	16'h	959b;
9645	:douta	=	16'h	959b;
9646	:douta	=	16'h	855a;
9647	:douta	=	16'h	8d5b;
9648	:douta	=	16'h	8d5a;
9649	:douta	=	16'h	959b;
9650	:douta	=	16'h	851a;
9651	:douta	=	16'h	84f9;
9652	:douta	=	16'h	8d5a;
9653	:douta	=	16'h	95bc;
9654	:douta	=	16'h	8d3a;
9655	:douta	=	16'h	959b;
9656	:douta	=	16'h	957b;
9657	:douta	=	16'h	959b;
9658	:douta	=	16'h	8d7b;
9659	:douta	=	16'h	8d5a;
9660	:douta	=	16'h	8d5b;
9661	:douta	=	16'h	851a;
9662	:douta	=	16'h	855a;
9663	:douta	=	16'h	95bc;
9664	:douta	=	16'h	8d5a;
9665	:douta	=	16'h	95bc;
9666	:douta	=	16'h	95dc;
9667	:douta	=	16'h	853b;
9668	:douta	=	16'h	6438;
9669	:douta	=	16'h	74da;
9670	:douta	=	16'h	8ddc;
9671	:douta	=	16'h	7d5b;
9672	:douta	=	16'h	74fb;
9673	:douta	=	16'h	6cda;
9674	:douta	=	16'h	64b9;
9675	:douta	=	16'h	85bd;
9676	:douta	=	16'h	7d5b;
9677	:douta	=	16'h	753a;
9678	:douta	=	16'h	7d5b;
9679	:douta	=	16'h	8ddc;
9680	:douta	=	16'h	855c;
9681	:douta	=	16'h	7d5b;
9682	:douta	=	16'h	7d3b;
9683	:douta	=	16'h	7d3b;
9684	:douta	=	16'h	753a;
9685	:douta	=	16'h	7d5b;
9686	:douta	=	16'h	7d5b;
9687	:douta	=	16'h	751a;
9688	:douta	=	16'h	8d9b;
9689	:douta	=	16'h	857b;
9690	:douta	=	16'h	6cda;
9691	:douta	=	16'h	6498;
9692	:douta	=	16'h	7d3b;
9693	:douta	=	16'h	7d5b;
9694	:douta	=	16'h	7d5b;
9695	:douta	=	16'h	74b9;
9696	:douta	=	16'h	74d9;
9697	:douta	=	16'h	74b9;
9698	:douta	=	16'h	7d3a;
9699	:douta	=	16'h	8d9c;
9700	:douta	=	16'h	74f9;
9701	:douta	=	16'h	6498;
9702	:douta	=	16'h	6499;
9703	:douta	=	16'h	6cda;
9704	:douta	=	16'h	7d3b;
9705	:douta	=	16'h	7d7b;
9706	:douta	=	16'h	7d3a;
9707	:douta	=	16'h	6cba;
9708	:douta	=	16'h	6bf6;
9709	:douta	=	16'h	2167;
9710	:douta	=	16'h	1968;
9711	:douta	=	16'h	21a9;
9712	:douta	=	16'h	21cb;
9713	:douta	=	16'h	7477;
9714	:douta	=	16'h	4352;
9715	:douta	=	16'h	32d2;
9716	:douta	=	16'h	8d5a;
9717	:douta	=	16'h	5bb4;
9718	:douta	=	16'h	9d9a;
9719	:douta	=	16'h	adba;
9720	:douta	=	16'h	7cd8;
9721	:douta	=	16'h	5bb4;
9722	:douta	=	16'h	959b;
9723	:douta	=	16'h	3290;
9724	:douta	=	16'h	5394;
9725	:douta	=	16'h	32b0;
9726	:douta	=	16'h	7c96;
9727	:douta	=	16'h	7c75;
9728	:douta	=	16'h	32f2;
9729	:douta	=	16'h	222e;
9730	:douta	=	16'h	32f1;
9731	:douta	=	16'h	5c37;
9732	:douta	=	16'h	53b4;
9733	:douta	=	16'h	6c98;
9734	:douta	=	16'h	6436;
9735	:douta	=	16'h	6c98;
9736	:douta	=	16'h	6c15;
9737	:douta	=	16'h	3a6e;
9738	:douta	=	16'h	4b11;
9739	:douta	=	16'h	4311;
9740	:douta	=	16'h	5b72;
9741	:douta	=	16'h	a537;
9742	:douta	=	16'h	94d6;
9743	:douta	=	16'h	9d17;
9744	:douta	=	16'h	73d3;
9745	:douta	=	16'h	73f2;
9746	:douta	=	16'h	8c95;
9747	:douta	=	16'h	ad98;
9748	:douta	=	16'h	6bd4;
9749	:douta	=	16'h	b595;
9750	:douta	=	16'h	d637;
9751	:douta	=	16'h	bdb6;
9752	:douta	=	16'h	8c73;
9753	:douta	=	16'h	ad54;
9754	:douta	=	16'h	73f2;
9755	:douta	=	16'h	7391;
9756	:douta	=	16'h	7c10;
9757	:douta	=	16'h	ad55;
9758	:douta	=	16'h	d657;
9759	:douta	=	16'h	de77;
9760	:douta	=	16'h	9cb2;
9761	:douta	=	16'h	8c10;
9762	:douta	=	16'h	b554;
9763	:douta	=	16'h	d636;
9764	:douta	=	16'h	83ef;
9765	:douta	=	16'h	ce16;
9766	:douta	=	16'h	c5f5;
9767	:douta	=	16'h	ef39;
9768	:douta	=	16'h	f75a;
9769	:douta	=	16'h	bd72;
9770	:douta	=	16'h	e676;
9771	:douta	=	16'h	c5d3;
9772	:douta	=	16'h	a48f;
9773	:douta	=	16'h	4a48;
9774	:douta	=	16'h	ef19;
9775	:douta	=	16'h	e6d8;
9776	:douta	=	16'h	b532;
9777	:douta	=	16'h	7bad;
9778	:douta	=	16'h	6289;
9779	:douta	=	16'h	d675;
9780	:douta	=	16'h	5aca;
9781	:douta	=	16'h	b570;
9782	:douta	=	16'h	83ab;
9783	:douta	=	16'h	730a;
9784	:douta	=	16'h	83ab;
9785	:douta	=	16'h	7b4b;
9786	:douta	=	16'h	6b2b;
9787	:douta	=	16'h	62c9;
9788	:douta	=	16'h	5a69;
9789	:douta	=	16'h	39e7;
9790	:douta	=	16'h	2986;
9791	:douta	=	16'h	10c4;
9792	:douta	=	16'h	2125;
9793	:douta	=	16'h	3187;
9794	:douta	=	16'h	10e5;
9795	:douta	=	16'h	10e4;
9796	:douta	=	16'h	10e5;
9797	:douta	=	16'h	2167;
9798	:douta	=	16'h	1126;
9799	:douta	=	16'h	10e5;
9800	:douta	=	16'h	0884;
9801	:douta	=	16'h	b4b1;
9802	:douta	=	16'h	42ab;
9803	:douta	=	16'h	4a29;
9804	:douta	=	16'h	7bad;
9805	:douta	=	16'h	5b2c;
9806	:douta	=	16'h	6b4e;
9807	:douta	=	16'h	5371;
9808	:douta	=	16'h	5b50;
9809	:douta	=	16'h	42ef;
9810	:douta	=	16'h	4a6b;
9811	:douta	=	16'h	6bf2;
9812	:douta	=	16'h	3a29;
9813	:douta	=	16'h	8c92;
9814	:douta	=	16'h	4a6a;
9815	:douta	=	16'h	ad33;
9816	:douta	=	16'h	1906;
9817	:douta	=	16'h	83ef;
9818	:douta	=	16'h	4b51;
9819	:douta	=	16'h	6371;
9820	:douta	=	16'h	3aae;
9821	:douta	=	16'h	8495;
9822	:douta	=	16'h	5bd3;
9823	:douta	=	16'h	3a6d;
9824	:douta	=	16'h	21ca;
9825	:douta	=	16'h	324d;
9826	:douta	=	16'h	3a09;
9827	:douta	=	16'h	1041;
9828	:douta	=	16'h	18a2;
9829	:douta	=	16'h	10a2;
9830	:douta	=	16'h	0861;
9831	:douta	=	16'h	0000;
9832	:douta	=	16'h	0000;
9833	:douta	=	16'h	4b0f;
9834	:douta	=	16'h	2a4e;
9835	:douta	=	16'h	32d1;
9836	:douta	=	16'h	1149;
9837	:douta	=	16'h	1989;
9838	:douta	=	16'h	53f5;
9839	:douta	=	16'h	53b3;
9840	:douta	=	16'h	53d5;
9841	:douta	=	16'h	42d1;
9842	:douta	=	16'h	5351;
9843	:douta	=	16'h	32d0;
9844	:douta	=	16'h	19ed;
9845	:douta	=	16'h	118b;
9846	:douta	=	16'h	63f4;
9847	:douta	=	16'h	7d1a;
9848	:douta	=	16'h	74b8;
9849	:douta	=	16'h	5c16;
9850	:douta	=	16'h	5c16;
9851	:douta	=	16'h	7d19;
9852	:douta	=	16'h	6cb9;
9853	:douta	=	16'h	52cd;
9854	:douta	=	16'h	422a;
9855	:douta	=	16'h	39c7;
9856	:douta	=	16'h	a42d;
9857	:douta	=	16'h	31a7;
9858	:douta	=	16'h	84d7;
9859	:douta	=	16'h	8d59;
9860	:douta	=	16'h	8497;
9861	:douta	=	16'h	7c97;
9862	:douta	=	16'h	8cd8;
9863	:douta	=	16'h	84f8;
9864	:douta	=	16'h	5bf5;
9865	:douta	=	16'h	6436;
9866	:douta	=	16'h	6c36;
9867	:douta	=	16'h	84f9;
9868	:douta	=	16'h	84f9;
9869	:douta	=	16'h	8d19;
9870	:douta	=	16'h	7c97;
9871	:douta	=	16'h	7c97;
9872	:douta	=	16'h	6c35;
9873	:douta	=	16'h	8d19;
9874	:douta	=	16'h	8d39;
9875	:douta	=	16'h	8d39;
9876	:douta	=	16'h	6c36;
9877	:douta	=	16'h	63f4;
9878	:douta	=	16'h	7c97;
9879	:douta	=	16'h	955a;
9880	:douta	=	16'h	8d7a;
9881	:douta	=	16'h	84f8;
9882	:douta	=	16'h	7c77;
9883	:douta	=	16'h	6c56;
9884	:douta	=	16'h	7c98;
9885	:douta	=	16'h	84f9;
9886	:douta	=	16'h	8519;
9887	:douta	=	16'h	8519;
9888	:douta	=	16'h	6c56;
9889	:douta	=	16'h	63d5;
9890	:douta	=	16'h	6c36;
9891	:douta	=	16'h	5bf5;
9892	:douta	=	16'h	6c57;
9893	:douta	=	16'h	7497;
9894	:douta	=	16'h	8d5a;
9895	:douta	=	16'h	8d7a;
9896	:douta	=	16'h	853a;
9897	:douta	=	16'h	8519;
9898	:douta	=	16'h	9dbc;
9899	:douta	=	16'h	8d5b;
9900	:douta	=	16'h	7cd9;
9901	:douta	=	16'h	95bc;
9902	:douta	=	16'h	959b;
9903	:douta	=	16'h	959c;
9904	:douta	=	16'h	95bc;
9905	:douta	=	16'h	8d5b;
9906	:douta	=	16'h	8d7b;
9907	:douta	=	16'h	853a;
9908	:douta	=	16'h	8d5a;
9909	:douta	=	16'h	853a;
9910	:douta	=	16'h	851a;
9911	:douta	=	16'h	8d5b;
9912	:douta	=	16'h	957b;
9913	:douta	=	16'h	8d7b;
9914	:douta	=	16'h	959b;
9915	:douta	=	16'h	959b;
9916	:douta	=	16'h	95bc;
9917	:douta	=	16'h	959b;
9918	:douta	=	16'h	7d19;
9919	:douta	=	16'h	8d5b;
9920	:douta	=	16'h	8d5a;
9921	:douta	=	16'h	95bc;
9922	:douta	=	16'h	8d9b;
9923	:douta	=	16'h	95bc;
9924	:douta	=	16'h	9ddc;
9925	:douta	=	16'h	6c79;
9926	:douta	=	16'h	7d3b;
9927	:douta	=	16'h	961d;
9928	:douta	=	16'h	6cba;
9929	:douta	=	16'h	859c;
9930	:douta	=	16'h	751b;
9931	:douta	=	16'h	6cba;
9932	:douta	=	16'h	7d3b;
9933	:douta	=	16'h	6cda;
9934	:douta	=	16'h	753b;
9935	:douta	=	16'h	7d5b;
9936	:douta	=	16'h	855c;
9937	:douta	=	16'h	8d9b;
9938	:douta	=	16'h	857c;
9939	:douta	=	16'h	74fa;
9940	:douta	=	16'h	74fa;
9941	:douta	=	16'h	857b;
9942	:douta	=	16'h	857b;
9943	:douta	=	16'h	74fa;
9944	:douta	=	16'h	751b;
9945	:douta	=	16'h	857b;
9946	:douta	=	16'h	857b;
9947	:douta	=	16'h	7d3b;
9948	:douta	=	16'h	6cba;
9949	:douta	=	16'h	753b;
9950	:douta	=	16'h	857c;
9951	:douta	=	16'h	7d3b;
9952	:douta	=	16'h	6c98;
9953	:douta	=	16'h	7d1a;
9954	:douta	=	16'h	74f9;
9955	:douta	=	16'h	855b;
9956	:douta	=	16'h	8dbc;
9957	:douta	=	16'h	855b;
9958	:douta	=	16'h	6499;
9959	:douta	=	16'h	6499;
9960	:douta	=	16'h	6478;
9961	:douta	=	16'h	755b;
9962	:douta	=	16'h	751b;
9963	:douta	=	16'h	7d7c;
9964	:douta	=	16'h	74fa;
9965	:douta	=	16'h	29aa;
9966	:douta	=	16'h	29ca;
9967	:douta	=	16'h	1968;
9968	:douta	=	16'h	1106;
9969	:douta	=	16'h	6c34;
9970	:douta	=	16'h	53d4;
9971	:douta	=	16'h	32d1;
9972	:douta	=	16'h	32d0;
9973	:douta	=	16'h	3b32;
9974	:douta	=	16'h	2ab1;
9975	:douta	=	16'h	adda;
9976	:douta	=	16'h	5bd4;
9977	:douta	=	16'h	9d79;
9978	:douta	=	16'h	8519;
9979	:douta	=	16'h	6435;
9980	:douta	=	16'h	63d4;
9981	:douta	=	16'h	7435;
9982	:douta	=	16'h	4353;
9983	:douta	=	16'h	322c;
9984	:douta	=	16'h	2ab0;
9985	:douta	=	16'h	32d2;
9986	:douta	=	16'h	4374;
9987	:douta	=	16'h	5c57;
9988	:douta	=	16'h	326f;
9989	:douta	=	16'h	4b32;
9990	:douta	=	16'h	4b52;
9991	:douta	=	16'h	5bd5;
9992	:douta	=	16'h	7c76;
9993	:douta	=	16'h	7c56;
9994	:douta	=	16'h	8497;
9995	:douta	=	16'h	9d59;
9996	:douta	=	16'h	84d7;
9997	:douta	=	16'h	7c12;
9998	:douta	=	16'h	4ad0;
9999	:douta	=	16'h	5b70;
10000	:douta	=	16'h	5b30;
10001	:douta	=	16'h	a516;
10002	:douta	=	16'h	a536;
10003	:douta	=	16'h	ce39;
10004	:douta	=	16'h	b5b8;
10005	:douta	=	16'h	a515;
10006	:douta	=	16'h	8c93;
10007	:douta	=	16'h	ad35;
10008	:douta	=	16'h	3a4d;
10009	:douta	=	16'h	8c52;
10010	:douta	=	16'h	c5f6;
10011	:douta	=	16'h	de77;
10012	:douta	=	16'h	ad75;
10013	:douta	=	16'h	8c72;
10014	:douta	=	16'h	ad56;
10015	:douta	=	16'h	6b4d;
10016	:douta	=	16'h	9cb2;
10017	:douta	=	16'h	8410;
10018	:douta	=	16'h	c5f6;
10019	:douta	=	16'h	de76;
10020	:douta	=	16'h	a4d1;
10021	:douta	=	16'h	ad33;
10022	:douta	=	16'h	8bf0;
10023	:douta	=	16'h	52ed;
10024	:douta	=	16'h	8c0f;
10025	:douta	=	16'h	9c90;
10026	:douta	=	16'h	9c6f;
10027	:douta	=	16'h	bdd3;
10028	:douta	=	16'h	de97;
10029	:douta	=	16'h	cdd3;
10030	:douta	=	16'h	a4d1;
10031	:douta	=	16'h	d636;
10032	:douta	=	16'h	736c;
10033	:douta	=	16'h	842e;
10034	:douta	=	16'h	c593;
10035	:douta	=	16'h	c614;
10036	:douta	=	16'h	b572;
10037	:douta	=	16'h	7b6c;
10038	:douta	=	16'h	836b;
10039	:douta	=	16'h	83ac;
10040	:douta	=	16'h	836b;
10041	:douta	=	16'h	7b4b;
10042	:douta	=	16'h	836b;
10043	:douta	=	16'h	62a9;
10044	:douta	=	16'h	5a68;
10045	:douta	=	16'h	4a49;
10046	:douta	=	16'h	31c8;
10047	:douta	=	16'h	2167;
10048	:douta	=	16'h	10c5;
10049	:douta	=	16'h	39a7;
10050	:douta	=	16'h	10a4;
10051	:douta	=	16'h	10e5;
10052	:douta	=	16'h	10a4;
10053	:douta	=	16'h	10e4;
10054	:douta	=	16'h	10e4;
10055	:douta	=	16'h	18e5;
10056	:douta	=	16'h	10e4;
10057	:douta	=	16'h	4229;
10058	:douta	=	16'h	31e9;
10059	:douta	=	16'h	39a8;
10060	:douta	=	16'h	9cf1;
10061	:douta	=	16'h	738d;
10062	:douta	=	16'h	63d1;
10063	:douta	=	16'h	63d2;
10064	:douta	=	16'h	6c33;
10065	:douta	=	16'h	5b0e;
10066	:douta	=	16'h	1927;
10067	:douta	=	16'h	1927;
10068	:douta	=	16'h	638e;
10069	:douta	=	16'h	530d;
10070	:douta	=	16'h	4a4a;
10071	:douta	=	16'h	8430;
10072	:douta	=	16'h	5acc;
10073	:douta	=	16'h	7bef;
10074	:douta	=	16'h	10e6;
10075	:douta	=	16'h	8474;
10076	:douta	=	16'h	3a8e;
10077	:douta	=	16'h	7c33;
10078	:douta	=	16'h	4b0f;
10079	:douta	=	16'h	5370;
10080	:douta	=	16'h	4b31;
10081	:douta	=	16'h	4b10;
10082	:douta	=	16'h	3a8f;
10083	:douta	=	16'h	5393;
10084	:douta	=	16'h	3aaf;
10085	:douta	=	16'h	0841;
10086	:douta	=	16'h	1081;
10087	:douta	=	16'h	10e3;
10088	:douta	=	16'h	18e4;
10089	:douta	=	16'h	1060;
10090	:douta	=	16'h	1926;
10091	:douta	=	16'h	428d;
10092	:douta	=	16'h	5330;
10093	:douta	=	16'h	220c;
10094	:douta	=	16'h	1169;
10095	:douta	=	16'h	4374;
10096	:douta	=	16'h	3b32;
10097	:douta	=	16'h	29ec;
10098	:douta	=	16'h	4b11;
10099	:douta	=	16'h	3b11;
10100	:douta	=	16'h	4312;
10101	:douta	=	16'h	4373;
10102	:douta	=	16'h	7cd8;
10103	:douta	=	16'h	53b4;
10104	:douta	=	16'h	74b8;
10105	:douta	=	16'h	198b;
10106	:douta	=	16'h	3a4e;
10107	:douta	=	16'h	6498;
10108	:douta	=	16'h	5372;
10109	:douta	=	16'h	4a4a;
10110	:douta	=	16'h	c48e;
10111	:douta	=	16'h	acaf;
10112	:douta	=	16'h	94b6;
10113	:douta	=	16'h	95bc;
10114	:douta	=	16'h	957b;
10115	:douta	=	16'h	6478;
10116	:douta	=	16'h	4bd6;
10117	:douta	=	16'h	7cd8;
10118	:douta	=	16'h	9dbb;
10119	:douta	=	16'h	957a;
10120	:douta	=	16'h	7498;
10121	:douta	=	16'h	6416;
10122	:douta	=	16'h	5bf5;
10123	:douta	=	16'h	5bb5;
10124	:douta	=	16'h	6c56;
10125	:douta	=	16'h	7457;
10126	:douta	=	16'h	7cb8;
10127	:douta	=	16'h	7c76;
10128	:douta	=	16'h	7476;
10129	:douta	=	16'h	7cb8;
10130	:douta	=	16'h	6415;
10131	:douta	=	16'h	6c36;
10132	:douta	=	16'h	5bd4;
10133	:douta	=	16'h	6415;
10134	:douta	=	16'h	95dc;
10135	:douta	=	16'h	8d1a;
10136	:douta	=	16'h	7cb8;
10137	:douta	=	16'h	84f9;
10138	:douta	=	16'h	8539;
10139	:douta	=	16'h	959b;
10140	:douta	=	16'h	84d8;
10141	:douta	=	16'h	7477;
10142	:douta	=	16'h	6c16;
10143	:douta	=	16'h	7cb8;
10144	:douta	=	16'h	84d8;
10145	:douta	=	16'h	7497;
10146	:douta	=	16'h	6415;
10147	:douta	=	16'h	6c56;
10148	:douta	=	16'h	63f5;
10149	:douta	=	16'h	7478;
10150	:douta	=	16'h	7cf9;
10151	:douta	=	16'h	851a;
10152	:douta	=	16'h	853a;
10153	:douta	=	16'h	7cd8;
10154	:douta	=	16'h	8d5a;
10155	:douta	=	16'h	8d7a;
10156	:douta	=	16'h	853a;
10157	:douta	=	16'h	8d3b;
10158	:douta	=	16'h	851a;
10159	:douta	=	16'h	7cd9;
10160	:douta	=	16'h	853a;
10161	:douta	=	16'h	959c;
10162	:douta	=	16'h	9ddc;
10163	:douta	=	16'h	8d5a;
10164	:douta	=	16'h	7cd9;
10165	:douta	=	16'h	7d19;
10166	:douta	=	16'h	8d3a;
10167	:douta	=	16'h	8d3a;
10168	:douta	=	16'h	8d5a;
10169	:douta	=	16'h	851a;
10170	:douta	=	16'h	8d7b;
10171	:douta	=	16'h	8d3a;
10172	:douta	=	16'h	8d7b;
10173	:douta	=	16'h	853a;
10174	:douta	=	16'h	8d3a;
10175	:douta	=	16'h	8d5b;
10176	:douta	=	16'h	959b;
10177	:douta	=	16'h	7cf9;
10178	:douta	=	16'h	851a;
10179	:douta	=	16'h	851a;
10180	:douta	=	16'h	853a;
10181	:douta	=	16'h	8d7b;
10182	:douta	=	16'h	8d7b;
10183	:douta	=	16'h	855a;
10184	:douta	=	16'h	855c;
10185	:douta	=	16'h	6499;
10186	:douta	=	16'h	5417;
10187	:douta	=	16'h	8e1e;
10188	:douta	=	16'h	9e3e;
10189	:douta	=	16'h	6478;
10190	:douta	=	16'h	5c58;
10191	:douta	=	16'h	6cfa;
10192	:douta	=	16'h	6cba;
10193	:douta	=	16'h	74da;
10194	:douta	=	16'h	7d3b;
10195	:douta	=	16'h	857c;
10196	:douta	=	16'h	7d3b;
10197	:douta	=	16'h	751a;
10198	:douta	=	16'h	7d1a;
10199	:douta	=	16'h	857b;
10200	:douta	=	16'h	857b;
10201	:douta	=	16'h	74d9;
10202	:douta	=	16'h	74ba;
10203	:douta	=	16'h	74fa;
10204	:douta	=	16'h	7d3a;
10205	:douta	=	16'h	751a;
10206	:douta	=	16'h	6cb9;
10207	:douta	=	16'h	6458;
10208	:douta	=	16'h	74da;
10209	:douta	=	16'h	859b;
10210	:douta	=	16'h	74f9;
10211	:douta	=	16'h	8d5b;
10212	:douta	=	16'h	7d3b;
10213	:douta	=	16'h	6c98;
10214	:douta	=	16'h	6cd9;
10215	:douta	=	16'h	6cfa;
10216	:douta	=	16'h	7d5c;
10217	:douta	=	16'h	6478;
10218	:douta	=	16'h	5c58;
10219	:douta	=	16'h	74fa;
10220	:douta	=	16'h	7d3b;
10221	:douta	=	16'h	751b;
10222	:douta	=	16'h	31ea;
10223	:douta	=	16'h	1906;
10224	:douta	=	16'h	2989;
10225	:douta	=	16'h	1107;
10226	:douta	=	16'h	957a;
10227	:douta	=	16'h	5353;
10228	:douta	=	16'h	9559;
10229	:douta	=	16'h	7497;
10230	:douta	=	16'h	9d7a;
10231	:douta	=	16'h	19cc;
10232	:douta	=	16'h	84d7;
10233	:douta	=	16'h	32d0;
10234	:douta	=	16'h	3290;
10235	:douta	=	16'h	4b51;
10236	:douta	=	16'h	7433;
10237	:douta	=	16'h	7c75;
10238	:douta	=	16'h	a597;
10239	:douta	=	16'h	42d0;
10240	:douta	=	16'h	3b53;
10241	:douta	=	16'h	32d1;
10242	:douta	=	16'h	32d1;
10243	:douta	=	16'h	74fa;
10244	:douta	=	16'h	5373;
10245	:douta	=	16'h	6c77;
10246	:douta	=	16'h	5bb4;
10247	:douta	=	16'h	6436;
10248	:douta	=	16'h	5373;
10249	:douta	=	16'h	428f;
10250	:douta	=	16'h	5351;
10251	:douta	=	16'h	8cf8;
10252	:douta	=	16'h	7c96;
10253	:douta	=	16'h	94b6;
10254	:douta	=	16'h	9d16;
10255	:douta	=	16'h	9cf5;
10256	:douta	=	16'h	6392;
10257	:douta	=	16'h	9cd6;
10258	:douta	=	16'h	8c94;
10259	:douta	=	16'h	bdf9;
10260	:douta	=	16'h	8454;
10261	:douta	=	16'h	d659;
10262	:douta	=	16'h	ce38;
10263	:douta	=	16'h	cdf6;
10264	:douta	=	16'h	8c53;
10265	:douta	=	16'h	6b70;
10266	:douta	=	16'h	ad55;
10267	:douta	=	16'h	ad34;
10268	:douta	=	16'h	9cd3;
10269	:douta	=	16'h	b555;
10270	:douta	=	16'h	d637;
10271	:douta	=	16'h	ee98;
10272	:douta	=	16'h	ef39;
10273	:douta	=	16'h	8410;
10274	:douta	=	16'h	83ef;
10275	:douta	=	16'h	c5d4;
10276	:douta	=	16'h	b593;
10277	:douta	=	16'h	ad32;
10278	:douta	=	16'h	eed8;
10279	:douta	=	16'h	bd52;
10280	:douta	=	16'h	e697;
10281	:douta	=	16'h	6b4c;
10282	:douta	=	16'h	6269;
10283	:douta	=	16'h	8cd1;
10284	:douta	=	16'h	cdf3;
10285	:douta	=	16'h	8c6f;
10286	:douta	=	16'h	eef8;
10287	:douta	=	16'h	deb7;
10288	:douta	=	16'h	c592;
10289	:douta	=	16'h	738c;
10290	:douta	=	16'h	ac91;
10291	:douta	=	16'h	94cf;
10292	:douta	=	16'h	736c;
10293	:douta	=	16'h	7b2b;
10294	:douta	=	16'h	8b8c;
10295	:douta	=	16'h	8bac;
10296	:douta	=	16'h	838b;
10297	:douta	=	16'h	838c;
10298	:douta	=	16'h	7b2a;
10299	:douta	=	16'h	62a9;
10300	:douta	=	16'h	4a49;
10301	:douta	=	16'h	4a29;
10302	:douta	=	16'h	4a6b;
10303	:douta	=	16'h	320a;
10304	:douta	=	16'h	29a8;
10305	:douta	=	16'h	31a7;
10306	:douta	=	16'h	1905;
10307	:douta	=	16'h	10e4;
10308	:douta	=	16'h	18e5;
10309	:douta	=	16'h	08a4;
10310	:douta	=	16'h	10c4;
10311	:douta	=	16'h	1105;
10312	:douta	=	16'h	10e4;
10313	:douta	=	16'h	4208;
10314	:douta	=	16'h	4a8a;
10315	:douta	=	16'h	528a;
10316	:douta	=	16'h	8c70;
10317	:douta	=	16'h	6b2b;
10318	:douta	=	16'h	63b1;
10319	:douta	=	16'h	63d2;
10320	:douta	=	16'h	5b6f;
10321	:douta	=	16'h	636e;
10322	:douta	=	16'h	7bae;
10323	:douta	=	16'h	2189;
10324	:douta	=	16'h	73d0;
10325	:douta	=	16'h	52cd;
10326	:douta	=	16'h	2189;
10327	:douta	=	16'h	3209;
10328	:douta	=	16'h	528b;
10329	:douta	=	16'h	6b8e;
10330	:douta	=	16'h	29aa;
10331	:douta	=	16'h	6bf1;
10332	:douta	=	16'h	2a2c;
10333	:douta	=	16'h	7453;
10334	:douta	=	16'h	5371;
10335	:douta	=	16'h	6391;
10336	:douta	=	16'h	21cb;
10337	:douta	=	16'h	428d;
10338	:douta	=	16'h	5330;
10339	:douta	=	16'h	63d2;
10340	:douta	=	16'h	53f6;
10341	:douta	=	16'h	4ace;
10342	:douta	=	16'h	2986;
10343	:douta	=	16'h	10a3;
10344	:douta	=	16'h	18e4;
10345	:douta	=	16'h	18c4;
10346	:douta	=	16'h	0841;
10347	:douta	=	16'h	0021;
10348	:douta	=	16'h	4aef;
10349	:douta	=	16'h	6393;
10350	:douta	=	16'h	00a6;
10351	:douta	=	16'h	2a8f;
10352	:douta	=	16'h	4311;
10353	:douta	=	16'h	4311;
10354	:douta	=	16'h	5bd5;
10355	:douta	=	16'h	3b32;
10356	:douta	=	16'h	00e9;
10357	:douta	=	16'h	118c;
10358	:douta	=	16'h	4b32;
10359	:douta	=	16'h	3af1;
10360	:douta	=	16'h	6497;
10361	:douta	=	16'h	4b11;
10362	:douta	=	16'h	6436;
10363	:douta	=	16'h	5bd4;
10364	:douta	=	16'h	5228;
10365	:douta	=	16'h	41e9;
10366	:douta	=	16'h	acce;
10367	:douta	=	16'h	41e8;
10368	:douta	=	16'h	9ddd;
10369	:douta	=	16'h	853b;
10370	:douta	=	16'h	8d5b;
10371	:douta	=	16'h	8d7b;
10372	:douta	=	16'h	7cd9;
10373	:douta	=	16'h	6c78;
10374	:douta	=	16'h	7498;
10375	:douta	=	16'h	959b;
10376	:douta	=	16'h	9ddc;
10377	:douta	=	16'h	8d3a;
10378	:douta	=	16'h	6c36;
10379	:douta	=	16'h	5bd5;
10380	:douta	=	16'h	6c57;
10381	:douta	=	16'h	7477;
10382	:douta	=	16'h	8d39;
10383	:douta	=	16'h	84f9;
10384	:douta	=	16'h	7cb8;
10385	:douta	=	16'h	8519;
10386	:douta	=	16'h	84d8;
10387	:douta	=	16'h	8d19;
10388	:douta	=	16'h	7c98;
10389	:douta	=	16'h	6415;
10390	:douta	=	16'h	6c36;
10391	:douta	=	16'h	9ddb;
10392	:douta	=	16'h	a61c;
10393	:douta	=	16'h	84f9;
10394	:douta	=	16'h	7cb8;
10395	:douta	=	16'h	84d9;
10396	:douta	=	16'h	8d5a;
10397	:douta	=	16'h	959b;
10398	:douta	=	16'h	84d8;
10399	:douta	=	16'h	7cb8;
10400	:douta	=	16'h	7477;
10401	:douta	=	16'h	84d8;
10402	:douta	=	16'h	7cd8;
10403	:douta	=	16'h	7457;
10404	:douta	=	16'h	63f5;
10405	:douta	=	16'h	7cb8;
10406	:douta	=	16'h	6416;
10407	:douta	=	16'h	6c57;
10408	:douta	=	16'h	8519;
10409	:douta	=	16'h	7cd8;
10410	:douta	=	16'h	8519;
10411	:douta	=	16'h	8539;
10412	:douta	=	16'h	8519;
10413	:douta	=	16'h	7498;
10414	:douta	=	16'h	8519;
10415	:douta	=	16'h	7cf9;
10416	:douta	=	16'h	7cf9;
10417	:douta	=	16'h	7d19;
10418	:douta	=	16'h	8d5b;
10419	:douta	=	16'h	9ddc;
10420	:douta	=	16'h	959b;
10421	:douta	=	16'h	853a;
10422	:douta	=	16'h	851a;
10423	:douta	=	16'h	8519;
10424	:douta	=	16'h	957a;
10425	:douta	=	16'h	957b;
10426	:douta	=	16'h	851a;
10427	:douta	=	16'h	957b;
10428	:douta	=	16'h	8d3a;
10429	:douta	=	16'h	8d7b;
10430	:douta	=	16'h	8519;
10431	:douta	=	16'h	8d3a;
10432	:douta	=	16'h	8d7b;
10433	:douta	=	16'h	8d7b;
10434	:douta	=	16'h	8d5b;
10435	:douta	=	16'h	851a;
10436	:douta	=	16'h	851a;
10437	:douta	=	16'h	8d9b;
10438	:douta	=	16'h	8d5b;
10439	:douta	=	16'h	8d7c;
10440	:douta	=	16'h	959c;
10441	:douta	=	16'h	95bc;
10442	:douta	=	16'h	53d7;
10443	:douta	=	16'h	4bd6;
10444	:douta	=	16'h	751a;
10445	:douta	=	16'h	ae7e;
10446	:douta	=	16'h	8d9c;
10447	:douta	=	16'h	6cfa;
10448	:douta	=	16'h	6cda;
10449	:douta	=	16'h	6cba;
10450	:douta	=	16'h	7d5b;
10451	:douta	=	16'h	859c;
10452	:douta	=	16'h	6cda;
10453	:douta	=	16'h	7d5b;
10454	:douta	=	16'h	855b;
10455	:douta	=	16'h	857b;
10456	:douta	=	16'h	855b;
10457	:douta	=	16'h	855b;
10458	:douta	=	16'h	6478;
10459	:douta	=	16'h	74b9;
10460	:douta	=	16'h	751a;
10461	:douta	=	16'h	74fa;
10462	:douta	=	16'h	74d9;
10463	:douta	=	16'h	74d9;
10464	:douta	=	16'h	74b9;
10465	:douta	=	16'h	7d3a;
10466	:douta	=	16'h	8dbc;
10467	:douta	=	16'h	8dbc;
10468	:douta	=	16'h	8d9c;
10469	:douta	=	16'h	855b;
10470	:douta	=	16'h	751a;
10471	:douta	=	16'h	6cd9;
10472	:douta	=	16'h	859b;
10473	:douta	=	16'h	7d7c;
10474	:douta	=	16'h	74fb;
10475	:douta	=	16'h	6478;
10476	:douta	=	16'h	6457;
10477	:douta	=	16'h	74f9;
10478	:douta	=	16'h	7457;
10479	:douta	=	16'h	29a9;
10480	:douta	=	16'h	2189;
10481	:douta	=	16'h	2989;
10482	:douta	=	16'h	2a8f;
10483	:douta	=	16'h	4b51;
10484	:douta	=	16'h	6c15;
10485	:douta	=	16'h	9d9a;
10486	:douta	=	16'h	ae1c;
10487	:douta	=	16'h	7435;
10488	:douta	=	16'h	84d7;
10489	:douta	=	16'h	4312;
10490	:douta	=	16'h	5393;
10491	:douta	=	16'h	0969;
10492	:douta	=	16'h	3a8d;
10493	:douta	=	16'h	324e;
10494	:douta	=	16'h	326e;
10495	:douta	=	16'h	6371;
10496	:douta	=	16'h	2ad1;
10497	:douta	=	16'h	4353;
10498	:douta	=	16'h	4374;
10499	:douta	=	16'h	6c99;
10500	:douta	=	16'h	4b53;
10501	:douta	=	16'h	324f;
10502	:douta	=	16'h	5bd5;
10503	:douta	=	16'h	4311;
10504	:douta	=	16'h	5373;
10505	:douta	=	16'h	6bd4;
10506	:douta	=	16'h	7c77;
10507	:douta	=	16'h	84d7;
10508	:douta	=	16'h	6c35;
10509	:douta	=	16'h	530f;
10510	:douta	=	16'h	4b0f;
10511	:douta	=	16'h	530f;
10512	:douta	=	16'h	8453;
10513	:douta	=	16'h	bd96;
10514	:douta	=	16'h	c639;
10515	:douta	=	16'h	d69a;
10516	:douta	=	16'h	bdf9;
10517	:douta	=	16'h	9c94;
10518	:douta	=	16'h	bdb7;
10519	:douta	=	16'h	6b8f;
10520	:douta	=	16'h	528b;
10521	:douta	=	16'h	bd95;
10522	:douta	=	16'h	c5d6;
10523	:douta	=	16'h	de78;
10524	:douta	=	16'h	b575;
10525	:douta	=	16'h	9cb3;
10526	:douta	=	16'h	d677;
10527	:douta	=	16'h	7bae;
10528	:douta	=	16'h	c594;
10529	:douta	=	16'h	632d;
10530	:douta	=	16'h	c5f6;
10531	:douta	=	16'h	b573;
10532	:douta	=	16'h	9cb1;
10533	:douta	=	16'h	acf2;
10534	:douta	=	16'h	6b0c;
10535	:douta	=	16'h	9491;
10536	:douta	=	16'h	bd73;
10537	:douta	=	16'h	83ed;
10538	:douta	=	16'h	9c6f;
10539	:douta	=	16'h	b572;
10540	:douta	=	16'h	ef39;
10541	:douta	=	16'h	bd93;
10542	:douta	=	16'h	ce14;
10543	:douta	=	16'h	deb7;
10544	:douta	=	16'h	8c0e;
10545	:douta	=	16'h	944e;
10546	:douta	=	16'h	bdd4;
10547	:douta	=	16'h	838b;
10548	:douta	=	16'h	836b;
10549	:douta	=	16'h	8bac;
10550	:douta	=	16'h	836b;
10551	:douta	=	16'h	8bcb;
10552	:douta	=	16'h	93cc;
10553	:douta	=	16'h	93ec;
10554	:douta	=	16'h	836b;
10555	:douta	=	16'h	62a9;
10556	:douta	=	16'h	4208;
10557	:douta	=	16'h	2147;
10558	:douta	=	16'h	2125;
10559	:douta	=	16'h	2946;
10560	:douta	=	16'h	2126;
10561	:douta	=	16'h	2126;
10562	:douta	=	16'h	3a28;
10563	:douta	=	16'h	10a4;
10564	:douta	=	16'h	10e5;
10565	:douta	=	16'h	10e5;
10566	:douta	=	16'h	10e5;
10567	:douta	=	16'h	10e4;
10568	:douta	=	16'h	18e5;
10569	:douta	=	16'h	10a4;
10570	:douta	=	16'h	2147;
10571	:douta	=	16'h	528a;
10572	:douta	=	16'h	7bac;
10573	:douta	=	16'h	8c2e;
10574	:douta	=	16'h	6bf3;
10575	:douta	=	16'h	5b71;
10576	:douta	=	16'h	6b8e;
10577	:douta	=	16'h	322b;
10578	:douta	=	16'h	3a2b;
10579	:douta	=	16'h	1988;
10580	:douta	=	16'h	738e;
10581	:douta	=	16'h	426b;
10582	:douta	=	16'h	9cb1;
10583	:douta	=	16'h	4acd;
10584	:douta	=	16'h	734d;
10585	:douta	=	16'h	9cf3;
10586	:douta	=	16'h	420a;
10587	:douta	=	16'h	08c6;
10588	:douta	=	16'h	18e6;
10589	:douta	=	16'h	6bb1;
10590	:douta	=	16'h	5b70;
10591	:douta	=	16'h	4b0f;
10592	:douta	=	16'h	530f;
10593	:douta	=	16'h	5b71;
10594	:douta	=	16'h	328e;
10595	:douta	=	16'h	5bb2;
10596	:douta	=	16'h	328f;
10597	:douta	=	16'h	2a0c;
10598	:douta	=	16'h	42f0;
10599	:douta	=	16'h	5b70;
10600	:douta	=	16'h	2168;
10601	:douta	=	16'h	10c2;
10602	:douta	=	16'h	18e3;
10603	:douta	=	16'h	10c4;
10604	:douta	=	16'h	0000;
10605	:douta	=	16'h	0000;
10606	:douta	=	16'h	428d;
10607	:douta	=	16'h	320c;
10608	:douta	=	16'h	0908;
10609	:douta	=	16'h	32af;
10610	:douta	=	16'h	32f1;
10611	:douta	=	16'h	3333;
10612	:douta	=	16'h	6457;
10613	:douta	=	16'h	6415;
10614	:douta	=	16'h	5c16;
10615	:douta	=	16'h	5394;
10616	:douta	=	16'h	4b93;
10617	:douta	=	16'h	4310;
10618	:douta	=	16'h	4aef;
10619	:douta	=	16'h	5a6a;
10620	:douta	=	16'h	39c9;
10621	:douta	=	16'h	c54f;
10622	:douta	=	16'h	8454;
10623	:douta	=	16'h	ae5e;
10624	:douta	=	16'h	8d5a;
10625	:douta	=	16'h	959b;
10626	:douta	=	16'h	959b;
10627	:douta	=	16'h	959b;
10628	:douta	=	16'h	959b;
10629	:douta	=	16'h	8519;
10630	:douta	=	16'h	959b;
10631	:douta	=	16'h	957a;
10632	:douta	=	16'h	8d5b;
10633	:douta	=	16'h	959c;
10634	:douta	=	16'h	8d7b;
10635	:douta	=	16'h	959b;
10636	:douta	=	16'h	9ddc;
10637	:douta	=	16'h	7cf8;
10638	:douta	=	16'h	7497;
10639	:douta	=	16'h	7cd8;
10640	:douta	=	16'h	7497;
10641	:douta	=	16'h	7498;
10642	:douta	=	16'h	7cd9;
10643	:douta	=	16'h	7cb8;
10644	:douta	=	16'h	7477;
10645	:douta	=	16'h	7478;
10646	:douta	=	16'h	8d7b;
10647	:douta	=	16'h	84d9;
10648	:douta	=	16'h	7c98;
10649	:douta	=	16'h	851a;
10650	:douta	=	16'h	95ba;
10651	:douta	=	16'h	957a;
10652	:douta	=	16'h	8d3a;
10653	:douta	=	16'h	6c35;
10654	:douta	=	16'h	7cb7;
10655	:douta	=	16'h	8d5a;
10656	:douta	=	16'h	9dbb;
10657	:douta	=	16'h	7cd8;
10658	:douta	=	16'h	6416;
10659	:douta	=	16'h	8d3a;
10660	:douta	=	16'h	9559;
10661	:douta	=	16'h	84f9;
10662	:douta	=	16'h	74d8;
10663	:douta	=	16'h	6435;
10664	:douta	=	16'h	5bd5;
10665	:douta	=	16'h	6c16;
10666	:douta	=	16'h	6c36;
10667	:douta	=	16'h	7477;
10668	:douta	=	16'h	7cd9;
10669	:douta	=	16'h	9ddc;
10670	:douta	=	16'h	8d5b;
10671	:douta	=	16'h	7cf9;
10672	:douta	=	16'h	95bc;
10673	:douta	=	16'h	959c;
10674	:douta	=	16'h	8d7b;
10675	:douta	=	16'h	853a;
10676	:douta	=	16'h	853a;
10677	:douta	=	16'h	855a;
10678	:douta	=	16'h	9dbc;
10679	:douta	=	16'h	95bc;
10680	:douta	=	16'h	8d7b;
10681	:douta	=	16'h	8519;
10682	:douta	=	16'h	8d7b;
10683	:douta	=	16'h	8519;
10684	:douta	=	16'h	7cd9;
10685	:douta	=	16'h	8d5a;
10686	:douta	=	16'h	95bc;
10687	:douta	=	16'h	959b;
10688	:douta	=	16'h	959b;
10689	:douta	=	16'h	8d5b;
10690	:douta	=	16'h	853a;
10691	:douta	=	16'h	8d5a;
10692	:douta	=	16'h	8d5b;
10693	:douta	=	16'h	853b;
10694	:douta	=	16'h	8d9c;
10695	:douta	=	16'h	959c;
10696	:douta	=	16'h	855b;
10697	:douta	=	16'h	855b;
10698	:douta	=	16'h	8d9c;
10699	:douta	=	16'h	959c;
10700	:douta	=	16'h	6c77;
10701	:douta	=	16'h	1a2f;
10702	:douta	=	16'h	3374;
10703	:douta	=	16'h	85bd;
10704	:douta	=	16'h	6cda;
10705	:douta	=	16'h	6cda;
10706	:douta	=	16'h	6c99;
10707	:douta	=	16'h	6c99;
10708	:douta	=	16'h	751a;
10709	:douta	=	16'h	74fa;
10710	:douta	=	16'h	751a;
10711	:douta	=	16'h	751a;
10712	:douta	=	16'h	857b;
10713	:douta	=	16'h	855b;
10714	:douta	=	16'h	8d9c;
10715	:douta	=	16'h	855b;
10716	:douta	=	16'h	6cb9;
10717	:douta	=	16'h	6cd9;
10718	:douta	=	16'h	74fa;
10719	:douta	=	16'h	7d3a;
10720	:douta	=	16'h	7d1a;
10721	:douta	=	16'h	7d3a;
10722	:douta	=	16'h	74d9;
10723	:douta	=	16'h	7d3a;
10724	:douta	=	16'h	8d9b;
10725	:douta	=	16'h	857b;
10726	:douta	=	16'h	74fa;
10727	:douta	=	16'h	95bc;
10728	:douta	=	16'h	8ddc;
10729	:douta	=	16'h	6c99;
10730	:douta	=	16'h	74fa;
10731	:douta	=	16'h	74da;
10732	:douta	=	16'h	7d7c;
10733	:douta	=	16'h	6c57;
10734	:douta	=	16'h	6436;
10735	:douta	=	16'h	7498;
10736	:douta	=	16'h	10e6;
10737	:douta	=	16'h	2168;
10738	:douta	=	16'h	1105;
10739	:douta	=	16'h	a5fc;
10740	:douta	=	16'h	7499;
10741	:douta	=	16'h	63f4;
10742	:douta	=	16'h	63b3;
10743	:douta	=	16'h	7496;
10744	:douta	=	16'h	5371;
10745	:douta	=	16'h	b5f8;
10746	:douta	=	16'h	4b31;
10747	:douta	=	16'h	7c33;
10748	:douta	=	16'h	6bf3;
10749	:douta	=	16'h	6416;
10750	:douta	=	16'h	326e;
10751	:douta	=	16'h	324e;
10752	:douta	=	16'h	3312;
10753	:douta	=	16'h	11cd;
10754	:douta	=	16'h	2a4f;
10755	:douta	=	16'h	4312;
10756	:douta	=	16'h	5bf5;
10757	:douta	=	16'h	5bd5;
10758	:douta	=	16'h	7cf9;
10759	:douta	=	16'h	4b53;
10760	:douta	=	16'h	5393;
10761	:douta	=	16'h	5310;
10762	:douta	=	16'h	5b72;
10763	:douta	=	16'h	84d7;
10764	:douta	=	16'h	7c96;
10765	:douta	=	16'h	8474;
10766	:douta	=	16'h	94b5;
10767	:douta	=	16'h	73f2;
10768	:douta	=	16'h	73f2;
10769	:douta	=	16'h	8c94;
10770	:douta	=	16'h	94d5;
10771	:douta	=	16'h	adb7;
10772	:douta	=	16'h	8c94;
10773	:douta	=	16'h	bdb6;
10774	:douta	=	16'h	c5d6;
10775	:douta	=	16'h	b554;
10776	:douta	=	16'h	6b70;
10777	:douta	=	16'h	83f1;
10778	:douta	=	16'h	b535;
10779	:douta	=	16'h	bdd6;
10780	:douta	=	16'h	9cd3;
10781	:douta	=	16'h	9cb2;
10782	:douta	=	16'h	ce36;
10783	:douta	=	16'h	c574;
10784	:douta	=	16'h	f6d8;
10785	:douta	=	16'h	52ad;
10786	:douta	=	16'h	736e;
10787	:douta	=	16'h	83d0;
10788	:douta	=	16'h	ad32;
10789	:douta	=	16'h	acf2;
10790	:douta	=	16'h	d636;
10791	:douta	=	16'h	a4d1;
10792	:douta	=	16'h	c593;
10793	:douta	=	16'h	6b4c;
10794	:douta	=	16'h	6aeb;
10795	:douta	=	16'h	532c;
10796	:douta	=	16'h	b551;
10797	:douta	=	16'h	9caf;
10798	:douta	=	16'h	f718;
10799	:douta	=	16'h	ef39;
10800	:douta	=	16'h	9caf;
10801	:douta	=	16'h	94b0;
10802	:douta	=	16'h	7b8c;
10803	:douta	=	16'h	8b8c;
10804	:douta	=	16'h	838c;
10805	:douta	=	16'h	8bac;
10806	:douta	=	16'h	836b;
10807	:douta	=	16'h	8bcc;
10808	:douta	=	16'h	93cc;
10809	:douta	=	16'h	8bab;
10810	:douta	=	16'h	8bac;
10811	:douta	=	16'h	5248;
10812	:douta	=	16'h	31a7;
10813	:douta	=	16'h	2126;
10814	:douta	=	16'h	18e5;
10815	:douta	=	16'h	2146;
10816	:douta	=	16'h	1906;
10817	:douta	=	16'h	10a4;
10818	:douta	=	16'h	3a08;
10819	:douta	=	16'h	10c5;
10820	:douta	=	16'h	10e5;
10821	:douta	=	16'h	10e4;
10822	:douta	=	16'h	10e5;
10823	:douta	=	16'h	10c4;
10824	:douta	=	16'h	10e5;
10825	:douta	=	16'h	10c4;
10826	:douta	=	16'h	39c8;
10827	:douta	=	16'h	2125;
10828	:douta	=	16'h	9c8f;
10829	:douta	=	16'h	9c91;
10830	:douta	=	16'h	5b72;
10831	:douta	=	16'h	5b71;
10832	:douta	=	16'h	9cb0;
10833	:douta	=	16'h	52cc;
10834	:douta	=	16'h	6b6e;
10835	:douta	=	16'h	1107;
10836	:douta	=	16'h	4acd;
10837	:douta	=	16'h	0085;
10838	:douta	=	16'h	73cf;
10839	:douta	=	16'h	4aac;
10840	:douta	=	16'h	5aec;
10841	:douta	=	16'h	8430;
10842	:douta	=	16'h	6b6e;
10843	:douta	=	16'h	29ca;
10844	:douta	=	16'h	52ac;
10845	:douta	=	16'h	5b4e;
10846	:douta	=	16'h	4acd;
10847	:douta	=	16'h	426d;
10848	:douta	=	16'h	5b4f;
10849	:douta	=	16'h	7c12;
10850	:douta	=	16'h	5bb3;
10851	:douta	=	16'h	6c14;
10852	:douta	=	16'h	4373;
10853	:douta	=	16'h	63f3;
10854	:douta	=	16'h	4b11;
10855	:douta	=	16'h	2a2d;
10856	:douta	=	16'h	2a2e;
10857	:douta	=	16'h	18e5;
10858	:douta	=	16'h	1061;
10859	:douta	=	16'h	1082;
10860	:douta	=	16'h	0001;
10861	:douta	=	16'h	0000;
10862	:douta	=	16'h	0000;
10863	:douta	=	16'h	5b50;
10864	:douta	=	16'h	4aef;
10865	:douta	=	16'h	32f1;
10866	:douta	=	16'h	224f;
10867	:douta	=	16'h	222d;
10868	:douta	=	16'h	5bb4;
10869	:douta	=	16'h	6c77;
10870	:douta	=	16'h	2a8f;
10871	:douta	=	16'h	326f;
10872	:douta	=	16'h	53f5;
10873	:douta	=	16'h	5394;
10874	:douta	=	16'h	5b50;
10875	:douta	=	16'h	39e9;
10876	:douta	=	16'h	830a;
10877	:douta	=	16'h	4a6a;
10878	:douta	=	16'h	9dfd;
10879	:douta	=	16'h	9ddc;
10880	:douta	=	16'h	8d7a;
10881	:douta	=	16'h	8d5a;
10882	:douta	=	16'h	959b;
10883	:douta	=	16'h	a5dc;
10884	:douta	=	16'h	a5fc;
10885	:douta	=	16'h	853a;
10886	:douta	=	16'h	8519;
10887	:douta	=	16'h	7cf9;
10888	:douta	=	16'h	853a;
10889	:douta	=	16'h	7cf9;
10890	:douta	=	16'h	8d7b;
10891	:douta	=	16'h	957b;
10892	:douta	=	16'h	8d7b;
10893	:douta	=	16'h	8d7a;
10894	:douta	=	16'h	8519;
10895	:douta	=	16'h	8d3a;
10896	:douta	=	16'h	8519;
10897	:douta	=	16'h	8519;
10898	:douta	=	16'h	7497;
10899	:douta	=	16'h	84f8;
10900	:douta	=	16'h	8519;
10901	:douta	=	16'h	7cd9;
10902	:douta	=	16'h	8d5a;
10903	:douta	=	16'h	74b8;
10904	:douta	=	16'h	855a;
10905	:douta	=	16'h	7498;
10906	:douta	=	16'h	7cd9;
10907	:douta	=	16'h	853a;
10908	:douta	=	16'h	95bb;
10909	:douta	=	16'h	8d59;
10910	:douta	=	16'h	6c15;
10911	:douta	=	16'h	7476;
10912	:douta	=	16'h	8d5a;
10913	:douta	=	16'h	95ba;
10914	:douta	=	16'h	8519;
10915	:douta	=	16'h	7478;
10916	:douta	=	16'h	7498;
10917	:douta	=	16'h	8d5a;
10918	:douta	=	16'h	8d5a;
10919	:douta	=	16'h	8d5a;
10920	:douta	=	16'h	7457;
10921	:douta	=	16'h	63f5;
10922	:douta	=	16'h	7cb8;
10923	:douta	=	16'h	7cf9;
10924	:douta	=	16'h	6c36;
10925	:douta	=	16'h	8519;
10926	:douta	=	16'h	959b;
10927	:douta	=	16'h	8d7b;
10928	:douta	=	16'h	8d7b;
10929	:douta	=	16'h	8519;
10930	:douta	=	16'h	8d7b;
10931	:douta	=	16'h	8d7b;
10932	:douta	=	16'h	8d7b;
10933	:douta	=	16'h	7cd9;
10934	:douta	=	16'h	9ddc;
10935	:douta	=	16'h	95bb;
10936	:douta	=	16'h	8d7b;
10937	:douta	=	16'h	957b;
10938	:douta	=	16'h	8d3a;
10939	:douta	=	16'h	957b;
10940	:douta	=	16'h	74b8;
10941	:douta	=	16'h	7cd9;
10942	:douta	=	16'h	8519;
10943	:douta	=	16'h	8d5b;
10944	:douta	=	16'h	8d7b;
10945	:douta	=	16'h	959c;
10946	:douta	=	16'h	8d5a;
10947	:douta	=	16'h	8d7b;
10948	:douta	=	16'h	959c;
10949	:douta	=	16'h	851a;
10950	:douta	=	16'h	7d1a;
10951	:douta	=	16'h	855b;
10952	:douta	=	16'h	95bc;
10953	:douta	=	16'h	8d7b;
10954	:douta	=	16'h	8d7b;
10955	:douta	=	16'h	855b;
10956	:douta	=	16'h	95bc;
10957	:douta	=	16'h	6c76;
10958	:douta	=	16'h	4b11;
10959	:douta	=	16'h	3b33;
10960	:douta	=	16'h	7d3b;
10961	:douta	=	16'h	857c;
10962	:douta	=	16'h	6458;
10963	:douta	=	16'h	6438;
10964	:douta	=	16'h	53d6;
10965	:douta	=	16'h	6478;
10966	:douta	=	16'h	6cd9;
10967	:douta	=	16'h	6cb9;
10968	:douta	=	16'h	74fa;
10969	:douta	=	16'h	7d7c;
10970	:douta	=	16'h	855b;
10971	:douta	=	16'h	8dbc;
10972	:douta	=	16'h	751a;
10973	:douta	=	16'h	74b9;
10974	:douta	=	16'h	6c99;
10975	:douta	=	16'h	74d9;
10976	:douta	=	16'h	7d3a;
10977	:douta	=	16'h	7d3b;
10978	:douta	=	16'h	7d1a;
10979	:douta	=	16'h	7d1a;
10980	:douta	=	16'h	855b;
10981	:douta	=	16'h	855b;
10982	:douta	=	16'h	7d1a;
10983	:douta	=	16'h	6cb9;
10984	:douta	=	16'h	95bc;
10985	:douta	=	16'h	74fa;
10986	:douta	=	16'h	6cba;
10987	:douta	=	16'h	6478;
10988	:douta	=	16'h	6c98;
10989	:douta	=	16'h	855b;
10990	:douta	=	16'h	6c97;
10991	:douta	=	16'h	6c77;
10992	:douta	=	16'h	4acf;
10993	:douta	=	16'h	1906;
10994	:douta	=	16'h	2189;
10995	:douta	=	16'h	7cb7;
10996	:douta	=	16'h	cebd;
10997	:douta	=	16'h	9d79;
10998	:douta	=	16'h	c65b;
10999	:douta	=	16'h	5bd4;
11000	:douta	=	16'h	3aaf;
11001	:douta	=	16'h	5330;
11002	:douta	=	16'h	63d2;
11003	:douta	=	16'h	ad77;
11004	:douta	=	16'h	a536;
11005	:douta	=	16'h	5b93;
11006	:douta	=	16'h	3ad0;
11007	:douta	=	16'h	4af0;
11008	:douta	=	16'h	4bb6;
11009	:douta	=	16'h	3b33;
11010	:douta	=	16'h	3b33;
11011	:douta	=	16'h	4333;
11012	:douta	=	16'h	5394;
11013	:douta	=	16'h	42d1;
11014	:douta	=	16'h	326f;
11015	:douta	=	16'h	322e;
11016	:douta	=	16'h	4311;
11017	:douta	=	16'h	63d3;
11018	:douta	=	16'h	5b93;
11019	:douta	=	16'h	84b7;
11020	:douta	=	16'h	8d39;
11021	:douta	=	16'h	6392;
11022	:douta	=	16'h	6bf3;
11023	:douta	=	16'h	7c35;
11024	:douta	=	16'h	5b70;
11025	:douta	=	16'h	9cd6;
11026	:douta	=	16'h	d659;
11027	:douta	=	16'h	d69b;
11028	:douta	=	16'h	b5f8;
11029	:douta	=	16'h	94b4;
11030	:douta	=	16'h	9472;
11031	:douta	=	16'h	bd95;
11032	:douta	=	16'h	8451;
11033	:douta	=	16'h	d657;
11034	:douta	=	16'h	d637;
11035	:douta	=	16'h	de97;
11036	:douta	=	16'h	ad34;
11037	:douta	=	16'h	b574;
11038	:douta	=	16'h	a512;
11039	:douta	=	16'h	5aed;
11040	:douta	=	16'h	83ae;
11041	:douta	=	16'h	7bcf;
11042	:douta	=	16'h	c5f4;
11043	:douta	=	16'h	bd94;
11044	:douta	=	16'h	c5d4;
11045	:douta	=	16'h	940f;
11046	:douta	=	16'h	acd1;
11047	:douta	=	16'h	8c4f;
11048	:douta	=	16'h	de56;
11049	:douta	=	16'h	62c9;
11050	:douta	=	16'h	c5b3;
11051	:douta	=	16'h	b530;
11052	:douta	=	16'h	ff9b;
11053	:douta	=	16'h	b592;
11054	:douta	=	16'h	a4b0;
11055	:douta	=	16'h	bd93;
11056	:douta	=	16'h	7bcd;
11057	:douta	=	16'h	7b2b;
11058	:douta	=	16'h	836b;
11059	:douta	=	16'h	8bcc;
11060	:douta	=	16'h	93ec;
11061	:douta	=	16'h	93cc;
11062	:douta	=	16'h	8bab;
11063	:douta	=	16'h	9c0d;
11064	:douta	=	16'h	9c0d;
11065	:douta	=	16'h	9c0d;
11066	:douta	=	16'h	9c0d;
11067	:douta	=	16'h	6aea;
11068	:douta	=	16'h	31a8;
11069	:douta	=	16'h	2125;
11070	:douta	=	16'h	2967;
11071	:douta	=	16'h	2987;
11072	:douta	=	16'h	2106;
11073	:douta	=	16'h	1905;
11074	:douta	=	16'h	39e9;
11075	:douta	=	16'h	1926;
11076	:douta	=	16'h	1105;
11077	:douta	=	16'h	18e5;
11078	:douta	=	16'h	18e5;
11079	:douta	=	16'h	18e5;
11080	:douta	=	16'h	18e5;
11081	:douta	=	16'h	1105;
11082	:douta	=	16'h	41e8;
11083	:douta	=	16'h	acd0;
11084	:douta	=	16'h	5aeb;
11085	:douta	=	16'h	0000;
11086	:douta	=	16'h	7c75;
11087	:douta	=	16'h	5b90;
11088	:douta	=	16'h	52cb;
11089	:douta	=	16'h	2147;
11090	:douta	=	16'h	636f;
11091	:douta	=	16'h	634d;
11092	:douta	=	16'h	52cc;
11093	:douta	=	16'h	3209;
11094	:douta	=	16'h	73cf;
11095	:douta	=	16'h	29a9;
11096	:douta	=	16'h	73d0;
11097	:douta	=	16'h	3a4c;
11098	:douta	=	16'h	4acc;
11099	:douta	=	16'h	1106;
11100	:douta	=	16'h	426a;
11101	:douta	=	16'h	5b2e;
11102	:douta	=	16'h	6b6f;
11103	:douta	=	16'h	29cb;
11104	:douta	=	16'h	6bd0;
11105	:douta	=	16'h	2a0c;
11106	:douta	=	16'h	6435;
11107	:douta	=	16'h	3b10;
11108	:douta	=	16'h	19ac;
11109	:douta	=	16'h	3acf;
11110	:douta	=	16'h	324d;
11111	:douta	=	16'h	42f1;
11112	:douta	=	16'h	5b91;
11113	:douta	=	16'h	5bf5;
11114	:douta	=	16'h	4b51;
11115	:douta	=	16'h	4acd;
11116	:douta	=	16'h	0800;
11117	:douta	=	16'h	0861;
11118	:douta	=	16'h	1061;
11119	:douta	=	16'h	0820;
11120	:douta	=	16'h	0000;
11121	:douta	=	16'h	31ea;
11122	:douta	=	16'h	4b31;
11123	:douta	=	16'h	3a8f;
11124	:douta	=	16'h	198a;
11125	:douta	=	16'h	5bf5;
11126	:douta	=	16'h	53f5;
11127	:douta	=	16'h	5c36;
11128	:douta	=	16'h	222e;
11129	:douta	=	16'h	524a;
11130	:douta	=	16'h	4a29;
11131	:douta	=	16'h	d550;
11132	:douta	=	16'h	734b;
11133	:douta	=	16'h	8d18;
11134	:douta	=	16'h	5bd5;
11135	:douta	=	16'h	5375;
11136	:douta	=	16'h	6c78;
11137	:douta	=	16'h	8d9b;
11138	:douta	=	16'h	84f9;
11139	:douta	=	16'h	853a;
11140	:douta	=	16'h	8519;
11141	:douta	=	16'h	8d7b;
11142	:douta	=	16'h	95bb;
11143	:douta	=	16'h	ae1c;
11144	:douta	=	16'h	957a;
11145	:douta	=	16'h	959b;
11146	:douta	=	16'h	7cd9;
11147	:douta	=	16'h	853a;
11148	:douta	=	16'h	8519;
11149	:douta	=	16'h	959b;
11150	:douta	=	16'h	a5fc;
11151	:douta	=	16'h	a5db;
11152	:douta	=	16'h	957a;
11153	:douta	=	16'h	7478;
11154	:douta	=	16'h	6c57;
11155	:douta	=	16'h	7cb8;
11156	:douta	=	16'h	8d5a;
11157	:douta	=	16'h	855a;
11158	:douta	=	16'h	8d5a;
11159	:douta	=	16'h	9dbb;
11160	:douta	=	16'h	8d5a;
11161	:douta	=	16'h	851a;
11162	:douta	=	16'h	8d39;
11163	:douta	=	16'h	7cd9;
11164	:douta	=	16'h	6c37;
11165	:douta	=	16'h	7cd8;
11166	:douta	=	16'h	9dbb;
11167	:douta	=	16'h	9ddb;
11168	:douta	=	16'h	8539;
11169	:douta	=	16'h	6c15;
11170	:douta	=	16'h	7497;
11171	:douta	=	16'h	957a;
11172	:douta	=	16'h	955a;
11173	:douta	=	16'h	6c16;
11174	:douta	=	16'h	7cb8;
11175	:douta	=	16'h	7cd8;
11176	:douta	=	16'h	95bb;
11177	:douta	=	16'h	8d5a;
11178	:douta	=	16'h	957b;
11179	:douta	=	16'h	74b8;
11180	:douta	=	16'h	855a;
11181	:douta	=	16'h	7cd9;
11182	:douta	=	16'h	7497;
11183	:douta	=	16'h	7cb8;
11184	:douta	=	16'h	7cf9;
11185	:douta	=	16'h	8d5b;
11186	:douta	=	16'h	7498;
11187	:douta	=	16'h	6c36;
11188	:douta	=	16'h	84f9;
11189	:douta	=	16'h	7cf9;
11190	:douta	=	16'h	84f9;
11191	:douta	=	16'h	8d5b;
11192	:douta	=	16'h	8d5b;
11193	:douta	=	16'h	853a;
11194	:douta	=	16'h	95bc;
11195	:douta	=	16'h	95bc;
11196	:douta	=	16'h	8d5b;
11197	:douta	=	16'h	853a;
11198	:douta	=	16'h	8d7b;
11199	:douta	=	16'h	959c;
11200	:douta	=	16'h	8d9b;
11201	:douta	=	16'h	8d5b;
11202	:douta	=	16'h	851a;
11203	:douta	=	16'h	959b;
11204	:douta	=	16'h	95bb;
11205	:douta	=	16'h	95bc;
11206	:douta	=	16'h	8d5b;
11207	:douta	=	16'h	8d7b;
11208	:douta	=	16'h	8d7b;
11209	:douta	=	16'h	853a;
11210	:douta	=	16'h	7cf9;
11211	:douta	=	16'h	857b;
11212	:douta	=	16'h	853a;
11213	:douta	=	16'h	851a;
11214	:douta	=	16'h	8d5b;
11215	:douta	=	16'h	95bd;
11216	:douta	=	16'h	853b;
11217	:douta	=	16'h	74d9;
11218	:douta	=	16'h	855b;
11219	:douta	=	16'h	857b;
11220	:douta	=	16'h	74fa;
11221	:douta	=	16'h	53f6;
11222	:douta	=	16'h	6458;
11223	:douta	=	16'h	751b;
11224	:douta	=	16'h	74fa;
11225	:douta	=	16'h	6498;
11226	:douta	=	16'h	6c99;
11227	:douta	=	16'h	751b;
11228	:douta	=	16'h	7d5b;
11229	:douta	=	16'h	859c;
11230	:douta	=	16'h	8ddc;
11231	:douta	=	16'h	6cb9;
11232	:douta	=	16'h	7d1a;
11233	:douta	=	16'h	6c79;
11234	:douta	=	16'h	74b9;
11235	:douta	=	16'h	7d5a;
11236	:douta	=	16'h	7d5b;
11237	:douta	=	16'h	859b;
11238	:douta	=	16'h	6cd9;
11239	:douta	=	16'h	8d7b;
11240	:douta	=	16'h	7d3a;
11241	:douta	=	16'h	74f9;
11242	:douta	=	16'h	7d5b;
11243	:douta	=	16'h	857b;
11244	:douta	=	16'h	7d5b;
11245	:douta	=	16'h	74da;
11246	:douta	=	16'h	74d9;
11247	:douta	=	16'h	74fa;
11248	:douta	=	16'h	74f9;
11249	:douta	=	16'h	6415;
11250	:douta	=	16'h	2127;
11251	:douta	=	16'h	2189;
11252	:douta	=	16'h	21ec;
11253	:douta	=	16'h	8cd5;
11254	:douta	=	16'h	7413;
11255	:douta	=	16'h	8cf5;
11256	:douta	=	16'h	73f3;
11257	:douta	=	16'h	6391;
11258	:douta	=	16'h	7c55;
11259	:douta	=	16'h	63b2;
11260	:douta	=	16'h	2a4f;
11261	:douta	=	16'h	5b91;
11262	:douta	=	16'h	63d3;
11263	:douta	=	16'h	8453;
11264	:douta	=	16'h	3b13;
11265	:douta	=	16'h	2ab1;
11266	:douta	=	16'h	2270;
11267	:douta	=	16'h	53d4;
11268	:douta	=	16'h	4332;
11269	:douta	=	16'h	7477;
11270	:douta	=	16'h	6416;
11271	:douta	=	16'h	6c36;
11272	:douta	=	16'h	6c77;
11273	:douta	=	16'h	3a8e;
11274	:douta	=	16'h	42cf;
11275	:douta	=	16'h	6bd4;
11276	:douta	=	16'h	7435;
11277	:douta	=	16'h	8475;
11278	:douta	=	16'h	9d17;
11279	:douta	=	16'h	8cb5;
11280	:douta	=	16'h	4b10;
11281	:douta	=	16'h	4aaf;
11282	:douta	=	16'h	be39;
11283	:douta	=	16'h	94b4;
11284	:douta	=	16'h	a576;
11285	:douta	=	16'h	ce17;
11286	:douta	=	16'h	c5d6;
11287	:douta	=	16'h	eeb8;
11288	:douta	=	16'h	8c52;
11289	:douta	=	16'h	ad34;
11290	:douta	=	16'h	b596;
11291	:douta	=	16'h	b596;
11292	:douta	=	16'h	9492;
11293	:douta	=	16'h	a4d2;
11294	:douta	=	16'h	bd94;
11295	:douta	=	16'h	8c10;
11296	:douta	=	16'h	eeb7;
11297	:douta	=	16'h	7bcf;
11298	:douta	=	16'h	9cd1;
11299	:douta	=	16'h	b574;
11300	:douta	=	16'h	83ef;
11301	:douta	=	16'h	83ce;
11302	:douta	=	16'h	de96;
11303	:douta	=	16'h	b512;
11304	:douta	=	16'h	eed7;
11305	:douta	=	16'h	738d;
11306	:douta	=	16'h	7b8d;
11307	:douta	=	16'h	948f;
11308	:douta	=	16'h	eef8;
11309	:douta	=	16'h	ad31;
11310	:douta	=	16'h	f737;
11311	:douta	=	16'h	f718;
11312	:douta	=	16'h	734a;
11313	:douta	=	16'h	836b;
11314	:douta	=	16'h	836b;
11315	:douta	=	16'h	93cc;
11316	:douta	=	16'h	940c;
11317	:douta	=	16'h	93ac;
11318	:douta	=	16'h	8bab;
11319	:douta	=	16'h	9c0c;
11320	:douta	=	16'h	ac6d;
11321	:douta	=	16'h	ac4d;
11322	:douta	=	16'h	a46d;
11323	:douta	=	16'h	9c0d;
11324	:douta	=	16'h	730b;
11325	:douta	=	16'h	5228;
11326	:douta	=	16'h	41e7;
11327	:douta	=	16'h	2946;
11328	:douta	=	16'h	1906;
11329	:douta	=	16'h	1905;
11330	:douta	=	16'h	2967;
11331	:douta	=	16'h	2968;
11332	:douta	=	16'h	1105;
11333	:douta	=	16'h	1906;
11334	:douta	=	16'h	1905;
11335	:douta	=	16'h	10e5;
11336	:douta	=	16'h	1905;
11337	:douta	=	16'h	1105;
11338	:douta	=	16'h	2125;
11339	:douta	=	16'h	840e;
11340	:douta	=	16'h	0001;
11341	:douta	=	16'h	0000;
11342	:douta	=	16'h	84d6;
11343	:douta	=	16'h	7c33;
11344	:douta	=	16'h	8470;
11345	:douta	=	16'h	7b8d;
11346	:douta	=	16'h	73ef;
11347	:douta	=	16'h	29a9;
11348	:douta	=	16'h	322a;
11349	:douta	=	16'h	2189;
11350	:douta	=	16'h	3209;
11351	:douta	=	16'h	1947;
11352	:douta	=	16'h	840f;
11353	:douta	=	16'h	21c9;
11354	:douta	=	16'h	73d0;
11355	:douta	=	16'h	3a0a;
11356	:douta	=	16'h	530d;
11357	:douta	=	16'h	3a2b;
11358	:douta	=	16'h	4acc;
11359	:douta	=	16'h	2148;
11360	:douta	=	16'h	5b4e;
11361	:douta	=	16'h	322c;
11362	:douta	=	16'h	7cd6;
11363	:douta	=	16'h	3b12;
11364	:douta	=	16'h	4b10;
11365	:douta	=	16'h	2a4f;
11366	:douta	=	16'h	32b0;
11367	:douta	=	16'h	21cc;
11368	:douta	=	16'h	42cf;
11369	:douta	=	16'h	3aaf;
11370	:douta	=	16'h	5393;
11371	:douta	=	16'h	4b94;
11372	:douta	=	16'h	39c8;
11373	:douta	=	16'h	18a2;
11374	:douta	=	16'h	1061;
11375	:douta	=	16'h	18a2;
11376	:douta	=	16'h	10a3;
11377	:douta	=	16'h	0000;
11378	:douta	=	16'h	18e4;
11379	:douta	=	16'h	7414;
11380	:douta	=	16'h	32af;
11381	:douta	=	16'h	2a4e;
11382	:douta	=	16'h	3ad1;
11383	:douta	=	16'h	5416;
11384	:douta	=	16'h	4374;
11385	:douta	=	16'h	5248;
11386	:douta	=	16'h	41a8;
11387	:douta	=	16'h	83cb;
11388	:douta	=	16'h	3967;
11389	:douta	=	16'h	a63e;
11390	:douta	=	16'h	8d7a;
11391	:douta	=	16'h	74b8;
11392	:douta	=	16'h	3af3;
11393	:douta	=	16'h	5bb5;
11394	:douta	=	16'h	8d7a;
11395	:douta	=	16'h	74b9;
11396	:douta	=	16'h	7cf9;
11397	:douta	=	16'h	7cd9;
11398	:douta	=	16'h	7d19;
11399	:douta	=	16'h	ae3c;
11400	:douta	=	16'h	ae3c;
11401	:douta	=	16'h	a61c;
11402	:douta	=	16'h	855a;
11403	:douta	=	16'h	95bb;
11404	:douta	=	16'h	7cd9;
11405	:douta	=	16'h	8d3a;
11406	:douta	=	16'h	8519;
11407	:douta	=	16'h	ae1c;
11408	:douta	=	16'h	a61c;
11409	:douta	=	16'h	9d9b;
11410	:douta	=	16'h	7c97;
11411	:douta	=	16'h	7c77;
11412	:douta	=	16'h	7457;
11413	:douta	=	16'h	8d5b;
11414	:douta	=	16'h	851a;
11415	:douta	=	16'h	8d3a;
11416	:douta	=	16'h	9ddc;
11417	:douta	=	16'h	8519;
11418	:douta	=	16'h	851a;
11419	:douta	=	16'h	851a;
11420	:douta	=	16'h	7cd8;
11421	:douta	=	16'h	7498;
11422	:douta	=	16'h	84f9;
11423	:douta	=	16'h	8d39;
11424	:douta	=	16'h	959a;
11425	:douta	=	16'h	8d39;
11426	:douta	=	16'h	6c36;
11427	:douta	=	16'h	7477;
11428	:douta	=	16'h	7cb8;
11429	:douta	=	16'h	955a;
11430	:douta	=	16'h	7477;
11431	:douta	=	16'h	6c15;
11432	:douta	=	16'h	7cb8;
11433	:douta	=	16'h	8d19;
11434	:douta	=	16'h	8d7b;
11435	:douta	=	16'h	8d5b;
11436	:douta	=	16'h	7cd9;
11437	:douta	=	16'h	84f9;
11438	:douta	=	16'h	7cb9;
11439	:douta	=	16'h	7cd8;
11440	:douta	=	16'h	7478;
11441	:douta	=	16'h	7cb9;
11442	:douta	=	16'h	853a;
11443	:douta	=	16'h	7cb8;
11444	:douta	=	16'h	7498;
11445	:douta	=	16'h	6416;
11446	:douta	=	16'h	8d5b;
11447	:douta	=	16'h	8d5b;
11448	:douta	=	16'h	959b;
11449	:douta	=	16'h	8519;
11450	:douta	=	16'h	7cd9;
11451	:douta	=	16'h	8d5a;
11452	:douta	=	16'h	9ddd;
11453	:douta	=	16'h	95bc;
11454	:douta	=	16'h	8d7b;
11455	:douta	=	16'h	853a;
11456	:douta	=	16'h	8d7b;
11457	:douta	=	16'h	9ddc;
11458	:douta	=	16'h	95bc;
11459	:douta	=	16'h	853a;
11460	:douta	=	16'h	855a;
11461	:douta	=	16'h	8d9b;
11462	:douta	=	16'h	855a;
11463	:douta	=	16'h	853a;
11464	:douta	=	16'h	855a;
11465	:douta	=	16'h	853a;
11466	:douta	=	16'h	853a;
11467	:douta	=	16'h	7d3a;
11468	:douta	=	16'h	7d1a;
11469	:douta	=	16'h	7d3a;
11470	:douta	=	16'h	7cfa;
11471	:douta	=	16'h	7d3b;
11472	:douta	=	16'h	95bc;
11473	:douta	=	16'h	9dfc;
11474	:douta	=	16'h	8d5b;
11475	:douta	=	16'h	853a;
11476	:douta	=	16'h	6c98;
11477	:douta	=	16'h	6458;
11478	:douta	=	16'h	53f6;
11479	:douta	=	16'h	6cb9;
11480	:douta	=	16'h	7d3b;
11481	:douta	=	16'h	751a;
11482	:douta	=	16'h	6c99;
11483	:douta	=	16'h	751b;
11484	:douta	=	16'h	74fb;
11485	:douta	=	16'h	74fa;
11486	:douta	=	16'h	8d9c;
11487	:douta	=	16'h	7d5b;
11488	:douta	=	16'h	7d3a;
11489	:douta	=	16'h	74b9;
11490	:douta	=	16'h	74b9;
11491	:douta	=	16'h	74da;
11492	:douta	=	16'h	7d3b;
11493	:douta	=	16'h	857c;
11494	:douta	=	16'h	74fa;
11495	:douta	=	16'h	7d1a;
11496	:douta	=	16'h	9dfd;
11497	:douta	=	16'h	751a;
11498	:douta	=	16'h	74da;
11499	:douta	=	16'h	6cda;
11500	:douta	=	16'h	751a;
11501	:douta	=	16'h	853b;
11502	:douta	=	16'h	7d1a;
11503	:douta	=	16'h	6c78;
11504	:douta	=	16'h	6cb8;
11505	:douta	=	16'h	7cfa;
11506	:douta	=	16'h	1906;
11507	:douta	=	16'h	2168;
11508	:douta	=	16'h	3aad;
11509	:douta	=	16'h	8c95;
11510	:douta	=	16'h	5b92;
11511	:douta	=	16'h	5371;
11512	:douta	=	16'h	3a8e;
11513	:douta	=	16'h	8494;
11514	:douta	=	16'h	7c54;
11515	:douta	=	16'h	c619;
11516	:douta	=	16'h	5373;
11517	:douta	=	16'h	326e;
11518	:douta	=	16'h	4b11;
11519	:douta	=	16'h	7c54;
11520	:douta	=	16'h	32f1;
11521	:douta	=	16'h	32f2;
11522	:douta	=	16'h	4bd5;
11523	:douta	=	16'h	4354;
11524	:douta	=	16'h	7cd9;
11525	:douta	=	16'h	4b52;
11526	:douta	=	16'h	6c57;
11527	:douta	=	16'h	5bb4;
11528	:douta	=	16'h	5bd4;
11529	:douta	=	16'h	5b72;
11530	:douta	=	16'h	6c35;
11531	:douta	=	16'h	84b7;
11532	:douta	=	16'h	8d18;
11533	:douta	=	16'h	5b31;
11534	:douta	=	16'h	8454;
11535	:douta	=	16'h	6bb2;
11536	:douta	=	16'h	6371;
11537	:douta	=	16'h	a537;
11538	:douta	=	16'h	ad36;
11539	:douta	=	16'h	c5d7;
11540	:douta	=	16'h	b597;
11541	:douta	=	16'h	8432;
11542	:douta	=	16'h	8c31;
11543	:douta	=	16'h	7c12;
11544	:douta	=	16'h	6370;
11545	:douta	=	16'h	8410;
11546	:douta	=	16'h	ce37;
11547	:douta	=	16'h	a534;
11548	:douta	=	16'h	b553;
11549	:douta	=	16'h	b553;
11550	:douta	=	16'h	b573;
11551	:douta	=	16'h	632d;
11552	:douta	=	16'h	942f;
11553	:douta	=	16'h	632d;
11554	:douta	=	16'h	9c90;
11555	:douta	=	16'h	942f;
11556	:douta	=	16'h	ce14;
11557	:douta	=	16'h	a4d0;
11558	:douta	=	16'h	de55;
11559	:douta	=	16'h	9490;
11560	:douta	=	16'h	83ee;
11561	:douta	=	16'h	942d;
11562	:douta	=	16'h	c592;
11563	:douta	=	16'h	acf0;
11564	:douta	=	16'h	ff5a;
11565	:douta	=	16'h	ce34;
11566	:douta	=	16'h	83cd;
11567	:douta	=	16'h	736b;
11568	:douta	=	16'h	838c;
11569	:douta	=	16'h	7b6b;
11570	:douta	=	16'h	838b;
11571	:douta	=	16'h	9c0c;
11572	:douta	=	16'h	9c0c;
11573	:douta	=	16'h	9c0c;
11574	:douta	=	16'h	9c0c;
11575	:douta	=	16'h	9c2d;
11576	:douta	=	16'h	b48d;
11577	:douta	=	16'h	b4ad;
11578	:douta	=	16'h	ac8e;
11579	:douta	=	16'h	836c;
11580	:douta	=	16'h	836b;
11581	:douta	=	16'h	838c;
11582	:douta	=	16'h	6b0a;
11583	:douta	=	16'h	5249;
11584	:douta	=	16'h	1105;
11585	:douta	=	16'h	1905;
11586	:douta	=	16'h	1906;
11587	:douta	=	16'h	1926;
11588	:douta	=	16'h	1905;
11589	:douta	=	16'h	1905;
11590	:douta	=	16'h	10e5;
11591	:douta	=	16'h	10e5;
11592	:douta	=	16'h	10e4;
11593	:douta	=	16'h	1905;
11594	:douta	=	16'h	10c3;
11595	:douta	=	16'h	10c3;
11596	:douta	=	16'h	0021;
11597	:douta	=	16'h	0000;
11598	:douta	=	16'h	6391;
11599	:douta	=	16'h	6c14;
11600	:douta	=	16'h	632e;
11601	:douta	=	16'h	4249;
11602	:douta	=	16'h	4a8b;
11603	:douta	=	16'h	5aeb;
11604	:douta	=	16'h	31c9;
11605	:douta	=	16'h	7bce;
11606	:douta	=	16'h	31eb;
11607	:douta	=	16'h	31ca;
11608	:douta	=	16'h	5b4f;
11609	:douta	=	16'h	29ea;
11610	:douta	=	16'h	3a4c;
11611	:douta	=	16'h	320a;
11612	:douta	=	16'h	73af;
11613	:douta	=	16'h	3a4a;
11614	:douta	=	16'h	5b0d;
11615	:douta	=	16'h	52cc;
11616	:douta	=	16'h	42ad;
11617	:douta	=	16'h	29aa;
11618	:douta	=	16'h	2a0b;
11619	:douta	=	16'h	322c;
11620	:douta	=	16'h	1949;
11621	:douta	=	16'h	73d1;
11622	:douta	=	16'h	6391;
11623	:douta	=	16'h	5351;
11624	:douta	=	16'h	5b91;
11625	:douta	=	16'h	326e;
11626	:douta	=	16'h	4b93;
11627	:douta	=	16'h	3ad1;
11628	:douta	=	16'h	3acf;
11629	:douta	=	16'h	328e;
11630	:douta	=	16'h	29c9;
11631	:douta	=	16'h	18c3;
11632	:douta	=	16'h	18c3;
11633	:douta	=	16'h	20e4;
11634	:douta	=	16'h	10e3;
11635	:douta	=	16'h	1061;
11636	:douta	=	16'h	3209;
11637	:douta	=	16'h	5350;
11638	:douta	=	16'h	32af;
11639	:douta	=	16'h	220c;
11640	:douta	=	16'h	3187;
11641	:douta	=	16'h	7289;
11642	:douta	=	16'h	cd70;
11643	:douta	=	16'h	5b0f;
11644	:douta	=	16'h	7d19;
11645	:douta	=	16'h	959a;
11646	:douta	=	16'h	8519;
11647	:douta	=	16'h	8d39;
11648	:douta	=	16'h	9d9a;
11649	:douta	=	16'h	8d7b;
11650	:douta	=	16'h	7477;
11651	:douta	=	16'h	851a;
11652	:douta	=	16'h	8d3a;
11653	:douta	=	16'h	53d6;
11654	:douta	=	16'h	6436;
11655	:douta	=	16'h	74d9;
11656	:douta	=	16'h	7cf9;
11657	:douta	=	16'h	ae1c;
11658	:douta	=	16'h	ae1b;
11659	:douta	=	16'h	95bb;
11660	:douta	=	16'h	95bb;
11661	:douta	=	16'h	959b;
11662	:douta	=	16'h	959b;
11663	:douta	=	16'h	8539;
11664	:douta	=	16'h	7477;
11665	:douta	=	16'h	7476;
11666	:douta	=	16'h	84f9;
11667	:douta	=	16'h	9d9a;
11668	:douta	=	16'h	9d7b;
11669	:douta	=	16'h	5311;
11670	:douta	=	16'h	957b;
11671	:douta	=	16'h	851a;
11672	:douta	=	16'h	84f9;
11673	:douta	=	16'h	8d7a;
11674	:douta	=	16'h	853a;
11675	:douta	=	16'h	8d5a;
11676	:douta	=	16'h	8d3a;
11677	:douta	=	16'h	84f9;
11678	:douta	=	16'h	957a;
11679	:douta	=	16'h	8d7a;
11680	:douta	=	16'h	7cb8;
11681	:douta	=	16'h	7497;
11682	:douta	=	16'h	84f9;
11683	:douta	=	16'h	8d3a;
11684	:douta	=	16'h	959b;
11685	:douta	=	16'h	84f9;
11686	:douta	=	16'h	63f5;
11687	:douta	=	16'h	63d4;
11688	:douta	=	16'h	8519;
11689	:douta	=	16'h	959a;
11690	:douta	=	16'h	7cd8;
11691	:douta	=	16'h	7cd8;
11692	:douta	=	16'h	959b;
11693	:douta	=	16'h	851a;
11694	:douta	=	16'h	7498;
11695	:douta	=	16'h	855a;
11696	:douta	=	16'h	7cf9;
11697	:douta	=	16'h	7cd8;
11698	:douta	=	16'h	7cd8;
11699	:douta	=	16'h	6c57;
11700	:douta	=	16'h	84d9;
11701	:douta	=	16'h	851a;
11702	:douta	=	16'h	8d3a;
11703	:douta	=	16'h	5bd5;
11704	:douta	=	16'h	6c16;
11705	:douta	=	16'h	851a;
11706	:douta	=	16'h	9ddc;
11707	:douta	=	16'h	959b;
11708	:douta	=	16'h	7cb9;
11709	:douta	=	16'h	7cf9;
11710	:douta	=	16'h	8d7b;
11711	:douta	=	16'h	8d7b;
11712	:douta	=	16'h	8d7c;
11713	:douta	=	16'h	7cd9;
11714	:douta	=	16'h	8519;
11715	:douta	=	16'h	95bc;
11716	:douta	=	16'h	959c;
11717	:douta	=	16'h	851a;
11718	:douta	=	16'h	8d5b;
11719	:douta	=	16'h	8d5a;
11720	:douta	=	16'h	8d7b;
11721	:douta	=	16'h	95dc;
11722	:douta	=	16'h	7d3a;
11723	:douta	=	16'h	8d7b;
11724	:douta	=	16'h	8d7b;
11725	:douta	=	16'h	853a;
11726	:douta	=	16'h	95bc;
11727	:douta	=	16'h	7cf9;
11728	:douta	=	16'h	853b;
11729	:douta	=	16'h	8d5b;
11730	:douta	=	16'h	8d7b;
11731	:douta	=	16'h	8d9b;
11732	:douta	=	16'h	9ddc;
11733	:douta	=	16'h	7d1a;
11734	:douta	=	16'h	751a;
11735	:douta	=	16'h	6498;
11736	:douta	=	16'h	4bd6;
11737	:douta	=	16'h	6cb9;
11738	:douta	=	16'h	855b;
11739	:douta	=	16'h	7d5b;
11740	:douta	=	16'h	6cda;
11741	:douta	=	16'h	6c99;
11742	:douta	=	16'h	6cda;
11743	:douta	=	16'h	6cd9;
11744	:douta	=	16'h	7d5c;
11745	:douta	=	16'h	859c;
11746	:douta	=	16'h	7d5b;
11747	:douta	=	16'h	7d5b;
11748	:douta	=	16'h	7d3b;
11749	:douta	=	16'h	6cda;
11750	:douta	=	16'h	6c99;
11751	:douta	=	16'h	74ba;
11752	:douta	=	16'h	751a;
11753	:douta	=	16'h	855b;
11754	:douta	=	16'h	753b;
11755	:douta	=	16'h	95dc;
11756	:douta	=	16'h	8dbc;
11757	:douta	=	16'h	5c17;
11758	:douta	=	16'h	7d3a;
11759	:douta	=	16'h	7d1a;
11760	:douta	=	16'h	7d1b;
11761	:douta	=	16'h	74f9;
11762	:douta	=	16'h	5b51;
11763	:douta	=	16'h	2988;
11764	:douta	=	16'h	2189;
11765	:douta	=	16'h	7c74;
11766	:douta	=	16'h	a536;
11767	:douta	=	16'h	6c35;
11768	:douta	=	16'h	94d6;
11769	:douta	=	16'h	4b11;
11770	:douta	=	16'h	5373;
11771	:douta	=	16'h	32b0;
11772	:douta	=	16'h	4b51;
11773	:douta	=	16'h	a598;
11774	:douta	=	16'h	9d58;
11775	:douta	=	16'h	5310;
11776	:douta	=	16'h	2ad1;
11777	:douta	=	16'h	224f;
11778	:douta	=	16'h	32d2;
11779	:douta	=	16'h	32f2;
11780	:douta	=	16'h	4311;
11781	:douta	=	16'h	4b52;
11782	:douta	=	16'h	7477;
11783	:douta	=	16'h	7477;
11784	:douta	=	16'h	7cd8;
11785	:douta	=	16'h	4b31;
11786	:douta	=	16'h	42f0;
11787	:douta	=	16'h	7c96;
11788	:douta	=	16'h	7435;
11789	:douta	=	16'h	7c33;
11790	:douta	=	16'h	a557;
11791	:douta	=	16'h	94d6;
11792	:douta	=	16'h	94b5;
11793	:douta	=	16'h	73f2;
11794	:douta	=	16'h	bdd8;
11795	:douta	=	16'h	8c93;
11796	:douta	=	16'h	a535;
11797	:douta	=	16'h	c5d5;
11798	:douta	=	16'h	cdf6;
11799	:douta	=	16'h	c5d6;
11800	:douta	=	16'h	94b2;
11801	:douta	=	16'h	8c52;
11802	:douta	=	16'h	bdb5;
11803	:douta	=	16'h	9cd2;
11804	:douta	=	16'h	9470;
11805	:douta	=	16'h	ad12;
11806	:douta	=	16'h	cdf5;
11807	:douta	=	16'h	52ab;
11808	:douta	=	16'h	ad12;
11809	:douta	=	16'h	a4b1;
11810	:douta	=	16'h	c5f4;
11811	:douta	=	16'h	ad11;
11812	:douta	=	16'h	7bad;
11813	:douta	=	16'h	7bad;
11814	:douta	=	16'h	f77a;
11815	:douta	=	16'h	630c;
11816	:douta	=	16'h	c594;
11817	:douta	=	16'h	62e9;
11818	:douta	=	16'h	8c2e;
11819	:douta	=	16'h	d614;
11820	:douta	=	16'h	bd72;
11821	:douta	=	16'h	c5f4;
11822	:douta	=	16'h	c613;
11823	:douta	=	16'h	838b;
11824	:douta	=	16'h	838b;
11825	:douta	=	16'h	836b;
11826	:douta	=	16'h	8b8b;
11827	:douta	=	16'h	9bec;
11828	:douta	=	16'h	9c0c;
11829	:douta	=	16'h	a42c;
11830	:douta	=	16'h	a44c;
11831	:douta	=	16'h	a46d;
11832	:douta	=	16'h	ac8d;
11833	:douta	=	16'h	b48d;
11834	:douta	=	16'h	ac8d;
11835	:douta	=	16'h	836c;
11836	:douta	=	16'h	836c;
11837	:douta	=	16'h	7b6b;
11838	:douta	=	16'h	6b2b;
11839	:douta	=	16'h	6aea;
11840	:douta	=	16'h	2167;
11841	:douta	=	16'h	1905;
11842	:douta	=	16'h	10c5;
11843	:douta	=	16'h	1105;
11844	:douta	=	16'h	2125;
11845	:douta	=	16'h	1905;
11846	:douta	=	16'h	10e5;
11847	:douta	=	16'h	10e5;
11848	:douta	=	16'h	10e5;
11849	:douta	=	16'h	1905;
11850	:douta	=	16'h	10c4;
11851	:douta	=	16'h	0021;
11852	:douta	=	16'h	0001;
11853	:douta	=	16'h	0000;
11854	:douta	=	16'h	5b2f;
11855	:douta	=	16'h	63f3;
11856	:douta	=	16'h	6bf2;
11857	:douta	=	16'h	7bac;
11858	:douta	=	16'h	4aab;
11859	:douta	=	16'h	528a;
11860	:douta	=	16'h	10c5;
11861	:douta	=	16'h	3a09;
11862	:douta	=	16'h	29a9;
11863	:douta	=	16'h	2168;
11864	:douta	=	16'h	52cd;
11865	:douta	=	16'h	29ca;
11866	:douta	=	16'h	530d;
11867	:douta	=	16'h	6b8e;
11868	:douta	=	16'h	5b4f;
11869	:douta	=	16'h	00a5;
11870	:douta	=	16'h	3a2a;
11871	:douta	=	16'h	29a8;
11872	:douta	=	16'h	3a4c;
11873	:douta	=	16'h	424b;
11874	:douta	=	16'h	42ef;
11875	:douta	=	16'h	324d;
11876	:douta	=	16'h	6370;
11877	:douta	=	16'h	3aaf;
11878	:douta	=	16'h	5372;
11879	:douta	=	16'h	324d;
11880	:douta	=	16'h	5351;
11881	:douta	=	16'h	3a4d;
11882	:douta	=	16'h	3ad0;
11883	:douta	=	16'h	2a6f;
11884	:douta	=	16'h	63f3;
11885	:douta	=	16'h	3acf;
11886	:douta	=	16'h	326d;
11887	:douta	=	16'h	2989;
11888	:douta	=	16'h	2124;
11889	:douta	=	16'h	18a3;
11890	:douta	=	16'h	1903;
11891	:douta	=	16'h	18e3;
11892	:douta	=	16'h	0841;
11893	:douta	=	16'h	2104;
11894	:douta	=	16'h	5b93;
11895	:douta	=	16'h	4b31;
11896	:douta	=	16'h	4a28;
11897	:douta	=	16'h	cd0f;
11898	:douta	=	16'h	7b8c;
11899	:douta	=	16'h	b63b;
11900	:douta	=	16'h	5c16;
11901	:douta	=	16'h	6416;
11902	:douta	=	16'h	8d79;
11903	:douta	=	16'h	8d5a;
11904	:douta	=	16'h	8d5a;
11905	:douta	=	16'h	9dbb;
11906	:douta	=	16'h	8519;
11907	:douta	=	16'h	7cf9;
11908	:douta	=	16'h	74b8;
11909	:douta	=	16'h	6c98;
11910	:douta	=	16'h	5bf6;
11911	:douta	=	16'h	6c77;
11912	:douta	=	16'h	6c57;
11913	:douta	=	16'h	74b8;
11914	:douta	=	16'h	ae3c;
11915	:douta	=	16'h	ae1c;
11916	:douta	=	16'h	9ddc;
11917	:douta	=	16'h	95bb;
11918	:douta	=	16'h	955a;
11919	:douta	=	16'h	a5db;
11920	:douta	=	16'h	9559;
11921	:douta	=	16'h	7cd7;
11922	:douta	=	16'h	6c16;
11923	:douta	=	16'h	6c56;
11924	:douta	=	16'h	8d3a;
11925	:douta	=	16'h	851a;
11926	:douta	=	16'h	8d5a;
11927	:douta	=	16'h	9dbb;
11928	:douta	=	16'h	ae1c;
11929	:douta	=	16'h	957b;
11930	:douta	=	16'h	8d5a;
11931	:douta	=	16'h	8539;
11932	:douta	=	16'h	8d5a;
11933	:douta	=	16'h	8d5a;
11934	:douta	=	16'h	8d5a;
11935	:douta	=	16'h	8d5a;
11936	:douta	=	16'h	8d39;
11937	:douta	=	16'h	7cf8;
11938	:douta	=	16'h	7cb8;
11939	:douta	=	16'h	6c36;
11940	:douta	=	16'h	7cb8;
11941	:douta	=	16'h	9d9b;
11942	:douta	=	16'h	84f8;
11943	:douta	=	16'h	6c35;
11944	:douta	=	16'h	7456;
11945	:douta	=	16'h	6c36;
11946	:douta	=	16'h	9dfc;
11947	:douta	=	16'h	95bb;
11948	:douta	=	16'h	957a;
11949	:douta	=	16'h	8d5a;
11950	:douta	=	16'h	8d7a;
11951	:douta	=	16'h	7cd9;
11952	:douta	=	16'h	7cb9;
11953	:douta	=	16'h	6c57;
11954	:douta	=	16'h	7cb8;
11955	:douta	=	16'h	7cb9;
11956	:douta	=	16'h	853a;
11957	:douta	=	16'h	7498;
11958	:douta	=	16'h	84f9;
11959	:douta	=	16'h	7cf9;
11960	:douta	=	16'h	7c98;
11961	:douta	=	16'h	6436;
11962	:douta	=	16'h	6416;
11963	:douta	=	16'h	957b;
11964	:douta	=	16'h	8d9c;
11965	:douta	=	16'h	8d7b;
11966	:douta	=	16'h	7d1a;
11967	:douta	=	16'h	851a;
11968	:douta	=	16'h	8d5b;
11969	:douta	=	16'h	8d5b;
11970	:douta	=	16'h	8d5a;
11971	:douta	=	16'h	7d1a;
11972	:douta	=	16'h	855b;
11973	:douta	=	16'h	8d7b;
11974	:douta	=	16'h	853a;
11975	:douta	=	16'h	7d1a;
11976	:douta	=	16'h	853a;
11977	:douta	=	16'h	855a;
11978	:douta	=	16'h	959b;
11979	:douta	=	16'h	853a;
11980	:douta	=	16'h	853b;
11981	:douta	=	16'h	855b;
11982	:douta	=	16'h	7d1a;
11983	:douta	=	16'h	8d9c;
11984	:douta	=	16'h	7cda;
11985	:douta	=	16'h	853a;
11986	:douta	=	16'h	855a;
11987	:douta	=	16'h	855a;
11988	:douta	=	16'h	8d7b;
11989	:douta	=	16'h	95bc;
11990	:douta	=	16'h	855a;
11991	:douta	=	16'h	7cf9;
11992	:douta	=	16'h	5c37;
11993	:douta	=	16'h	4374;
11994	:douta	=	16'h	74fa;
11995	:douta	=	16'h	751a;
11996	:douta	=	16'h	74f9;
11997	:douta	=	16'h	6cb9;
11998	:douta	=	16'h	6cba;
11999	:douta	=	16'h	5c38;
12000	:douta	=	16'h	6479;
12001	:douta	=	16'h	7d5c;
12002	:douta	=	16'h	85bc;
12003	:douta	=	16'h	74fa;
12004	:douta	=	16'h	857c;
12005	:douta	=	16'h	753b;
12006	:douta	=	16'h	7d1b;
12007	:douta	=	16'h	6cb9;
12008	:douta	=	16'h	7d5b;
12009	:douta	=	16'h	7d5c;
12010	:douta	=	16'h	7d3b;
12011	:douta	=	16'h	855b;
12012	:douta	=	16'h	8ddc;
12013	:douta	=	16'h	7cd9;
12014	:douta	=	16'h	6c78;
12015	:douta	=	16'h	74da;
12016	:douta	=	16'h	857b;
12017	:douta	=	16'h	859c;
12018	:douta	=	16'h	74b8;
12019	:douta	=	16'h	1906;
12020	:douta	=	16'h	2988;
12021	:douta	=	16'h	5372;
12022	:douta	=	16'h	4310;
12023	:douta	=	16'h	4b31;
12024	:douta	=	16'h	8cd6;
12025	:douta	=	16'h	a558;
12026	:douta	=	16'h	7cb8;
12027	:douta	=	16'h	5bb4;
12028	:douta	=	16'h	3290;
12029	:douta	=	16'h	63d3;
12030	:douta	=	16'h	7c33;
12031	:douta	=	16'h	7c75;
12032	:douta	=	16'h	4b94;
12033	:douta	=	16'h	3b54;
12034	:douta	=	16'h	3b32;
12035	:douta	=	16'h	4b95;
12036	:douta	=	16'h	3290;
12037	:douta	=	16'h	3ab0;
12038	:douta	=	16'h	3af1;
12039	:douta	=	16'h	2a2e;
12040	:douta	=	16'h	3ab0;
12041	:douta	=	16'h	7cb7;
12042	:douta	=	16'h	5351;
12043	:douta	=	16'h	7c76;
12044	:douta	=	16'h	9539;
12045	:douta	=	16'h	7414;
12046	:douta	=	16'h	7c33;
12047	:douta	=	16'h	8cb5;
12048	:douta	=	16'h	6c13;
12049	:douta	=	16'h	6bd3;
12050	:douta	=	16'h	9d15;
12051	:douta	=	16'h	9c93;
12052	:douta	=	16'h	c5f7;
12053	:douta	=	16'h	a4d4;
12054	:douta	=	16'h	9c92;
12055	:douta	=	16'h	39eb;
12056	:douta	=	16'h	6bb0;
12057	:douta	=	16'h	8451;
12058	:douta	=	16'h	a4b1;
12059	:douta	=	16'h	9470;
12060	:douta	=	16'h	cdf6;
12061	:douta	=	16'h	bd73;
12062	:douta	=	16'h	a4f2;
12063	:douta	=	16'h	9450;
12064	:douta	=	16'h	c5b3;
12065	:douta	=	16'h	5acb;
12066	:douta	=	16'h	a4b0;
12067	:douta	=	16'h	a4d0;
12068	:douta	=	16'h	e6b6;
12069	:douta	=	16'h	9c6f;
12070	:douta	=	16'h	de96;
12071	:douta	=	16'h	b572;
12072	:douta	=	16'h	ce14;
12073	:douta	=	16'h	83ad;
12074	:douta	=	16'h	b50f;
12075	:douta	=	16'h	ce34;
12076	:douta	=	16'h	eed7;
12077	:douta	=	16'h	a4f1;
12078	:douta	=	16'h	8bab;
12079	:douta	=	16'h	8bac;
12080	:douta	=	16'h	8bac;
12081	:douta	=	16'h	93cb;
12082	:douta	=	16'h	9c0c;
12083	:douta	=	16'h	9c0c;
12084	:douta	=	16'h	a40c;
12085	:douta	=	16'h	a44c;
12086	:douta	=	16'h	b48d;
12087	:douta	=	16'h	b4ad;
12088	:douta	=	16'h	ac6d;
12089	:douta	=	16'h	ac8d;
12090	:douta	=	16'h	b48e;
12091	:douta	=	16'h	ac6d;
12092	:douta	=	16'h	93cc;
12093	:douta	=	16'h	6aea;
12094	:douta	=	16'h	6aea;
12095	:douta	=	16'h	6b0a;
12096	:douta	=	16'h	524a;
12097	:douta	=	16'h	39c8;
12098	:douta	=	16'h	18e5;
12099	:douta	=	16'h	18e5;
12100	:douta	=	16'h	10e5;
12101	:douta	=	16'h	18e5;
12102	:douta	=	16'h	18e5;
12103	:douta	=	16'h	1905;
12104	:douta	=	16'h	1905;
12105	:douta	=	16'h	1905;
12106	:douta	=	16'h	1905;
12107	:douta	=	16'h	0883;
12108	:douta	=	16'h	0000;
12109	:douta	=	16'h	0002;
12110	:douta	=	16'h	3125;
12111	:douta	=	16'h	84b6;
12112	:douta	=	16'h	7cb6;
12113	:douta	=	16'h	3186;
12114	:douta	=	16'h	29a7;
12115	:douta	=	16'h	4229;
12116	:douta	=	16'h	10c5;
12117	:douta	=	16'h	630b;
12118	:douta	=	16'h	29a9;
12119	:douta	=	16'h	632d;
12120	:douta	=	16'h	42ac;
12121	:douta	=	16'h	422a;
12122	:douta	=	16'h	3a6b;
12123	:douta	=	16'h	428c;
12124	:douta	=	16'h	5b4e;
12125	:douta	=	16'h	5b0d;
12126	:douta	=	16'h	322b;
12127	:douta	=	16'h	6b6f;
12128	:douta	=	16'h	322b;
12129	:douta	=	16'h	2189;
12130	:douta	=	16'h	326d;
12131	:douta	=	16'h	1927;
12132	:douta	=	16'h	21cb;
12133	:douta	=	16'h	636f;
12134	:douta	=	16'h	21ca;
12135	:douta	=	16'h	6bd2;
12136	:douta	=	16'h	4b31;
12137	:douta	=	16'h	5372;
12138	:douta	=	16'h	4353;
12139	:douta	=	16'h	328f;
12140	:douta	=	16'h	326e;
12141	:douta	=	16'h	1969;
12142	:douta	=	16'h	320a;
12143	:douta	=	16'h	3a4b;
12144	:douta	=	16'h	5b50;
12145	:douta	=	16'h	532f;
12146	:douta	=	16'h	31a8;
12147	:douta	=	16'h	18c3;
12148	:douta	=	16'h	18e3;
12149	:douta	=	16'h	10c2;
12150	:douta	=	16'h	0840;
12151	:douta	=	16'h	0860;
12152	:douta	=	16'h	6a49;
12153	:douta	=	16'h	5269;
12154	:douta	=	16'h	73d2;
12155	:douta	=	16'h	9579;
12156	:douta	=	16'h	7498;
12157	:douta	=	16'h	959a;
12158	:douta	=	16'h	8d19;
12159	:douta	=	16'h	7cd7;
12160	:douta	=	16'h	84f9;
12161	:douta	=	16'h	7c98;
12162	:douta	=	16'h	7cb8;
12163	:douta	=	16'h	8d5a;
12164	:douta	=	16'h	8d5a;
12165	:douta	=	16'h	63d5;
12166	:douta	=	16'h	5394;
12167	:douta	=	16'h	84f9;
12168	:douta	=	16'h	7cb8;
12169	:douta	=	16'h	7cf8;
12170	:douta	=	16'h	5c16;
12171	:douta	=	16'h	7cd9;
12172	:douta	=	16'h	95bc;
12173	:douta	=	16'h	a5db;
12174	:douta	=	16'h	959a;
12175	:douta	=	16'h	8519;
12176	:douta	=	16'h	84d8;
12177	:douta	=	16'h	7c97;
12178	:douta	=	16'h	8d39;
12179	:douta	=	16'h	84b8;
12180	:douta	=	16'h	adfb;
12181	:douta	=	16'h	a5ba;
12182	:douta	=	16'h	6cb9;
12183	:douta	=	16'h	a5fc;
12184	:douta	=	16'h	9ddb;
12185	:douta	=	16'h	ae1c;
12186	:douta	=	16'h	b65c;
12187	:douta	=	16'h	957a;
12188	:douta	=	16'h	9dbb;
12189	:douta	=	16'h	957a;
12190	:douta	=	16'h	8519;
12191	:douta	=	16'h	84f9;
12192	:douta	=	16'h	8d5a;
12193	:douta	=	16'h	7cf9;
12194	:douta	=	16'h	851a;
12195	:douta	=	16'h	8d5a;
12196	:douta	=	16'h	8d39;
12197	:douta	=	16'h	7cd8;
12198	:douta	=	16'h	851a;
12199	:douta	=	16'h	8d3a;
12200	:douta	=	16'h	8d5a;
12201	:douta	=	16'h	95bb;
12202	:douta	=	16'h	7cb8;
12203	:douta	=	16'h	7477;
12204	:douta	=	16'h	7477;
12205	:douta	=	16'h	8d39;
12206	:douta	=	16'h	8d79;
12207	:douta	=	16'h	8d5a;
12208	:douta	=	16'h	853a;
12209	:douta	=	16'h	8519;
12210	:douta	=	16'h	7456;
12211	:douta	=	16'h	6c15;
12212	:douta	=	16'h	5bd5;
12213	:douta	=	16'h	6c57;
12214	:douta	=	16'h	7cd9;
12215	:douta	=	16'h	8d3a;
12216	:douta	=	16'h	7cd8;
12217	:douta	=	16'h	8d5a;
12218	:douta	=	16'h	9ddc;
12219	:douta	=	16'h	853a;
12220	:douta	=	16'h	6c36;
12221	:douta	=	16'h	6c16;
12222	:douta	=	16'h	7cf9;
12223	:douta	=	16'h	7cf9;
12224	:douta	=	16'h	851a;
12225	:douta	=	16'h	851a;
12226	:douta	=	16'h	853a;
12227	:douta	=	16'h	957b;
12228	:douta	=	16'h	959c;
12229	:douta	=	16'h	8d7b;
12230	:douta	=	16'h	853a;
12231	:douta	=	16'h	851a;
12232	:douta	=	16'h	8d9c;
12233	:douta	=	16'h	95bc;
12234	:douta	=	16'h	7d3a;
12235	:douta	=	16'h	7d3a;
12236	:douta	=	16'h	8d7b;
12237	:douta	=	16'h	8d7b;
12238	:douta	=	16'h	95dc;
12239	:douta	=	16'h	7d1b;
12240	:douta	=	16'h	853a;
12241	:douta	=	16'h	7cfa;
12242	:douta	=	16'h	853a;
12243	:douta	=	16'h	7d1a;
12244	:douta	=	16'h	8d7b;
12245	:douta	=	16'h	853a;
12246	:douta	=	16'h	855b;
12247	:douta	=	16'h	7cfa;
12248	:douta	=	16'h	8d9c;
12249	:douta	=	16'h	95dd;
12250	:douta	=	16'h	6c37;
12251	:douta	=	16'h	53b5;
12252	:douta	=	16'h	53b6;
12253	:douta	=	16'h	74da;
12254	:douta	=	16'h	74da;
12255	:douta	=	16'h	8dfd;
12256	:douta	=	16'h	7d5b;
12257	:douta	=	16'h	74fb;
12258	:douta	=	16'h	6cda;
12259	:douta	=	16'h	6cba;
12260	:douta	=	16'h	859c;
12261	:douta	=	16'h	7d5b;
12262	:douta	=	16'h	7d5b;
12263	:douta	=	16'h	859c;
12264	:douta	=	16'h	74fa;
12265	:douta	=	16'h	74fa;
12266	:douta	=	16'h	74d9;
12267	:douta	=	16'h	8dbc;
12268	:douta	=	16'h	857b;
12269	:douta	=	16'h	7d5b;
12270	:douta	=	16'h	857b;
12271	:douta	=	16'h	7d1a;
12272	:douta	=	16'h	855b;
12273	:douta	=	16'h	8d9c;
12274	:douta	=	16'h	6c77;
12275	:douta	=	16'h	5b72;
12276	:douta	=	16'h	18a4;
12277	:douta	=	16'h	326d;
12278	:douta	=	16'h	8cf6;
12279	:douta	=	16'h	8496;
12280	:douta	=	16'h	5b72;
12281	:douta	=	16'h	3aaf;
12282	:douta	=	16'h	42f1;
12283	:douta	=	16'h	6c13;
12284	:douta	=	16'h	9d37;
12285	:douta	=	16'h	6c14;
12286	:douta	=	16'h	8cd6;
12287	:douta	=	16'h	5331;
12288	:douta	=	16'h	4353;
12289	:douta	=	16'h	224f;
12290	:douta	=	16'h	220e;
12291	:douta	=	16'h	6479;
12292	:douta	=	16'h	4b73;
12293	:douta	=	16'h	5373;
12294	:douta	=	16'h	6c36;
12295	:douta	=	16'h	7497;
12296	:douta	=	16'h	5373;
12297	:douta	=	16'h	4b31;
12298	:douta	=	16'h	3a6e;
12299	:douta	=	16'h	5b72;
12300	:douta	=	16'h	5372;
12301	:douta	=	16'h	7414;
12302	:douta	=	16'h	8c74;
12303	:douta	=	16'h	a538;
12304	:douta	=	16'h	b5b9;
12305	:douta	=	16'h	7c34;
12306	:douta	=	16'h	9d35;
12307	:douta	=	16'h	3a4d;
12308	:douta	=	16'h	7413;
12309	:douta	=	16'h	c5d5;
12310	:douta	=	16'h	c5f6;
12311	:douta	=	16'h	bd55;
12312	:douta	=	16'h	bdd6;
12313	:douta	=	16'h	8c30;
12314	:douta	=	16'h	8431;
12315	:douta	=	16'h	428d;
12316	:douta	=	16'h	6b6e;
12317	:douta	=	16'h	83cf;
12318	:douta	=	16'h	bd74;
12319	:douta	=	16'h	b512;
12320	:douta	=	16'h	de76;
12321	:douta	=	16'h	944f;
12322	:douta	=	16'h	bdd3;
12323	:douta	=	16'h	842f;
12324	:douta	=	16'h	944e;
12325	:douta	=	16'h	acd0;
12326	:douta	=	16'h	e6d9;
12327	:douta	=	16'h	ce14;
12328	:douta	=	16'h	de96;
12329	:douta	=	16'h	5268;
12330	:douta	=	16'h	942d;
12331	:douta	=	16'h	ad11;
12332	:douta	=	16'h	ad10;
12333	:douta	=	16'h	9c8f;
12334	:douta	=	16'h	8bab;
12335	:douta	=	16'h	8bac;
12336	:douta	=	16'h	8bec;
12337	:douta	=	16'h	93ec;
12338	:douta	=	16'h	a42c;
12339	:douta	=	16'h	a44c;
12340	:douta	=	16'h	ac6d;
12341	:douta	=	16'h	ac6c;
12342	:douta	=	16'h	b4ad;
12343	:douta	=	16'h	bcce;
12344	:douta	=	16'h	a44c;
12345	:douta	=	16'h	ac4d;
12346	:douta	=	16'h	b48d;
12347	:douta	=	16'h	b4ae;
12348	:douta	=	16'h	9c0c;
12349	:douta	=	16'h	6aea;
12350	:douta	=	16'h	62ca;
12351	:douta	=	16'h	62a9;
12352	:douta	=	16'h	4a29;
12353	:douta	=	16'h	39e9;
12354	:douta	=	16'h	2167;
12355	:douta	=	16'h	10e5;
12356	:douta	=	16'h	1926;
12357	:douta	=	16'h	1905;
12358	:douta	=	16'h	18e5;
12359	:douta	=	16'h	1905;
12360	:douta	=	16'h	2106;
12361	:douta	=	16'h	1906;
12362	:douta	=	16'h	1925;
12363	:douta	=	16'h	1905;
12364	:douta	=	16'h	0000;
12365	:douta	=	16'h	0001;
12366	:douta	=	16'h	0000;
12367	:douta	=	16'h	7c95;
12368	:douta	=	16'h	63f2;
12369	:douta	=	16'h	638f;
12370	:douta	=	16'h	2187;
12371	:douta	=	16'h	630b;
12372	:douta	=	16'h	31a7;
12373	:douta	=	16'h	3208;
12374	:douta	=	16'h	18e5;
12375	:douta	=	16'h	31a7;
12376	:douta	=	16'h	322a;
12377	:douta	=	16'h	630e;
12378	:douta	=	16'h	322a;
12379	:douta	=	16'h	6bb0;
12380	:douta	=	16'h	2a2b;
12381	:douta	=	16'h	3a4b;
12382	:douta	=	16'h	2188;
12383	:douta	=	16'h	424b;
12384	:douta	=	16'h	4a8c;
12385	:douta	=	16'h	6b6e;
12386	:douta	=	16'h	2a4d;
12387	:douta	=	16'h	52ee;
12388	:douta	=	16'h	3a8d;
12389	:douta	=	16'h	2a2c;
12390	:douta	=	16'h	1989;
12391	:douta	=	16'h	5351;
12392	:douta	=	16'h	4b31;
12393	:douta	=	16'h	530f;
12394	:douta	=	16'h	3aaf;
12395	:douta	=	16'h	5b72;
12396	:douta	=	16'h	3b11;
12397	:douta	=	16'h	2a2c;
12398	:douta	=	16'h	3a6d;
12399	:douta	=	16'h	428c;
12400	:douta	=	16'h	5b50;
12401	:douta	=	16'h	324c;
12402	:douta	=	16'h	6bb2;
12403	:douta	=	16'h	10e3;
12404	:douta	=	16'h	1082;
12405	:douta	=	16'h	18c3;
12406	:douta	=	16'h	1062;
12407	:douta	=	16'h	2924;
12408	:douta	=	16'h	ac2c;
12409	:douta	=	16'h	528b;
12410	:douta	=	16'h	b5da;
12411	:douta	=	16'h	84d8;
12412	:douta	=	16'h	955a;
12413	:douta	=	16'h	8d19;
12414	:douta	=	16'h	84d8;
12415	:douta	=	16'h	8d3a;
12416	:douta	=	16'h	957a;
12417	:douta	=	16'h	8519;
12418	:douta	=	16'h	7cd8;
12419	:douta	=	16'h	6c57;
12420	:douta	=	16'h	7457;
12421	:douta	=	16'h	957a;
12422	:douta	=	16'h	6c77;
12423	:douta	=	16'h	6415;
12424	:douta	=	16'h	84d8;
12425	:douta	=	16'h	957a;
12426	:douta	=	16'h	6c77;
12427	:douta	=	16'h	6c36;
12428	:douta	=	16'h	84f9;
12429	:douta	=	16'h	957a;
12430	:douta	=	16'h	8d19;
12431	:douta	=	16'h	9d9a;
12432	:douta	=	16'h	9d9a;
12433	:douta	=	16'h	84b8;
12434	:douta	=	16'h	84f8;
12435	:douta	=	16'h	63f4;
12436	:douta	=	16'h	8d5a;
12437	:douta	=	16'h	ae1b;
12438	:douta	=	16'h	957b;
12439	:douta	=	16'h	b67d;
12440	:douta	=	16'h	ae3c;
12441	:douta	=	16'h	9dfb;
12442	:douta	=	16'h	a61c;
12443	:douta	=	16'h	8d7a;
12444	:douta	=	16'h	a61c;
12445	:douta	=	16'h	8d7a;
12446	:douta	=	16'h	9dfb;
12447	:douta	=	16'h	957b;
12448	:douta	=	16'h	8d3a;
12449	:douta	=	16'h	8d3a;
12450	:douta	=	16'h	8519;
12451	:douta	=	16'h	851a;
12452	:douta	=	16'h	959a;
12453	:douta	=	16'h	8d5a;
12454	:douta	=	16'h	7cf9;
12455	:douta	=	16'h	8d3a;
12456	:douta	=	16'h	8519;
12457	:douta	=	16'h	8519;
12458	:douta	=	16'h	84d9;
12459	:douta	=	16'h	8d3a;
12460	:douta	=	16'h	8d7a;
12461	:douta	=	16'h	7c97;
12462	:douta	=	16'h	7477;
12463	:douta	=	16'h	853a;
12464	:douta	=	16'h	7cf9;
12465	:douta	=	16'h	853a;
12466	:douta	=	16'h	95bc;
12467	:douta	=	16'h	7d19;
12468	:douta	=	16'h	7457;
12469	:douta	=	16'h	63f5;
12470	:douta	=	16'h	7cd9;
12471	:douta	=	16'h	8539;
12472	:douta	=	16'h	8519;
12473	:douta	=	16'h	6c36;
12474	:douta	=	16'h	74b8;
12475	:douta	=	16'h	8d7b;
12476	:douta	=	16'h	855a;
12477	:douta	=	16'h	84f9;
12478	:douta	=	16'h	7498;
12479	:douta	=	16'h	6456;
12480	:douta	=	16'h	7477;
12481	:douta	=	16'h	7cb8;
12482	:douta	=	16'h	95bc;
12483	:douta	=	16'h	74b8;
12484	:douta	=	16'h	7d1a;
12485	:douta	=	16'h	8d7b;
12486	:douta	=	16'h	8d7b;
12487	:douta	=	16'h	8d7b;
12488	:douta	=	16'h	853a;
12489	:douta	=	16'h	8d5b;
12490	:douta	=	16'h	95bc;
12491	:douta	=	16'h	7d1a;
12492	:douta	=	16'h	7cd9;
12493	:douta	=	16'h	8d5b;
12494	:douta	=	16'h	8d5b;
12495	:douta	=	16'h	95bc;
12496	:douta	=	16'h	8d7b;
12497	:douta	=	16'h	855b;
12498	:douta	=	16'h	74b8;
12499	:douta	=	16'h	7d1a;
12500	:douta	=	16'h	7d1a;
12501	:douta	=	16'h	855b;
12502	:douta	=	16'h	855b;
12503	:douta	=	16'h	851b;
12504	:douta	=	16'h	855b;
12505	:douta	=	16'h	8dbc;
12506	:douta	=	16'h	95dd;
12507	:douta	=	16'h	8dbc;
12508	:douta	=	16'h	5394;
12509	:douta	=	16'h	3ad1;
12510	:douta	=	16'h	53f6;
12511	:douta	=	16'h	7d7c;
12512	:douta	=	16'h	8ddd;
12513	:douta	=	16'h	857c;
12514	:douta	=	16'h	7d7c;
12515	:douta	=	16'h	5c78;
12516	:douta	=	16'h	859c;
12517	:douta	=	16'h	85bc;
12518	:douta	=	16'h	7d3b;
12519	:douta	=	16'h	751a;
12520	:douta	=	16'h	751a;
12521	:douta	=	16'h	751a;
12522	:douta	=	16'h	74fa;
12523	:douta	=	16'h	74d9;
12524	:douta	=	16'h	8dbc;
12525	:douta	=	16'h	853b;
12526	:douta	=	16'h	7d5b;
12527	:douta	=	16'h	859b;
12528	:douta	=	16'h	857b;
12529	:douta	=	16'h	7d3a;
12530	:douta	=	16'h	7d19;
12531	:douta	=	16'h	6416;
12532	:douta	=	16'h	31c9;
12533	:douta	=	16'h	29e9;
12534	:douta	=	16'h	5351;
12535	:douta	=	16'h	9d36;
12536	:douta	=	16'h	7c76;
12537	:douta	=	16'h	5bb3;
12538	:douta	=	16'h	7c55;
12539	:douta	=	16'h	326e;
12540	:douta	=	16'h	6c14;
12541	:douta	=	16'h	42cf;
12542	:douta	=	16'h	8cd6;
12543	:douta	=	16'h	adb8;
12544	:douta	=	16'h	3b33;
12545	:douta	=	16'h	4354;
12546	:douta	=	16'h	3b53;
12547	:douta	=	16'h	2a6f;
12548	:douta	=	16'h	5c16;
12549	:douta	=	16'h	4333;
12550	:douta	=	16'h	6c36;
12551	:douta	=	16'h	6c15;
12552	:douta	=	16'h	6c16;
12553	:douta	=	16'h	42f1;
12554	:douta	=	16'h	7415;
12555	:douta	=	16'h	73f4;
12556	:douta	=	16'h	9518;
12557	:douta	=	16'h	5330;
12558	:douta	=	16'h	7c33;
12559	:douta	=	16'h	8cb5;
12560	:douta	=	16'h	6bb2;
12561	:douta	=	16'h	6371;
12562	:douta	=	16'h	8411;
12563	:douta	=	16'h	ad56;
12564	:douta	=	16'h	bdd6;
12565	:douta	=	16'h	ad15;
12566	:douta	=	16'h	b555;
12567	:douta	=	16'h	a4f4;
12568	:douta	=	16'h	8c71;
12569	:douta	=	16'h	73af;
12570	:douta	=	16'h	9c91;
12571	:douta	=	16'h	ad13;
12572	:douta	=	16'h	9491;
12573	:douta	=	16'h	bd93;
12574	:douta	=	16'h	b574;
12575	:douta	=	16'h	a4b0;
12576	:douta	=	16'h	cdd3;
12577	:douta	=	16'h	5269;
12578	:douta	=	16'h	bdb3;
12579	:douta	=	16'h	8c6f;
12580	:douta	=	16'h	bd72;
12581	:douta	=	16'h	942e;
12582	:douta	=	16'h	ef1a;
12583	:douta	=	16'h	940e;
12584	:douta	=	16'h	bd92;
12585	:douta	=	16'h	940d;
12586	:douta	=	16'h	d614;
12587	:douta	=	16'h	c614;
12588	:douta	=	16'h	7b4b;
12589	:douta	=	16'h	838b;
12590	:douta	=	16'h	8bac;
12591	:douta	=	16'h	93cc;
12592	:douta	=	16'h	9c0c;
12593	:douta	=	16'h	9c0c;
12594	:douta	=	16'h	9c2b;
12595	:douta	=	16'h	ac6c;
12596	:douta	=	16'h	ac6c;
12597	:douta	=	16'h	b48d;
12598	:douta	=	16'h	bcce;
12599	:douta	=	16'h	bcce;
12600	:douta	=	16'h	b4cd;
12601	:douta	=	16'h	b46d;
12602	:douta	=	16'h	a42c;
12603	:douta	=	16'h	9c0c;
12604	:douta	=	16'h	9c0c;
12605	:douta	=	16'h	9c0d;
12606	:douta	=	16'h	838c;
12607	:douta	=	16'h	732b;
12608	:douta	=	16'h	524a;
12609	:douta	=	16'h	4a29;
12610	:douta	=	16'h	31a8;
12611	:douta	=	16'h	2987;
12612	:douta	=	16'h	4a29;
12613	:douta	=	16'h	0884;
12614	:douta	=	16'h	18e5;
12615	:douta	=	16'h	2126;
12616	:douta	=	16'h	1905;
12617	:douta	=	16'h	18e5;
12618	:douta	=	16'h	10e4;
12619	:douta	=	16'h	1105;
12620	:douta	=	16'h	0001;
12621	:douta	=	16'h	0000;
12622	:douta	=	16'h	0001;
12623	:douta	=	16'h	528c;
12624	:douta	=	16'h	6c12;
12625	:douta	=	16'h	530e;
12626	:douta	=	16'h	2147;
12627	:douta	=	16'h	2987;
12628	:douta	=	16'h	6b2c;
12629	:douta	=	16'h	7bef;
12630	:douta	=	16'h	1925;
12631	:douta	=	16'h	6b4c;
12632	:douta	=	16'h	42ac;
12633	:douta	=	16'h	426b;
12634	:douta	=	16'h	2188;
12635	:douta	=	16'h	3a8c;
12636	:douta	=	16'h	1106;
12637	:douta	=	16'h	5b2e;
12638	:douta	=	16'h	320b;
12639	:douta	=	16'h	5b0d;
12640	:douta	=	16'h	3a2b;
12641	:douta	=	16'h	4a8c;
12642	:douta	=	16'h	218a;
12643	:douta	=	16'h	29c9;
12644	:douta	=	16'h	2a0b;
12645	:douta	=	16'h	2a0b;
12646	:douta	=	16'h	2168;
12647	:douta	=	16'h	5b4f;
12648	:douta	=	16'h	530f;
12649	:douta	=	16'h	5bd3;
12650	:douta	=	16'h	4b30;
12651	:douta	=	16'h	5372;
12652	:douta	=	16'h	324e;
12653	:douta	=	16'h	428e;
12654	:douta	=	16'h	08a5;
12655	:douta	=	16'h	5b2f;
12656	:douta	=	16'h	530f;
12657	:douta	=	16'h	5b70;
12658	:douta	=	16'h	42f0;
12659	:douta	=	16'h	4b0f;
12660	:douta	=	16'h	42cf;
12661	:douta	=	16'h	29a8;
12662	:douta	=	16'h	18a2;
12663	:douta	=	16'h	3166;
12664	:douta	=	16'h	836b;
12665	:douta	=	16'h	9d39;
12666	:douta	=	16'h	7497;
12667	:douta	=	16'h	8d59;
12668	:douta	=	16'h	8539;
12669	:douta	=	16'h	8539;
12670	:douta	=	16'h	7477;
12671	:douta	=	16'h	7cb8;
12672	:douta	=	16'h	7cb8;
12673	:douta	=	16'h	7cb8;
12674	:douta	=	16'h	8519;
12675	:douta	=	16'h	957a;
12676	:douta	=	16'h	8d39;
12677	:douta	=	16'h	7477;
12678	:douta	=	16'h	8d19;
12679	:douta	=	16'h	8d5a;
12680	:douta	=	16'h	8538;
12681	:douta	=	16'h	6415;
12682	:douta	=	16'h	6c36;
12683	:douta	=	16'h	7cd8;
12684	:douta	=	16'h	95bb;
12685	:douta	=	16'h	7c77;
12686	:douta	=	16'h	7477;
12687	:douta	=	16'h	7cd8;
12688	:douta	=	16'h	8d59;
12689	:douta	=	16'h	8518;
12690	:douta	=	16'h	84b7;
12691	:douta	=	16'h	8cf8;
12692	:douta	=	16'h	7c97;
12693	:douta	=	16'h	8cf8;
12694	:douta	=	16'h	ae3c;
12695	:douta	=	16'h	9ddc;
12696	:douta	=	16'h	9dbb;
12697	:douta	=	16'h	b63d;
12698	:douta	=	16'h	95bb;
12699	:douta	=	16'h	959b;
12700	:douta	=	16'h	b65d;
12701	:douta	=	16'h	b65d;
12702	:douta	=	16'h	9dfc;
12703	:douta	=	16'h	9dbc;
12704	:douta	=	16'h	7cd8;
12705	:douta	=	16'h	8d7b;
12706	:douta	=	16'h	8519;
12707	:douta	=	16'h	8d3a;
12708	:douta	=	16'h	7cd9;
12709	:douta	=	16'h	7cd8;
12710	:douta	=	16'h	959b;
12711	:douta	=	16'h	853a;
12712	:douta	=	16'h	8519;
12713	:douta	=	16'h	84f9;
12714	:douta	=	16'h	8d5a;
12715	:douta	=	16'h	95bb;
12716	:douta	=	16'h	8d5a;
12717	:douta	=	16'h	84f9;
12718	:douta	=	16'h	8d3a;
12719	:douta	=	16'h	853a;
12720	:douta	=	16'h	8d5b;
12721	:douta	=	16'h	7497;
12722	:douta	=	16'h	63d5;
12723	:douta	=	16'h	7477;
12724	:douta	=	16'h	7cf9;
12725	:douta	=	16'h	8d5a;
12726	:douta	=	16'h	74b8;
12727	:douta	=	16'h	6c16;
12728	:douta	=	16'h	5bd4;
12729	:douta	=	16'h	84f9;
12730	:douta	=	16'h	851a;
12731	:douta	=	16'h	63f5;
12732	:douta	=	16'h	74b8;
12733	:douta	=	16'h	7cf9;
12734	:douta	=	16'h	7d19;
12735	:douta	=	16'h	8d5b;
12736	:douta	=	16'h	8d3a;
12737	:douta	=	16'h	7498;
12738	:douta	=	16'h	7498;
12739	:douta	=	16'h	6c57;
12740	:douta	=	16'h	6c78;
12741	:douta	=	16'h	7d1a;
12742	:douta	=	16'h	74b9;
12743	:douta	=	16'h	74d9;
12744	:douta	=	16'h	8d7b;
12745	:douta	=	16'h	8d9b;
12746	:douta	=	16'h	857b;
12747	:douta	=	16'h	74b8;
12748	:douta	=	16'h	7d19;
12749	:douta	=	16'h	8d7c;
12750	:douta	=	16'h	8d5b;
12751	:douta	=	16'h	74b9;
12752	:douta	=	16'h	853b;
12753	:douta	=	16'h	959c;
12754	:douta	=	16'h	853a;
12755	:douta	=	16'h	853a;
12756	:douta	=	16'h	8d5b;
12757	:douta	=	16'h	8d5b;
12758	:douta	=	16'h	7d1a;
12759	:douta	=	16'h	7d1a;
12760	:douta	=	16'h	851b;
12761	:douta	=	16'h	855a;
12762	:douta	=	16'h	853b;
12763	:douta	=	16'h	855b;
12764	:douta	=	16'h	7d5b;
12765	:douta	=	16'h	8ddd;
12766	:douta	=	16'h	855b;
12767	:douta	=	16'h	5bd5;
12768	:douta	=	16'h	6437;
12769	:douta	=	16'h	74fa;
12770	:douta	=	16'h	74fa;
12771	:douta	=	16'h	6cda;
12772	:douta	=	16'h	751b;
12773	:douta	=	16'h	6cda;
12774	:douta	=	16'h	7d5b;
12775	:douta	=	16'h	7d5b;
12776	:douta	=	16'h	74fa;
12777	:douta	=	16'h	857b;
12778	:douta	=	16'h	857b;
12779	:douta	=	16'h	7d5b;
12780	:douta	=	16'h	7d3a;
12781	:douta	=	16'h	7d3b;
12782	:douta	=	16'h	7d5b;
12783	:douta	=	16'h	7d3b;
12784	:douta	=	16'h	857c;
12785	:douta	=	16'h	855b;
12786	:douta	=	16'h	7d1a;
12787	:douta	=	16'h	7cd9;
12788	:douta	=	16'h	63d3;
12789	:douta	=	16'h	10c5;
12790	:douta	=	16'h	63b2;
12791	:douta	=	16'h	6bf4;
12792	:douta	=	16'h	63b2;
12793	:douta	=	16'h	7434;
12794	:douta	=	16'h	5351;
12795	:douta	=	16'h	9d78;
12796	:douta	=	16'h	63b2;
12797	:douta	=	16'h	a5b9;
12798	:douta	=	16'h	6c13;
12799	:douta	=	16'h	42d0;
12800	:douta	=	16'h	220d;
12801	:douta	=	16'h	3b12;
12802	:douta	=	16'h	2ab0;
12803	:douta	=	16'h	224f;
12804	:douta	=	16'h	6457;
12805	:douta	=	16'h	6416;
12806	:douta	=	16'h	7436;
12807	:douta	=	16'h	7456;
12808	:douta	=	16'h	6436;
12809	:douta	=	16'h	5b94;
12810	:douta	=	16'h	4b11;
12811	:douta	=	16'h	7435;
12812	:douta	=	16'h	8496;
12813	:douta	=	16'h	6bf3;
12814	:douta	=	16'h	9d37;
12815	:douta	=	16'h	adba;
12816	:douta	=	16'h	9d16;
12817	:douta	=	16'h	9d37;
12818	:douta	=	16'h	9493;
12819	:douta	=	16'h	4aef;
12820	:douta	=	16'h	6370;
12821	:douta	=	16'h	c617;
12822	:douta	=	16'h	bdb5;
12823	:douta	=	16'h	cdd6;
12824	:douta	=	16'h	b573;
12825	:douta	=	16'h	bd53;
12826	:douta	=	16'h	9c91;
12827	:douta	=	16'h	9cf2;
12828	:douta	=	16'h	7c10;
12829	:douta	=	16'h	632c;
12830	:douta	=	16'h	736d;
12831	:douta	=	16'h	bd72;
12832	:douta	=	16'h	f737;
12833	:douta	=	16'h	942e;
12834	:douta	=	16'h	9cb0;
12835	:douta	=	16'h	840e;
12836	:douta	=	16'h	83ee;
12837	:douta	=	16'h	8c0e;
12838	:douta	=	16'h	de56;
12839	:douta	=	16'h	d655;
12840	:douta	=	16'h	eef8;
12841	:douta	=	16'h	838c;
12842	:douta	=	16'h	8bed;
12843	:douta	=	16'h	ad32;
12844	:douta	=	16'h	838b;
12845	:douta	=	16'h	93cc;
12846	:douta	=	16'h	93cb;
12847	:douta	=	16'h	940c;
12848	:douta	=	16'h	a42c;
12849	:douta	=	16'h	9c0c;
12850	:douta	=	16'h	a42c;
12851	:douta	=	16'h	ac6c;
12852	:douta	=	16'h	b48c;
12853	:douta	=	16'h	bcee;
12854	:douta	=	16'h	bcee;
12855	:douta	=	16'h	bccd;
12856	:douta	=	16'h	c50e;
12857	:douta	=	16'h	bced;
12858	:douta	=	16'h	ac4d;
12859	:douta	=	16'h	9bec;
12860	:douta	=	16'h	8bab;
12861	:douta	=	16'h	8b6c;
12862	:douta	=	16'h	8b8d;
12863	:douta	=	16'h	838b;
12864	:douta	=	16'h	5a69;
12865	:douta	=	16'h	4a29;
12866	:douta	=	16'h	41e9;
12867	:douta	=	16'h	29a8;
12868	:douta	=	16'h	2946;
12869	:douta	=	16'h	10e4;
12870	:douta	=	16'h	18e5;
12871	:douta	=	16'h	2126;
12872	:douta	=	16'h	18e5;
12873	:douta	=	16'h	10e4;
12874	:douta	=	16'h	18e5;
12875	:douta	=	16'h	1104;
12876	:douta	=	16'h	10a4;
12877	:douta	=	16'h	0000;
12878	:douta	=	16'h	0022;
12879	:douta	=	16'h	2125;
12880	:douta	=	16'h	6370;
12881	:douta	=	16'h	63b1;
12882	:douta	=	16'h	426c;
12883	:douta	=	16'h	3a08;
12884	:douta	=	16'h	4269;
12885	:douta	=	16'h	31e8;
12886	:douta	=	16'h	10e4;
12887	:douta	=	16'h	39a8;
12888	:douta	=	16'h	2987;
12889	:douta	=	16'h	4aab;
12890	:douta	=	16'h	3a2a;
12891	:douta	=	16'h	42ce;
12892	:douta	=	16'h	1107;
12893	:douta	=	16'h	29ea;
12894	:douta	=	16'h	1968;
12895	:douta	=	16'h	4a8b;
12896	:douta	=	16'h	1126;
12897	:douta	=	16'h	5b0d;
12898	:douta	=	16'h	08e6;
12899	:douta	=	16'h	4aac;
12900	:douta	=	16'h	42ad;
12901	:douta	=	16'h	1169;
12902	:douta	=	16'h	1927;
12903	:douta	=	16'h	3a6d;
12904	:douta	=	16'h	322b;
12905	:douta	=	16'h	3a4c;
12906	:douta	=	16'h	6390;
12907	:douta	=	16'h	6bd2;
12908	:douta	=	16'h	42cf;
12909	:douta	=	16'h	3aae;
12910	:douta	=	16'h	2a0c;
12911	:douta	=	16'h	3aae;
12912	:douta	=	16'h	2a2c;
12913	:douta	=	16'h	3a8d;
12914	:douta	=	16'h	1128;
12915	:douta	=	16'h	6391;
12916	:douta	=	16'h	3a4c;
12917	:douta	=	16'h	73f2;
12918	:douta	=	16'h	39e8;
12919	:douta	=	16'h	6227;
12920	:douta	=	16'h	4a29;
12921	:douta	=	16'h	ae7c;
12922	:douta	=	16'h	7cd7;
12923	:douta	=	16'h	7cb7;
12924	:douta	=	16'h	7477;
12925	:douta	=	16'h	7456;
12926	:douta	=	16'h	8d5a;
12927	:douta	=	16'h	8d39;
12928	:douta	=	16'h	6c57;
12929	:douta	=	16'h	6415;
12930	:douta	=	16'h	74b8;
12931	:douta	=	16'h	7cd8;
12932	:douta	=	16'h	84d8;
12933	:douta	=	16'h	8d19;
12934	:douta	=	16'h	7477;
12935	:douta	=	16'h	8539;
12936	:douta	=	16'h	8d5a;
12937	:douta	=	16'h	959b;
12938	:douta	=	16'h	6c35;
12939	:douta	=	16'h	5bd5;
12940	:douta	=	16'h	7457;
12941	:douta	=	16'h	9559;
12942	:douta	=	16'h	8d19;
12943	:douta	=	16'h	6416;
12944	:douta	=	16'h	7c98;
12945	:douta	=	16'h	8d39;
12946	:douta	=	16'h	7c96;
12947	:douta	=	16'h	9559;
12948	:douta	=	16'h	9d7a;
12949	:douta	=	16'h	adfb;
12950	:douta	=	16'h	9d9a;
12951	:douta	=	16'h	b67d;
12952	:douta	=	16'h	ae3d;
12953	:douta	=	16'h	a5fc;
12954	:douta	=	16'h	ae3d;
12955	:douta	=	16'h	7d1a;
12956	:douta	=	16'h	9ddc;
12957	:douta	=	16'h	b67d;
12958	:douta	=	16'h	ae3d;
12959	:douta	=	16'h	a61c;
12960	:douta	=	16'h	959b;
12961	:douta	=	16'h	7cd9;
12962	:douta	=	16'h	95bb;
12963	:douta	=	16'h	8519;
12964	:douta	=	16'h	7cd8;
12965	:douta	=	16'h	957b;
12966	:douta	=	16'h	8d3a;
12967	:douta	=	16'h	853a;
12968	:douta	=	16'h	8d5a;
12969	:douta	=	16'h	957b;
12970	:douta	=	16'h	8519;
12971	:douta	=	16'h	8d5a;
12972	:douta	=	16'h	8d3a;
12973	:douta	=	16'h	853a;
12974	:douta	=	16'h	8519;
12975	:douta	=	16'h	8d3a;
12976	:douta	=	16'h	957b;
12977	:douta	=	16'h	7cd8;
12978	:douta	=	16'h	84f9;
12979	:douta	=	16'h	7457;
12980	:douta	=	16'h	5bf5;
12981	:douta	=	16'h	7477;
12982	:douta	=	16'h	6c56;
12983	:douta	=	16'h	853a;
12984	:douta	=	16'h	74b8;
12985	:douta	=	16'h	6c77;
12986	:douta	=	16'h	851a;
12987	:douta	=	16'h	6c37;
12988	:douta	=	16'h	74b8;
12989	:douta	=	16'h	84fa;
12990	:douta	=	16'h	7498;
12991	:douta	=	16'h	7cf9;
12992	:douta	=	16'h	851a;
12993	:douta	=	16'h	84f9;
12994	:douta	=	16'h	7cd9;
12995	:douta	=	16'h	74b8;
12996	:douta	=	16'h	6c57;
12997	:douta	=	16'h	6c98;
12998	:douta	=	16'h	6c57;
12999	:douta	=	16'h	6c77;
13000	:douta	=	16'h	7cfa;
13001	:douta	=	16'h	7d1a;
13002	:douta	=	16'h	8d5a;
13003	:douta	=	16'h	8d5a;
13004	:douta	=	16'h	7cf9;
13005	:douta	=	16'h	74d9;
13006	:douta	=	16'h	855b;
13007	:douta	=	16'h	853b;
13008	:douta	=	16'h	851a;
13009	:douta	=	16'h	855a;
13010	:douta	=	16'h	855b;
13011	:douta	=	16'h	8d9b;
13012	:douta	=	16'h	8d7b;
13013	:douta	=	16'h	853a;
13014	:douta	=	16'h	853b;
13015	:douta	=	16'h	7d1a;
13016	:douta	=	16'h	74b9;
13017	:douta	=	16'h	855b;
13018	:douta	=	16'h	7d3b;
13019	:douta	=	16'h	855b;
13020	:douta	=	16'h	7d1a;
13021	:douta	=	16'h	855b;
13022	:douta	=	16'h	7d3b;
13023	:douta	=	16'h	857c;
13024	:douta	=	16'h	7d3a;
13025	:douta	=	16'h	74da;
13026	:douta	=	16'h	6cba;
13027	:douta	=	16'h	7d1b;
13028	:douta	=	16'h	751a;
13029	:douta	=	16'h	6cd9;
13030	:douta	=	16'h	6cba;
13031	:douta	=	16'h	6cba;
13032	:douta	=	16'h	6c99;
13033	:douta	=	16'h	6cb9;
13034	:douta	=	16'h	7d3b;
13035	:douta	=	16'h	8ddc;
13036	:douta	=	16'h	74d9;
13037	:douta	=	16'h	751b;
13038	:douta	=	16'h	859c;
13039	:douta	=	16'h	8d9b;
13040	:douta	=	16'h	8dbc;
13041	:douta	=	16'h	8ddc;
13042	:douta	=	16'h	74f9;
13043	:douta	=	16'h	74d9;
13044	:douta	=	16'h	74d8;
13045	:douta	=	16'h	0884;
13046	:douta	=	16'h	4ace;
13047	:douta	=	16'h	42cf;
13048	:douta	=	16'h	add9;
13049	:douta	=	16'h	9d58;
13050	:douta	=	16'h	8495;
13051	:douta	=	16'h	5b92;
13052	:douta	=	16'h	7c54;
13053	:douta	=	16'h	6bd2;
13054	:douta	=	16'h	ad78;
13055	:douta	=	16'h	6371;
13056	:douta	=	16'h	2ab0;
13057	:douta	=	16'h	4b95;
13058	:douta	=	16'h	32f2;
13059	:douta	=	16'h	4312;
13060	:douta	=	16'h	5c36;
13061	:douta	=	16'h	4b74;
13062	:douta	=	16'h	7c76;
13063	:douta	=	16'h	7477;
13064	:douta	=	16'h	63f4;
13065	:douta	=	16'h	5352;
13066	:douta	=	16'h	7cb8;
13067	:douta	=	16'h	6bf3;
13068	:douta	=	16'h	84b7;
13069	:douta	=	16'h	5b92;
13070	:douta	=	16'h	7413;
13071	:douta	=	16'h	8cb5;
13072	:douta	=	16'h	7c13;
13073	:douta	=	16'h	6bd2;
13074	:douta	=	16'h	a514;
13075	:douta	=	16'h	b535;
13076	:douta	=	16'h	deb9;
13077	:douta	=	16'h	7c12;
13078	:douta	=	16'h	ad14;
13079	:douta	=	16'h	7b90;
13080	:douta	=	16'h	8451;
13081	:douta	=	16'h	4a6c;
13082	:douta	=	16'h	a4d1;
13083	:douta	=	16'h	a4f2;
13084	:douta	=	16'h	9cd1;
13085	:douta	=	16'h	b552;
13086	:douta	=	16'h	e696;
13087	:douta	=	16'h	944f;
13088	:douta	=	16'h	9c6f;
13089	:douta	=	16'h	7bac;
13090	:douta	=	16'h	ce34;
13091	:douta	=	16'h	bd92;
13092	:douta	=	16'h	7c0d;
13093	:douta	=	16'h	7b4c;
13094	:douta	=	16'h	e6b7;
13095	:douta	=	16'h	b531;
13096	:douta	=	16'h	bdb2;
13097	:douta	=	16'h	accf;
13098	:douta	=	16'h	b571;
13099	:douta	=	16'h	7309;
13100	:douta	=	16'h	93ec;
13101	:douta	=	16'h	9c0d;
13102	:douta	=	16'h	9c0c;
13103	:douta	=	16'h	9c0d;
13104	:douta	=	16'h	ac4d;
13105	:douta	=	16'h	ac4c;
13106	:douta	=	16'h	b48d;
13107	:douta	=	16'h	b4cd;
13108	:douta	=	16'h	bced;
13109	:douta	=	16'h	cd4e;
13110	:douta	=	16'h	cd4f;
13111	:douta	=	16'h	d570;
13112	:douta	=	16'h	cd4f;
13113	:douta	=	16'h	cd6f;
13114	:douta	=	16'h	c50f;
13115	:douta	=	16'h	ac4d;
13116	:douta	=	16'h	9c0d;
13117	:douta	=	16'h	8b8c;
13118	:douta	=	16'h	72ca;
13119	:douta	=	16'h	5a68;
13120	:douta	=	16'h	62ca;
13121	:douta	=	16'h	5a6a;
13122	:douta	=	16'h	31c8;
13123	:douta	=	16'h	2967;
13124	:douta	=	16'h	2146;
13125	:douta	=	16'h	528a;
13126	:douta	=	16'h	630c;
13127	:douta	=	16'h	08a4;
13128	:douta	=	16'h	18e4;
13129	:douta	=	16'h	10e5;
13130	:douta	=	16'h	10e4;
13131	:douta	=	16'h	10e4;
13132	:douta	=	16'h	1905;
13133	:douta	=	16'h	1926;
13134	:douta	=	16'h	0000;
13135	:douta	=	16'h	0000;
13136	:douta	=	16'h	0020;
13137	:douta	=	16'h	6391;
13138	:douta	=	16'h	6bf1;
13139	:douta	=	16'h	428b;
13140	:douta	=	16'h	732b;
13141	:douta	=	16'h	52cb;
13142	:douta	=	16'h	940e;
13143	:douta	=	16'h	6b4d;
13144	:douta	=	16'h	2966;
13145	:douta	=	16'h	3a2a;
13146	:douta	=	16'h	29a9;
13147	:douta	=	16'h	29ea;
13148	:douta	=	16'h	422b;
13149	:douta	=	16'h	29a8;
13150	:douta	=	16'h	320a;
13151	:douta	=	16'h	73ae;
13152	:douta	=	16'h	632e;
13153	:douta	=	16'h	4aee;
13154	:douta	=	16'h	424b;
13155	:douta	=	16'h	42ce;
13156	:douta	=	16'h	1968;
13157	:douta	=	16'h	08a5;
13158	:douta	=	16'h	1106;
13159	:douta	=	16'h	29c9;
13160	:douta	=	16'h	4a8c;
13161	:douta	=	16'h	2189;
13162	:douta	=	16'h	4aee;
13163	:douta	=	16'h	32ae;
13164	:douta	=	16'h	3a4d;
13165	:douta	=	16'h	3a6d;
13166	:douta	=	16'h	21ca;
13167	:douta	=	16'h	3a4c;
13168	:douta	=	16'h	322c;
13169	:douta	=	16'h	3aaf;
13170	:douta	=	16'h	4ad0;
13171	:douta	=	16'h	5371;
13172	:douta	=	16'h	428d;
13173	:douta	=	16'h	4aaf;
13174	:douta	=	16'h	49a7;
13175	:douta	=	16'h	b48d;
13176	:douta	=	16'h	9cb5;
13177	:douta	=	16'h	84f9;
13178	:douta	=	16'h	7c97;
13179	:douta	=	16'h	84d8;
13180	:douta	=	16'h	84d8;
13181	:douta	=	16'h	955a;
13182	:douta	=	16'h	7497;
13183	:douta	=	16'h	7477;
13184	:douta	=	16'h	7cb7;
13185	:douta	=	16'h	84d8;
13186	:douta	=	16'h	84b7;
13187	:douta	=	16'h	7477;
13188	:douta	=	16'h	8d19;
13189	:douta	=	16'h	955a;
13190	:douta	=	16'h	8519;
13191	:douta	=	16'h	8cf8;
13192	:douta	=	16'h	8519;
13193	:douta	=	16'h	84d8;
13194	:douta	=	16'h	8519;
13195	:douta	=	16'h	8d3a;
13196	:douta	=	16'h	84d8;
13197	:douta	=	16'h	6415;
13198	:douta	=	16'h	6c57;
13199	:douta	=	16'h	7cb7;
13200	:douta	=	16'h	8d19;
13201	:douta	=	16'h	8d39;
13202	:douta	=	16'h	955a;
13203	:douta	=	16'h	84f8;
13204	:douta	=	16'h	b61b;
13205	:douta	=	16'h	ae1b;
13206	:douta	=	16'h	7cd8;
13207	:douta	=	16'h	957b;
13208	:douta	=	16'h	7498;
13209	:douta	=	16'h	9dfb;
13210	:douta	=	16'h	9dbc;
13211	:douta	=	16'h	7d19;
13212	:douta	=	16'h	8d5a;
13213	:douta	=	16'h	84f9;
13214	:douta	=	16'h	8d5a;
13215	:douta	=	16'h	95db;
13216	:douta	=	16'h	959b;
13217	:douta	=	16'h	9ddb;
13218	:douta	=	16'h	7498;
13219	:douta	=	16'h	7cd9;
13220	:douta	=	16'h	957b;
13221	:douta	=	16'h	8d7a;
13222	:douta	=	16'h	9ddc;
13223	:douta	=	16'h	8d7a;
13224	:douta	=	16'h	7cd9;
13225	:douta	=	16'h	8519;
13226	:douta	=	16'h	8d5a;
13227	:douta	=	16'h	8d39;
13228	:douta	=	16'h	8d3a;
13229	:douta	=	16'h	957b;
13230	:douta	=	16'h	8d7a;
13231	:douta	=	16'h	8d5a;
13232	:douta	=	16'h	853a;
13233	:douta	=	16'h	74b8;
13234	:douta	=	16'h	6c57;
13235	:douta	=	16'h	853a;
13236	:douta	=	16'h	851a;
13237	:douta	=	16'h	7cd9;
13238	:douta	=	16'h	8519;
13239	:douta	=	16'h	7477;
13240	:douta	=	16'h	6c16;
13241	:douta	=	16'h	7498;
13242	:douta	=	16'h	7498;
13243	:douta	=	16'h	8d3a;
13244	:douta	=	16'h	853a;
13245	:douta	=	16'h	851a;
13246	:douta	=	16'h	7cd9;
13247	:douta	=	16'h	851a;
13248	:douta	=	16'h	5bf6;
13249	:douta	=	16'h	7498;
13250	:douta	=	16'h	853a;
13251	:douta	=	16'h	74b8;
13252	:douta	=	16'h	851a;
13253	:douta	=	16'h	7cfa;
13254	:douta	=	16'h	7498;
13255	:douta	=	16'h	6c77;
13256	:douta	=	16'h	6c57;
13257	:douta	=	16'h	6c77;
13258	:douta	=	16'h	6437;
13259	:douta	=	16'h	6436;
13260	:douta	=	16'h	6436;
13261	:douta	=	16'h	95dc;
13262	:douta	=	16'h	95bc;
13263	:douta	=	16'h	855b;
13264	:douta	=	16'h	7cb9;
13265	:douta	=	16'h	7cf9;
13266	:douta	=	16'h	857b;
13267	:douta	=	16'h	7d1a;
13268	:douta	=	16'h	7d3a;
13269	:douta	=	16'h	8d5b;
13270	:douta	=	16'h	95bc;
13271	:douta	=	16'h	95dc;
13272	:douta	=	16'h	853b;
13273	:douta	=	16'h	855c;
13274	:douta	=	16'h	7d1b;
13275	:douta	=	16'h	7cfa;
13276	:douta	=	16'h	7d1b;
13277	:douta	=	16'h	853b;
13278	:douta	=	16'h	7d1b;
13279	:douta	=	16'h	857c;
13280	:douta	=	16'h	7d3a;
13281	:douta	=	16'h	74f9;
13282	:douta	=	16'h	74f9;
13283	:douta	=	16'h	8d9c;
13284	:douta	=	16'h	6c99;
13285	:douta	=	16'h	6479;
13286	:douta	=	16'h	751a;
13287	:douta	=	16'h	7d3b;
13288	:douta	=	16'h	74fa;
13289	:douta	=	16'h	6cb9;
13290	:douta	=	16'h	7d5b;
13291	:douta	=	16'h	7d5a;
13292	:douta	=	16'h	7d5a;
13293	:douta	=	16'h	95dc;
13294	:douta	=	16'h	6cb8;
13295	:douta	=	16'h	7cf9;
13296	:douta	=	16'h	7d5b;
13297	:douta	=	16'h	7d5b;
13298	:douta	=	16'h	855b;
13299	:douta	=	16'h	7d3a;
13300	:douta	=	16'h	7cf9;
13301	:douta	=	16'h	2167;
13302	:douta	=	16'h	1928;
13303	:douta	=	16'h	b5d9;
13304	:douta	=	16'h	2a0c;
13305	:douta	=	16'h	5b72;
13306	:douta	=	16'h	5b71;
13307	:douta	=	16'h	8474;
13308	:douta	=	16'h	7c33;
13309	:douta	=	16'h	9cf5;
13310	:douta	=	16'h	3a4c;
13311	:douta	=	16'h	73b0;
13312	:douta	=	16'h	2a6f;
13313	:douta	=	16'h	2a2f;
13314	:douta	=	16'h	19ee;
13315	:douta	=	16'h	32f1;
13316	:douta	=	16'h	4b74;
13317	:douta	=	16'h	4b74;
13318	:douta	=	16'h	7c96;
13319	:douta	=	16'h	7cb8;
13320	:douta	=	16'h	6c16;
13321	:douta	=	16'h	5372;
13322	:douta	=	16'h	5bb3;
13323	:douta	=	16'h	5310;
13324	:douta	=	16'h	6c14;
13325	:douta	=	16'h	5331;
13326	:douta	=	16'h	8433;
13327	:douta	=	16'h	9d16;
13328	:douta	=	16'h	9cd6;
13329	:douta	=	16'h	9d16;
13330	:douta	=	16'h	a4f3;
13331	:douta	=	16'h	ad75;
13332	:douta	=	16'h	b555;
13333	:douta	=	16'h	9493;
13334	:douta	=	16'h	bd75;
13335	:douta	=	16'h	ad33;
13336	:douta	=	16'h	ce35;
13337	:douta	=	16'h	a4b2;
13338	:douta	=	16'h	ad13;
13339	:douta	=	16'h	8c70;
13340	:douta	=	16'h	8c50;
13341	:douta	=	16'h	630c;
13342	:douta	=	16'h	8c30;
13343	:douta	=	16'h	a4b0;
13344	:douta	=	16'h	c5d4;
13345	:douta	=	16'h	cdf4;
13346	:douta	=	16'h	de56;
13347	:douta	=	16'h	ad11;
13348	:douta	=	16'h	9c8f;
13349	:douta	=	16'h	62ca;
13350	:douta	=	16'h	d655;
13351	:douta	=	16'h	d635;
13352	:douta	=	16'h	d676;
13353	:douta	=	16'h	948e;
13354	:douta	=	16'h	732a;
13355	:douta	=	16'h	7b4b;
13356	:douta	=	16'h	9bec;
13357	:douta	=	16'h	9c2d;
13358	:douta	=	16'h	a44d;
13359	:douta	=	16'h	9c0c;
13360	:douta	=	16'h	a44c;
13361	:douta	=	16'h	b4ad;
13362	:douta	=	16'h	bcce;
13363	:douta	=	16'h	bcee;
13364	:douta	=	16'h	c50e;
13365	:douta	=	16'h	cd4e;
13366	:douta	=	16'h	d590;
13367	:douta	=	16'h	d590;
13368	:douta	=	16'h	cd70;
13369	:douta	=	16'h	d571;
13370	:douta	=	16'h	d591;
13371	:douta	=	16'h	bcee;
13372	:douta	=	16'h	ac6d;
13373	:douta	=	16'h	9c0d;
13374	:douta	=	16'h	93ed;
13375	:douta	=	16'h	6aa9;
13376	:douta	=	16'h	5a69;
13377	:douta	=	16'h	5228;
13378	:douta	=	16'h	526b;
13379	:douta	=	16'h	39c8;
13380	:douta	=	16'h	2987;
13381	:douta	=	16'h	29a8;
13382	:douta	=	16'h	5aaa;
13383	:douta	=	16'h	2125;
13384	:douta	=	16'h	10a4;
13385	:douta	=	16'h	18e5;
13386	:douta	=	16'h	10e4;
13387	:douta	=	16'h	18e5;
13388	:douta	=	16'h	18e5;
13389	:douta	=	16'h	1925;
13390	:douta	=	16'h	0000;
13391	:douta	=	16'h	0001;
13392	:douta	=	16'h	0000;
13393	:douta	=	16'h	52cd;
13394	:douta	=	16'h	7412;
13395	:douta	=	16'h	4a8c;
13396	:douta	=	16'h	52a9;
13397	:douta	=	16'h	4a69;
13398	:douta	=	16'h	5aaa;
13399	:douta	=	16'h	8c2e;
13400	:douta	=	16'h	734d;
13401	:douta	=	16'h	424b;
13402	:douta	=	16'h	4a8b;
13403	:douta	=	16'h	3a4c;
13404	:douta	=	16'h	424b;
13405	:douta	=	16'h	21a9;
13406	:douta	=	16'h	31ea;
13407	:douta	=	16'h	320a;
13408	:douta	=	16'h	73cf;
13409	:douta	=	16'h	42ad;
13410	:douta	=	16'h	6b4e;
13411	:douta	=	16'h	73b0;
13412	:douta	=	16'h	3a2b;
13413	:douta	=	16'h	29a9;
13414	:douta	=	16'h	29ca;
13415	:douta	=	16'h	1148;
13416	:douta	=	16'h	2168;
13417	:douta	=	16'h	0023;
13418	:douta	=	16'h	532f;
13419	:douta	=	16'h	21aa;
13420	:douta	=	16'h	3a2b;
13421	:douta	=	16'h	322c;
13422	:douta	=	16'h	326d;
13423	:douta	=	16'h	19aa;
13424	:douta	=	16'h	1969;
13425	:douta	=	16'h	21eb;
13426	:douta	=	16'h	0908;
13427	:douta	=	16'h	4b2f;
13428	:douta	=	16'h	630d;
13429	:douta	=	16'h	73d1;
13430	:douta	=	16'h	9b8d;
13431	:douta	=	16'h	9c0c;
13432	:douta	=	16'h	b63c;
13433	:douta	=	16'h	957a;
13434	:douta	=	16'h	a5db;
13435	:douta	=	16'h	8d39;
13436	:douta	=	16'h	7cb8;
13437	:douta	=	16'h	84f8;
13438	:douta	=	16'h	959a;
13439	:douta	=	16'h	9559;
13440	:douta	=	16'h	6c37;
13441	:douta	=	16'h	5bf5;
13442	:douta	=	16'h	7497;
13443	:douta	=	16'h	84d8;
13444	:douta	=	16'h	7c97;
13445	:douta	=	16'h	9dbb;
13446	:douta	=	16'h	9dba;
13447	:douta	=	16'h	7cb8;
13448	:douta	=	16'h	7cf8;
13449	:douta	=	16'h	8d5a;
13450	:douta	=	16'h	957a;
13451	:douta	=	16'h	955a;
13452	:douta	=	16'h	8d3a;
13453	:douta	=	16'h	84d8;
13454	:douta	=	16'h	6c57;
13455	:douta	=	16'h	7456;
13456	:douta	=	16'h	7497;
13457	:douta	=	16'h	84f9;
13458	:douta	=	16'h	84f9;
13459	:douta	=	16'h	8d19;
13460	:douta	=	16'h	be7c;
13461	:douta	=	16'h	b63b;
13462	:douta	=	16'h	84f9;
13463	:douta	=	16'h	9dbb;
13464	:douta	=	16'h	9d9a;
13465	:douta	=	16'h	7498;
13466	:douta	=	16'h	959a;
13467	:douta	=	16'h	8d7b;
13468	:douta	=	16'h	7cb8;
13469	:douta	=	16'h	8d3a;
13470	:douta	=	16'h	853a;
13471	:douta	=	16'h	851a;
13472	:douta	=	16'h	855a;
13473	:douta	=	16'h	8d5a;
13474	:douta	=	16'h	7d19;
13475	:douta	=	16'h	6c57;
13476	:douta	=	16'h	6c98;
13477	:douta	=	16'h	8d5b;
13478	:douta	=	16'h	8d7b;
13479	:douta	=	16'h	959b;
13480	:douta	=	16'h	8539;
13481	:douta	=	16'h	853a;
13482	:douta	=	16'h	84f9;
13483	:douta	=	16'h	84f9;
13484	:douta	=	16'h	7cd8;
13485	:douta	=	16'h	8539;
13486	:douta	=	16'h	853a;
13487	:douta	=	16'h	8d7b;
13488	:douta	=	16'h	959b;
13489	:douta	=	16'h	851a;
13490	:douta	=	16'h	63f5;
13491	:douta	=	16'h	5b94;
13492	:douta	=	16'h	7cb8;
13493	:douta	=	16'h	853a;
13494	:douta	=	16'h	7477;
13495	:douta	=	16'h	84f9;
13496	:douta	=	16'h	84f9;
13497	:douta	=	16'h	6c57;
13498	:douta	=	16'h	6457;
13499	:douta	=	16'h	7cf9;
13500	:douta	=	16'h	7cf9;
13501	:douta	=	16'h	8d5b;
13502	:douta	=	16'h	7498;
13503	:douta	=	16'h	7cd9;
13504	:douta	=	16'h	853a;
13505	:douta	=	16'h	7cd9;
13506	:douta	=	16'h	6c57;
13507	:douta	=	16'h	7cd9;
13508	:douta	=	16'h	7cd9;
13509	:douta	=	16'h	7cd9;
13510	:douta	=	16'h	7cfa;
13511	:douta	=	16'h	7d1a;
13512	:douta	=	16'h	6436;
13513	:douta	=	16'h	6c77;
13514	:douta	=	16'h	7498;
13515	:douta	=	16'h	6c57;
13516	:douta	=	16'h	6416;
13517	:douta	=	16'h	7498;
13518	:douta	=	16'h	7498;
13519	:douta	=	16'h	857b;
13520	:douta	=	16'h	8d9b;
13521	:douta	=	16'h	8dbb;
13522	:douta	=	16'h	7cd9;
13523	:douta	=	16'h	7cfa;
13524	:douta	=	16'h	7d3a;
13525	:douta	=	16'h	7d1a;
13526	:douta	=	16'h	7d3a;
13527	:douta	=	16'h	8d9c;
13528	:douta	=	16'h	95dd;
13529	:douta	=	16'h	8d9c;
13530	:douta	=	16'h	857c;
13531	:douta	=	16'h	7cfa;
13532	:douta	=	16'h	7d1a;
13533	:douta	=	16'h	7cfa;
13534	:douta	=	16'h	7d3b;
13535	:douta	=	16'h	855b;
13536	:douta	=	16'h	8dbc;
13537	:douta	=	16'h	7d1a;
13538	:douta	=	16'h	74fa;
13539	:douta	=	16'h	857b;
13540	:douta	=	16'h	857c;
13541	:douta	=	16'h	7d1a;
13542	:douta	=	16'h	6458;
13543	:douta	=	16'h	6478;
13544	:douta	=	16'h	7d3b;
13545	:douta	=	16'h	6458;
13546	:douta	=	16'h	6cd9;
13547	:douta	=	16'h	8dbc;
13548	:douta	=	16'h	857b;
13549	:douta	=	16'h	859b;
13550	:douta	=	16'h	857b;
13551	:douta	=	16'h	7d1b;
13552	:douta	=	16'h	74d9;
13553	:douta	=	16'h	7d1a;
13554	:douta	=	16'h	7d3b;
13555	:douta	=	16'h	7d3a;
13556	:douta	=	16'h	74d9;
13557	:douta	=	16'h	4aef;
13558	:douta	=	16'h	08a4;
13559	:douta	=	16'h	7c54;
13560	:douta	=	16'h	9cf6;
13561	:douta	=	16'h	7434;
13562	:douta	=	16'h	8cd6;
13563	:douta	=	16'h	6bd3;
13564	:douta	=	16'h	6bd3;
13565	:douta	=	16'h	636f;
13566	:douta	=	16'h	8433;
13567	:douta	=	16'h	a4f4;
13568	:douta	=	16'h	2a2f;
13569	:douta	=	16'h	4394;
13570	:douta	=	16'h	4374;
13571	:douta	=	16'h	2a8f;
13572	:douta	=	16'h	53d4;
13573	:douta	=	16'h	5c36;
13574	:douta	=	16'h	3ab0;
13575	:douta	=	16'h	7497;
13576	:douta	=	16'h	42d0;
13577	:douta	=	16'h	5b93;
13578	:douta	=	16'h	5372;
13579	:douta	=	16'h	7414;
13580	:douta	=	16'h	63b3;
13581	:douta	=	16'h	8cd7;
13582	:douta	=	16'h	8cd6;
13583	:douta	=	16'h	9537;
13584	:douta	=	16'h	9cf5;
13585	:douta	=	16'h	9d36;
13586	:douta	=	16'h	7bf1;
13587	:douta	=	16'h	9492;
13588	:douta	=	16'h	9cb3;
13589	:douta	=	16'h	9cf3;
13590	:douta	=	16'h	c5d5;
13591	:douta	=	16'h	a4d2;
13592	:douta	=	16'h	ad33;
13593	:douta	=	16'h	4aad;
13594	:douta	=	16'h	9cb1;
13595	:douta	=	16'h	9c90;
13596	:douta	=	16'h	c5d3;
13597	:douta	=	16'h	bd72;
13598	:douta	=	16'h	bd93;
13599	:douta	=	16'h	c5b3;
13600	:douta	=	16'h	de76;
13601	:douta	=	16'h	bd72;
13602	:douta	=	16'h	9cae;
13603	:douta	=	16'h	b552;
13604	:douta	=	16'h	a4d0;
13605	:douta	=	16'h	83cd;
13606	:douta	=	16'h	eed8;
13607	:douta	=	16'h	cdf3;
13608	:douta	=	16'h	ad32;
13609	:douta	=	16'h	7b0a;
13610	:douta	=	16'h	834b;
13611	:douta	=	16'h	838b;
13612	:douta	=	16'h	8bcb;
13613	:douta	=	16'h	93cc;
13614	:douta	=	16'h	ac6d;
13615	:douta	=	16'h	ac6c;
13616	:douta	=	16'h	b4ad;
13617	:douta	=	16'h	bd0e;
13618	:douta	=	16'h	cd4f;
13619	:douta	=	16'h	cd6f;
13620	:douta	=	16'h	d570;
13621	:douta	=	16'h	ddd2;
13622	:douta	=	16'h	ddd1;
13623	:douta	=	16'h	ddd1;
13624	:douta	=	16'h	ddd2;
13625	:douta	=	16'h	d5b1;
13626	:douta	=	16'h	ddd1;
13627	:douta	=	16'h	ddf3;
13628	:douta	=	16'h	ddf2;
13629	:douta	=	16'h	c50e;
13630	:douta	=	16'h	b48e;
13631	:douta	=	16'h	940d;
13632	:douta	=	16'h	5b0d;
13633	:douta	=	16'h	4a2a;
13634	:douta	=	16'h	5aab;
13635	:douta	=	16'h	52ab;
13636	:douta	=	16'h	2988;
13637	:douta	=	16'h	62cb;
13638	:douta	=	16'h	5acb;
13639	:douta	=	16'h	2967;
13640	:douta	=	16'h	31a8;
13641	:douta	=	16'h	10e5;
13642	:douta	=	16'h	18e5;
13643	:douta	=	16'h	1905;
13644	:douta	=	16'h	1904;
13645	:douta	=	16'h	1904;
13646	:douta	=	16'h	2145;
13647	:douta	=	16'h	0000;
13648	:douta	=	16'h	0000;
13649	:douta	=	16'h	0000;
13650	:douta	=	16'h	1906;
13651	:douta	=	16'h	6370;
13652	:douta	=	16'h	6370;
13653	:douta	=	16'h	2987;
13654	:douta	=	16'h	8c0d;
13655	:douta	=	16'h	6b0b;
13656	:douta	=	16'h	2105;
13657	:douta	=	16'h	18e4;
13658	:douta	=	16'h	2146;
13659	:douta	=	16'h	10e5;
13660	:douta	=	16'h	2127;
13661	:douta	=	16'h	1106;
13662	:douta	=	16'h	424b;
13663	:douta	=	16'h	4a8d;
13664	:douta	=	16'h	5b4e;
13665	:douta	=	16'h	2a0c;
13666	:douta	=	16'h	4acd;
13667	:douta	=	16'h	118a;
13668	:douta	=	16'h	428d;
13669	:douta	=	16'h	2188;
13670	:douta	=	16'h	532e;
13671	:douta	=	16'h	4a8a;
13672	:douta	=	16'h	3a4b;
13673	:douta	=	16'h	6baf;
13674	:douta	=	16'h	21eb;
13675	:douta	=	16'h	1947;
13676	:douta	=	16'h	3a6c;
13677	:douta	=	16'h	29a9;
13678	:douta	=	16'h	2189;
13679	:douta	=	16'h	320b;
13680	:douta	=	16'h	428d;
13681	:douta	=	16'h	0927;
13682	:douta	=	16'h	29ea;
13683	:douta	=	16'h	2a0c;
13684	:douta	=	16'h	5b50;
13685	:douta	=	16'h	326d;
13686	:douta	=	16'h	a42c;
13687	:douta	=	16'h	5acb;
13688	:douta	=	16'h	959a;
13689	:douta	=	16'h	84d8;
13690	:douta	=	16'h	84f9;
13691	:douta	=	16'h	7cd8;
13692	:douta	=	16'h	7cf8;
13693	:douta	=	16'h	8d39;
13694	:douta	=	16'h	8519;
13695	:douta	=	16'h	74b8;
13696	:douta	=	16'h	7cd8;
13697	:douta	=	16'h	957a;
13698	:douta	=	16'h	8d39;
13699	:douta	=	16'h	7477;
13700	:douta	=	16'h	7457;
13701	:douta	=	16'h	6c36;
13702	:douta	=	16'h	84f9;
13703	:douta	=	16'h	8518;
13704	:douta	=	16'h	84f9;
13705	:douta	=	16'h	84d9;
13706	:douta	=	16'h	74b8;
13707	:douta	=	16'h	7cb8;
13708	:douta	=	16'h	9ddb;
13709	:douta	=	16'h	a5db;
13710	:douta	=	16'h	9dbb;
13711	:douta	=	16'h	6416;
13712	:douta	=	16'h	8519;
13713	:douta	=	16'h	8d39;
13714	:douta	=	16'h	a5db;
13715	:douta	=	16'h	a5fc;
13716	:douta	=	16'h	9d9b;
13717	:douta	=	16'h	a5fb;
13718	:douta	=	16'h	957b;
13719	:douta	=	16'h	8d3a;
13720	:douta	=	16'h	8d5a;
13721	:douta	=	16'h	9dbc;
13722	:douta	=	16'h	853a;
13723	:douta	=	16'h	851a;
13724	:douta	=	16'h	8519;
13725	:douta	=	16'h	a61d;
13726	:douta	=	16'h	7cf9;
13727	:douta	=	16'h	7cf9;
13728	:douta	=	16'h	7d1a;
13729	:douta	=	16'h	6c97;
13730	:douta	=	16'h	6456;
13731	:douta	=	16'h	a5fb;
13732	:douta	=	16'h	b65d;
13733	:douta	=	16'h	851a;
13734	:douta	=	16'h	8d59;
13735	:douta	=	16'h	8519;
13736	:douta	=	16'h	853a;
13737	:douta	=	16'h	7cd9;
13738	:douta	=	16'h	8519;
13739	:douta	=	16'h	9ddc;
13740	:douta	=	16'h	8d39;
13741	:douta	=	16'h	7cd9;
13742	:douta	=	16'h	8d5a;
13743	:douta	=	16'h	8519;
13744	:douta	=	16'h	7477;
13745	:douta	=	16'h	7cf9;
13746	:douta	=	16'h	8d9b;
13747	:douta	=	16'h	855a;
13748	:douta	=	16'h	853a;
13749	:douta	=	16'h	7498;
13750	:douta	=	16'h	7457;
13751	:douta	=	16'h	851a;
13752	:douta	=	16'h	7cd9;
13753	:douta	=	16'h	6c57;
13754	:douta	=	16'h	7498;
13755	:douta	=	16'h	6c77;
13756	:douta	=	16'h	7cf9;
13757	:douta	=	16'h	7478;
13758	:douta	=	16'h	6c57;
13759	:douta	=	16'h	6456;
13760	:douta	=	16'h	8d5b;
13761	:douta	=	16'h	6416;
13762	:douta	=	16'h	7cd9;
13763	:douta	=	16'h	6c77;
13764	:douta	=	16'h	6415;
13765	:douta	=	16'h	6c36;
13766	:douta	=	16'h	7498;
13767	:douta	=	16'h	6416;
13768	:douta	=	16'h	5bb4;
13769	:douta	=	16'h	7477;
13770	:douta	=	16'h	6c77;
13771	:douta	=	16'h	7498;
13772	:douta	=	16'h	6c56;
13773	:douta	=	16'h	6c36;
13774	:douta	=	16'h	7cf9;
13775	:douta	=	16'h	6c77;
13776	:douta	=	16'h	74d9;
13777	:douta	=	16'h	6c98;
13778	:douta	=	16'h	8dbc;
13779	:douta	=	16'h	8d9c;
13780	:douta	=	16'h	855b;
13781	:douta	=	16'h	7d3b;
13782	:douta	=	16'h	7d1b;
13783	:douta	=	16'h	853b;
13784	:douta	=	16'h	7cfb;
13785	:douta	=	16'h	7d1b;
13786	:douta	=	16'h	8d7c;
13787	:douta	=	16'h	8dbc;
13788	:douta	=	16'h	7d1b;
13789	:douta	=	16'h	853b;
13790	:douta	=	16'h	6c99;
13791	:douta	=	16'h	8d7c;
13792	:douta	=	16'h	8d9d;
13793	:douta	=	16'h	7d3a;
13794	:douta	=	16'h	7d3a;
13795	:douta	=	16'h	7d3a;
13796	:douta	=	16'h	6c98;
13797	:douta	=	16'h	74b9;
13798	:douta	=	16'h	857b;
13799	:douta	=	16'h	857b;
13800	:douta	=	16'h	855b;
13801	:douta	=	16'h	74da;
13802	:douta	=	16'h	6cb9;
13803	:douta	=	16'h	6458;
13804	:douta	=	16'h	74da;
13805	:douta	=	16'h	857b;
13806	:douta	=	16'h	7d3a;
13807	:douta	=	16'h	857b;
13808	:douta	=	16'h	857b;
13809	:douta	=	16'h	8d9c;
13810	:douta	=	16'h	7d3a;
13811	:douta	=	16'h	74fa;
13812	:douta	=	16'h	7cfa;
13813	:douta	=	16'h	6c77;
13814	:douta	=	16'h	2169;
13815	:douta	=	16'h	7c75;
13816	:douta	=	16'h	5351;
13817	:douta	=	16'h	7433;
13818	:douta	=	16'h	4b0f;
13819	:douta	=	16'h	7413;
13820	:douta	=	16'h	ad57;
13821	:douta	=	16'h	94b4;
13822	:douta	=	16'h	8453;
13823	:douta	=	16'h	3a4c;
13824	:douta	=	16'h	3312;
13825	:douta	=	16'h	4395;
13826	:douta	=	16'h	4b95;
13827	:douta	=	16'h	220d;
13828	:douta	=	16'h	4b73;
13829	:douta	=	16'h	3b12;
13830	:douta	=	16'h	5bb3;
13831	:douta	=	16'h	7477;
13832	:douta	=	16'h	63f4;
13833	:douta	=	16'h	5b93;
13834	:douta	=	16'h	428f;
13835	:douta	=	16'h	5310;
13836	:douta	=	16'h	42af;
13837	:douta	=	16'h	4b10;
13838	:douta	=	16'h	6392;
13839	:douta	=	16'h	6bb2;
13840	:douta	=	16'h	a557;
13841	:douta	=	16'h	a557;
13842	:douta	=	16'h	bd96;
13843	:douta	=	16'h	b556;
13844	:douta	=	16'h	bdb6;
13845	:douta	=	16'h	6b6f;
13846	:douta	=	16'h	9450;
13847	:douta	=	16'h	acf2;
13848	:douta	=	16'h	bdb4;
13849	:douta	=	16'h	9451;
13850	:douta	=	16'h	a4f2;
13851	:douta	=	16'h	b533;
13852	:douta	=	16'h	8c2f;
13853	:douta	=	16'h	736d;
13854	:douta	=	16'h	9c91;
13855	:douta	=	16'h	b532;
13856	:douta	=	16'h	bd73;
13857	:douta	=	16'h	c593;
13858	:douta	=	16'h	e6b7;
13859	:douta	=	16'h	cdf4;
13860	:douta	=	16'h	9cb0;
13861	:douta	=	16'h	8c0d;
13862	:douta	=	16'h	bdb3;
13863	:douta	=	16'h	e6b6;
13864	:douta	=	16'h	b592;
13865	:douta	=	16'h	7b2a;
13866	:douta	=	16'h	7b4a;
13867	:douta	=	16'h	93cb;
13868	:douta	=	16'h	93cb;
13869	:douta	=	16'h	93cc;
13870	:douta	=	16'h	ac6c;
13871	:douta	=	16'h	ac8d;
13872	:douta	=	16'h	b4ad;
13873	:douta	=	16'h	c50e;
13874	:douta	=	16'h	cd6f;
13875	:douta	=	16'h	d5b1;
13876	:douta	=	16'h	d591;
13877	:douta	=	16'h	ddd2;
13878	:douta	=	16'h	ddf2;
13879	:douta	=	16'h	ddd2;
13880	:douta	=	16'h	ddf2;
13881	:douta	=	16'h	ddd1;
13882	:douta	=	16'h	ddd1;
13883	:douta	=	16'h	e613;
13884	:douta	=	16'h	e654;
13885	:douta	=	16'h	cd4f;
13886	:douta	=	16'h	c50f;
13887	:douta	=	16'h	8c0f;
13888	:douta	=	16'h	4a08;
13889	:douta	=	16'h	7b2a;
13890	:douta	=	16'h	7bce;
13891	:douta	=	16'h	4a6b;
13892	:douta	=	16'h	31a8;
13893	:douta	=	16'h	6b0c;
13894	:douta	=	16'h	4a4a;
13895	:douta	=	16'h	2166;
13896	:douta	=	16'h	2126;
13897	:douta	=	16'h	1906;
13898	:douta	=	16'h	2125;
13899	:douta	=	16'h	1905;
13900	:douta	=	16'h	10e4;
13901	:douta	=	16'h	1904;
13902	:douta	=	16'h	2125;
13903	:douta	=	16'h	0000;
13904	:douta	=	16'h	0000;
13905	:douta	=	16'h	0022;
13906	:douta	=	16'h	0062;
13907	:douta	=	16'h	5b2f;
13908	:douta	=	16'h	29c9;
13909	:douta	=	16'h	1926;
13910	:douta	=	16'h	2126;
13911	:douta	=	16'h	83cd;
13912	:douta	=	16'h	5269;
13913	:douta	=	16'h	62aa;
13914	:douta	=	16'h	632c;
13915	:douta	=	16'h	2146;
13916	:douta	=	16'h	31c9;
13917	:douta	=	16'h	2168;
13918	:douta	=	16'h	21a8;
13919	:douta	=	16'h	2147;
13920	:douta	=	16'h	324a;
13921	:douta	=	16'h	00a5;
13922	:douta	=	16'h	73b0;
13923	:douta	=	16'h	4aad;
13924	:douta	=	16'h	322c;
13925	:douta	=	16'h	322a;
13926	:douta	=	16'h	324c;
13927	:douta	=	16'h	1968;
13928	:douta	=	16'h	29a9;
13929	:douta	=	16'h	5aec;
13930	:douta	=	16'h	2189;
13931	:douta	=	16'h	3a09;
13932	:douta	=	16'h	320b;
13933	:douta	=	16'h	426c;
13934	:douta	=	16'h	1969;
13935	:douta	=	16'h	2189;
13936	:douta	=	16'h	29ec;
13937	:douta	=	16'h	324d;
13938	:douta	=	16'h	0908;
13939	:douta	=	16'h	198a;
13940	:douta	=	16'h	322c;
13941	:douta	=	16'h	218a;
13942	:douta	=	16'h	8bab;
13943	:douta	=	16'h	52cd;
13944	:douta	=	16'h	957a;
13945	:douta	=	16'h	6c76;
13946	:douta	=	16'h	7497;
13947	:douta	=	16'h	84d8;
13948	:douta	=	16'h	8d19;
13949	:douta	=	16'h	84d8;
13950	:douta	=	16'h	7cb8;
13951	:douta	=	16'h	959b;
13952	:douta	=	16'h	6c36;
13953	:douta	=	16'h	6c57;
13954	:douta	=	16'h	84f9;
13955	:douta	=	16'h	957a;
13956	:douta	=	16'h	8518;
13957	:douta	=	16'h	8d39;
13958	:douta	=	16'h	7457;
13959	:douta	=	16'h	84f9;
13960	:douta	=	16'h	84f9;
13961	:douta	=	16'h	84f9;
13962	:douta	=	16'h	853a;
13963	:douta	=	16'h	7497;
13964	:douta	=	16'h	84f9;
13965	:douta	=	16'h	8d39;
13966	:douta	=	16'h	8d79;
13967	:douta	=	16'h	7cd8;
13968	:douta	=	16'h	7cb8;
13969	:douta	=	16'h	7cb8;
13970	:douta	=	16'h	8519;
13971	:douta	=	16'h	9d9b;
13972	:douta	=	16'h	9ddc;
13973	:douta	=	16'h	a5db;
13974	:douta	=	16'h	7cd9;
13975	:douta	=	16'h	8d7a;
13976	:douta	=	16'h	8519;
13977	:douta	=	16'h	a5dc;
13978	:douta	=	16'h	9ddb;
13979	:douta	=	16'h	8519;
13980	:douta	=	16'h	84f8;
13981	:douta	=	16'h	84f9;
13982	:douta	=	16'h	8539;
13983	:douta	=	16'h	959b;
13984	:douta	=	16'h	7498;
13985	:douta	=	16'h	6c98;
13986	:douta	=	16'h	6437;
13987	:douta	=	16'h	6c77;
13988	:douta	=	16'h	5c37;
13989	:douta	=	16'h	95bb;
13990	:douta	=	16'h	959b;
13991	:douta	=	16'h	8d5a;
13992	:douta	=	16'h	74b8;
13993	:douta	=	16'h	95bc;
13994	:douta	=	16'h	5bd5;
13995	:douta	=	16'h	6416;
13996	:douta	=	16'h	9dbb;
13997	:douta	=	16'h	8d3a;
13998	:douta	=	16'h	84f9;
13999	:douta	=	16'h	8d5b;
14000	:douta	=	16'h	855a;
14001	:douta	=	16'h	7477;
14002	:douta	=	16'h	7cd9;
14003	:douta	=	16'h	7cd9;
14004	:douta	=	16'h	8d7b;
14005	:douta	=	16'h	8d9c;
14006	:douta	=	16'h	74b8;
14007	:douta	=	16'h	5bd4;
14008	:douta	=	16'h	6c36;
14009	:douta	=	16'h	853a;
14010	:douta	=	16'h	7cf9;
14011	:douta	=	16'h	5bb4;
14012	:douta	=	16'h	7cd9;
14013	:douta	=	16'h	851a;
14014	:douta	=	16'h	6c57;
14015	:douta	=	16'h	5bb4;
14016	:douta	=	16'h	7cf9;
14017	:douta	=	16'h	74b8;
14018	:douta	=	16'h	855b;
14019	:douta	=	16'h	7477;
14020	:douta	=	16'h	7457;
14021	:douta	=	16'h	6436;
14022	:douta	=	16'h	5bd4;
14023	:douta	=	16'h	6c97;
14024	:douta	=	16'h	6415;
14025	:douta	=	16'h	6415;
14026	:douta	=	16'h	6415;
14027	:douta	=	16'h	7498;
14028	:douta	=	16'h	74b8;
14029	:douta	=	16'h	5bb4;
14030	:douta	=	16'h	6416;
14031	:douta	=	16'h	7cd9;
14032	:douta	=	16'h	74f9;
14033	:douta	=	16'h	7cf9;
14034	:douta	=	16'h	7d1a;
14035	:douta	=	16'h	7cfa;
14036	:douta	=	16'h	855b;
14037	:douta	=	16'h	855b;
14038	:douta	=	16'h	857b;
14039	:douta	=	16'h	853c;
14040	:douta	=	16'h	7d1a;
14041	:douta	=	16'h	7d3b;
14042	:douta	=	16'h	74da;
14043	:douta	=	16'h	7cfb;
14044	:douta	=	16'h	8dbd;
14045	:douta	=	16'h	857c;
14046	:douta	=	16'h	8d7c;
14047	:douta	=	16'h	74b9;
14048	:douta	=	16'h	7cfa;
14049	:douta	=	16'h	7d3a;
14050	:douta	=	16'h	6cb9;
14051	:douta	=	16'h	74fa;
14052	:douta	=	16'h	7d3a;
14053	:douta	=	16'h	857b;
14054	:douta	=	16'h	7cfa;
14055	:douta	=	16'h	7d1a;
14056	:douta	=	16'h	7d3a;
14057	:douta	=	16'h	8d9c;
14058	:douta	=	16'h	74fa;
14059	:douta	=	16'h	6458;
14060	:douta	=	16'h	5c37;
14061	:douta	=	16'h	857b;
14062	:douta	=	16'h	857b;
14063	:douta	=	16'h	857b;
14064	:douta	=	16'h	855b;
14065	:douta	=	16'h	855b;
14066	:douta	=	16'h	8dbc;
14067	:douta	=	16'h	751a;
14068	:douta	=	16'h	74d9;
14069	:douta	=	16'h	7498;
14070	:douta	=	16'h	3a4c;
14071	:douta	=	16'h	7474;
14072	:douta	=	16'h	8cb5;
14073	:douta	=	16'h	7c54;
14074	:douta	=	16'h	4b0f;
14075	:douta	=	16'h	42ae;
14076	:douta	=	16'h	6391;
14077	:douta	=	16'h	ad55;
14078	:douta	=	16'h	9d15;
14079	:douta	=	16'h	3a8d;
14080	:douta	=	16'h	222f;
14081	:douta	=	16'h	3b32;
14082	:douta	=	16'h	32d1;
14083	:douta	=	16'h	2a2e;
14084	:douta	=	16'h	4333;
14085	:douta	=	16'h	6417;
14086	:douta	=	16'h	5393;
14087	:douta	=	16'h	84b8;
14088	:douta	=	16'h	4b10;
14089	:douta	=	16'h	6c76;
14090	:douta	=	16'h	42af;
14091	:douta	=	16'h	7c75;
14092	:douta	=	16'h	7454;
14093	:douta	=	16'h	8cd7;
14094	:douta	=	16'h	94d6;
14095	:douta	=	16'h	9d16;
14096	:douta	=	16'h	8c95;
14097	:douta	=	16'h	8475;
14098	:douta	=	16'h	5b2f;
14099	:douta	=	16'h	7bf1;
14100	:douta	=	16'h	9cf3;
14101	:douta	=	16'h	c5b5;
14102	:douta	=	16'h	cdd6;
14103	:douta	=	16'h	c5f5;
14104	:douta	=	16'h	9cd2;
14105	:douta	=	16'h	632c;
14106	:douta	=	16'h	62cb;
14107	:douta	=	16'h	8bee;
14108	:douta	=	16'h	83ee;
14109	:douta	=	16'h	a4d1;
14110	:douta	=	16'h	ce36;
14111	:douta	=	16'h	eef8;
14112	:douta	=	16'h	d677;
14113	:douta	=	16'h	732b;
14114	:douta	=	16'h	bd92;
14115	:douta	=	16'h	b531;
14116	:douta	=	16'h	bdb3;
14117	:douta	=	16'h	946d;
14118	:douta	=	16'h	ff7a;
14119	:douta	=	16'h	6ae9;
14120	:douta	=	16'h	7b0a;
14121	:douta	=	16'h	72ea;
14122	:douta	=	16'h	8b8b;
14123	:douta	=	16'h	93eb;
14124	:douta	=	16'h	9bec;
14125	:douta	=	16'h	93cb;
14126	:douta	=	16'h	ac6c;
14127	:douta	=	16'h	b48d;
14128	:douta	=	16'h	bccd;
14129	:douta	=	16'h	cd6f;
14130	:douta	=	16'h	cd70;
14131	:douta	=	16'h	ddf3;
14132	:douta	=	16'h	e613;
14133	:douta	=	16'h	de13;
14134	:douta	=	16'h	de13;
14135	:douta	=	16'h	e634;
14136	:douta	=	16'h	ddf3;
14137	:douta	=	16'h	ddf3;
14138	:douta	=	16'h	e633;
14139	:douta	=	16'h	cd6f;
14140	:douta	=	16'h	cd90;
14141	:douta	=	16'h	e653;
14142	:douta	=	16'h	b4f0;
14143	:douta	=	16'h	3165;
14144	:douta	=	16'h	a46f;
14145	:douta	=	16'h	acd0;
14146	:douta	=	16'h	62eb;
14147	:douta	=	16'h	39e9;
14148	:douta	=	16'h	4209;
14149	:douta	=	16'h	6aeb;
14150	:douta	=	16'h	39e9;
14151	:douta	=	16'h	29a8;
14152	:douta	=	16'h	29a8;
14153	:douta	=	16'h	2126;
14154	:douta	=	16'h	2946;
14155	:douta	=	16'h	10a3;
14156	:douta	=	16'h	1905;
14157	:douta	=	16'h	18e4;
14158	:douta	=	16'h	18e4;
14159	:douta	=	16'h	2145;
14160	:douta	=	16'h	0883;
14161	:douta	=	16'h	0001;
14162	:douta	=	16'h	0022;
14163	:douta	=	16'h	1106;
14164	:douta	=	16'h	1968;
14165	:douta	=	16'h	1905;
14166	:douta	=	16'h	1926;
14167	:douta	=	16'h	10e5;
14168	:douta	=	16'h	08c4;
14169	:douta	=	16'h	0842;
14170	:douta	=	16'h	4a48;
14171	:douta	=	16'h	4208;
14172	:douta	=	16'h	2966;
14173	:douta	=	16'h	4208;
14174	:douta	=	16'h	8c0e;
14175	:douta	=	16'h	630d;
14176	:douta	=	16'h	324d;
14177	:douta	=	16'h	4aac;
14178	:douta	=	16'h	21cb;
14179	:douta	=	16'h	1948;
14180	:douta	=	16'h	29a9;
14181	:douta	=	16'h	31c9;
14182	:douta	=	16'h	320a;
14183	:douta	=	16'h	4aab;
14184	:douta	=	16'h	29ca;
14185	:douta	=	16'h	8410;
14186	:douta	=	16'h	29a9;
14187	:douta	=	16'h	3a09;
14188	:douta	=	16'h	29a8;
14189	:douta	=	16'h	1947;
14190	:douta	=	16'h	4acc;
14191	:douta	=	16'h	29ca;
14192	:douta	=	16'h	322a;
14193	:douta	=	16'h	3187;
14194	:douta	=	16'h	8452;
14195	:douta	=	16'h	530f;
14196	:douta	=	16'h	32af;
14197	:douta	=	16'h	6ace;
14198	:douta	=	16'h	5aed;
14199	:douta	=	16'h	a598;
14200	:douta	=	16'h	959b;
14201	:douta	=	16'h	6436;
14202	:douta	=	16'h	8519;
14203	:douta	=	16'h	9dbb;
14204	:douta	=	16'h	8d38;
14205	:douta	=	16'h	8519;
14206	:douta	=	16'h	8d5a;
14207	:douta	=	16'h	8519;
14208	:douta	=	16'h	addc;
14209	:douta	=	16'h	9d9a;
14210	:douta	=	16'h	7477;
14211	:douta	=	16'h	7cd8;
14212	:douta	=	16'h	84f9;
14213	:douta	=	16'h	6c56;
14214	:douta	=	16'h	8d19;
14215	:douta	=	16'h	a5dc;
14216	:douta	=	16'h	5bb4;
14217	:douta	=	16'h	5bf5;
14218	:douta	=	16'h	8519;
14219	:douta	=	16'h	9dbb;
14220	:douta	=	16'h	8539;
14221	:douta	=	16'h	8519;
14222	:douta	=	16'h	84d9;
14223	:douta	=	16'h	9559;
14224	:douta	=	16'h	8d7a;
14225	:douta	=	16'h	8d39;
14226	:douta	=	16'h	959b;
14227	:douta	=	16'h	8d3a;
14228	:douta	=	16'h	957a;
14229	:douta	=	16'h	7cd8;
14230	:douta	=	16'h	a5db;
14231	:douta	=	16'h	853a;
14232	:douta	=	16'h	8519;
14233	:douta	=	16'h	957a;
14234	:douta	=	16'h	8d3a;
14235	:douta	=	16'h	959a;
14236	:douta	=	16'h	84d8;
14237	:douta	=	16'h	84f9;
14238	:douta	=	16'h	84f9;
14239	:douta	=	16'h	7cd9;
14240	:douta	=	16'h	853a;
14241	:douta	=	16'h	ae1c;
14242	:douta	=	16'h	957a;
14243	:douta	=	16'h	6417;
14244	:douta	=	16'h	74b8;
14245	:douta	=	16'h	851a;
14246	:douta	=	16'h	74b8;
14247	:douta	=	16'h	959b;
14248	:douta	=	16'h	9d9c;
14249	:douta	=	16'h	84f9;
14250	:douta	=	16'h	7cd8;
14251	:douta	=	16'h	955a;
14252	:douta	=	16'h	5bd5;
14253	:douta	=	16'h	53b4;
14254	:douta	=	16'h	5c16;
14255	:douta	=	16'h	853a;
14256	:douta	=	16'h	7d3a;
14257	:douta	=	16'h	6cb8;
14258	:douta	=	16'h	7d1a;
14259	:douta	=	16'h	7d3b;
14260	:douta	=	16'h	7498;
14261	:douta	=	16'h	7cd9;
14262	:douta	=	16'h	74d9;
14263	:douta	=	16'h	7d1a;
14264	:douta	=	16'h	7cf9;
14265	:douta	=	16'h	6c36;
14266	:douta	=	16'h	5bf5;
14267	:douta	=	16'h	6c57;
14268	:douta	=	16'h	8d39;
14269	:douta	=	16'h	7477;
14270	:douta	=	16'h	6c56;
14271	:douta	=	16'h	6c77;
14272	:douta	=	16'h	7cd9;
14273	:douta	=	16'h	7cf9;
14274	:douta	=	16'h	5b94;
14275	:douta	=	16'h	6436;
14276	:douta	=	16'h	6cb8;
14277	:douta	=	16'h	7498;
14278	:douta	=	16'h	7456;
14279	:douta	=	16'h	6c15;
14280	:douta	=	16'h	63f5;
14281	:douta	=	16'h	853a;
14282	:douta	=	16'h	6c77;
14283	:douta	=	16'h	6415;
14284	:douta	=	16'h	63f4;
14285	:douta	=	16'h	5bd4;
14286	:douta	=	16'h	5bd5;
14287	:douta	=	16'h	6c78;
14288	:douta	=	16'h	6c98;
14289	:douta	=	16'h	855a;
14290	:douta	=	16'h	74d9;
14291	:douta	=	16'h	6c78;
14292	:douta	=	16'h	6c78;
14293	:douta	=	16'h	8d9c;
14294	:douta	=	16'h	855b;
14295	:douta	=	16'h	855c;
14296	:douta	=	16'h	857c;
14297	:douta	=	16'h	74fa;
14298	:douta	=	16'h	855c;
14299	:douta	=	16'h	859c;
14300	:douta	=	16'h	7cfa;
14301	:douta	=	16'h	7d3a;
14302	:douta	=	16'h	855b;
14303	:douta	=	16'h	7cfa;
14304	:douta	=	16'h	7d3b;
14305	:douta	=	16'h	855c;
14306	:douta	=	16'h	855b;
14307	:douta	=	16'h	857b;
14308	:douta	=	16'h	6c98;
14309	:douta	=	16'h	74d9;
14310	:douta	=	16'h	7d1a;
14311	:douta	=	16'h	7d1a;
14312	:douta	=	16'h	8d9c;
14313	:douta	=	16'h	6c99;
14314	:douta	=	16'h	6478;
14315	:douta	=	16'h	857c;
14316	:douta	=	16'h	8dbc;
14317	:douta	=	16'h	53f6;
14318	:douta	=	16'h	6458;
14319	:douta	=	16'h	7d3a;
14320	:douta	=	16'h	7d5b;
14321	:douta	=	16'h	857b;
14322	:douta	=	16'h	74d9;
14323	:douta	=	16'h	8dbc;
14324	:douta	=	16'h	857c;
14325	:douta	=	16'h	7d1b;
14326	:douta	=	16'h	5b73;
14327	:douta	=	16'h	52cd;
14328	:douta	=	16'h	5350;
14329	:douta	=	16'h	8453;
14330	:douta	=	16'h	8cb5;
14331	:douta	=	16'h	63b2;
14332	:douta	=	16'h	8c73;
14333	:douta	=	16'h	42cf;
14334	:douta	=	16'h	21aa;
14335	:douta	=	16'h	73d2;
14336	:douta	=	16'h	3b33;
14337	:douta	=	16'h	4354;
14338	:douta	=	16'h	4bd6;
14339	:douta	=	16'h	198b;
14340	:douta	=	16'h	3b12;
14341	:douta	=	16'h	3ad1;
14342	:douta	=	16'h	42d0;
14343	:douta	=	16'h	5352;
14344	:douta	=	16'h	6c35;
14345	:douta	=	16'h	6c16;
14346	:douta	=	16'h	6bf4;
14347	:douta	=	16'h	5b51;
14348	:douta	=	16'h	6bf3;
14349	:douta	=	16'h	6bf4;
14350	:douta	=	16'h	7413;
14351	:douta	=	16'h	9d17;
14352	:douta	=	16'h	9d36;
14353	:douta	=	16'h	a578;
14354	:douta	=	16'h	9493;
14355	:douta	=	16'h	7c11;
14356	:douta	=	16'h	73b0;
14357	:douta	=	16'h	8c30;
14358	:douta	=	16'h	9c71;
14359	:douta	=	16'h	b574;
14360	:douta	=	16'h	e677;
14361	:douta	=	16'h	b573;
14362	:douta	=	16'h	b553;
14363	:douta	=	16'h	a4d1;
14364	:douta	=	16'h	730c;
14365	:douta	=	16'h	4a6b;
14366	:douta	=	16'h	8c30;
14367	:douta	=	16'h	ad12;
14368	:douta	=	16'h	e696;
14369	:douta	=	16'h	a4f1;
14370	:douta	=	16'h	eef8;
14371	:douta	=	16'h	c5d3;
14372	:douta	=	16'h	8c4f;
14373	:douta	=	16'h	4a49;
14374	:douta	=	16'h	ce14;
14375	:douta	=	16'h	6ac9;
14376	:douta	=	16'h	732a;
14377	:douta	=	16'h	7b4a;
14378	:douta	=	16'h	93ab;
14379	:douta	=	16'h	93eb;
14380	:douta	=	16'h	9c0c;
14381	:douta	=	16'h	9beb;
14382	:douta	=	16'h	b48d;
14383	:douta	=	16'h	bccd;
14384	:douta	=	16'h	bced;
14385	:douta	=	16'h	d590;
14386	:douta	=	16'h	d5b1;
14387	:douta	=	16'h	ddf2;
14388	:douta	=	16'h	de33;
14389	:douta	=	16'h	e634;
14390	:douta	=	16'h	ddf2;
14391	:douta	=	16'h	ddf3;
14392	:douta	=	16'h	e613;
14393	:douta	=	16'h	de13;
14394	:douta	=	16'h	de12;
14395	:douta	=	16'h	c56f;
14396	:douta	=	16'h	c50f;
14397	:douta	=	16'h	ddd1;
14398	:douta	=	16'h	c531;
14399	:douta	=	16'h	6aa9;
14400	:douta	=	16'h	9c2e;
14401	:douta	=	16'h	a48e;
14402	:douta	=	16'h	5acb;
14403	:douta	=	16'h	29a9;
14404	:douta	=	16'h	62cb;
14405	:douta	=	16'h	6b0b;
14406	:douta	=	16'h	4229;
14407	:douta	=	16'h	31a8;
14408	:douta	=	16'h	2967;
14409	:douta	=	16'h	1925;
14410	:douta	=	16'h	4229;
14411	:douta	=	16'h	2966;
14412	:douta	=	16'h	1904;
14413	:douta	=	16'h	10e4;
14414	:douta	=	16'h	10e4;
14415	:douta	=	16'h	18c4;
14416	:douta	=	16'h	1905;
14417	:douta	=	16'h	0000;
14418	:douta	=	16'h	0001;
14419	:douta	=	16'h	10a5;
14420	:douta	=	16'h	2a0b;
14421	:douta	=	16'h	21c9;
14422	:douta	=	16'h	10e5;
14423	:douta	=	16'h	10e5;
14424	:douta	=	16'h	1946;
14425	:douta	=	16'h	62a9;
14426	:douta	=	16'h	630a;
14427	:douta	=	16'h	62ea;
14428	:douta	=	16'h	41e7;
14429	:douta	=	16'h	1084;
14430	:douta	=	16'h	4249;
14431	:douta	=	16'h	6b2b;
14432	:douta	=	16'h	320b;
14433	:douta	=	16'h	52ac;
14434	:douta	=	16'h	4aee;
14435	:douta	=	16'h	29ea;
14436	:douta	=	16'h	3a2b;
14437	:douta	=	16'h	1149;
14438	:douta	=	16'h	1148;
14439	:douta	=	16'h	1127;
14440	:douta	=	16'h	0084;
14441	:douta	=	16'h	5acb;
14442	:douta	=	16'h	426b;
14443	:douta	=	16'h	52ac;
14444	:douta	=	16'h	29a9;
14445	:douta	=	16'h	52ec;
14446	:douta	=	16'h	29ea;
14447	:douta	=	16'h	3a2c;
14448	:douta	=	16'h	1148;
14449	:douta	=	16'h	1926;
14450	:douta	=	16'h	29ea;
14451	:douta	=	16'h	31a9;
14452	:douta	=	16'h	21cb;
14453	:douta	=	16'h	8bae;
14454	:douta	=	16'h	5b0d;
14455	:douta	=	16'h	9dba;
14456	:douta	=	16'h	6c77;
14457	:douta	=	16'h	8d19;
14458	:douta	=	16'h	84f9;
14459	:douta	=	16'h	9d9a;
14460	:douta	=	16'h	9d9a;
14461	:douta	=	16'h	84f9;
14462	:douta	=	16'h	7cd8;
14463	:douta	=	16'h	8d19;
14464	:douta	=	16'h	a5bb;
14465	:douta	=	16'h	a5da;
14466	:douta	=	16'h	957a;
14467	:douta	=	16'h	8d19;
14468	:douta	=	16'h	7477;
14469	:douta	=	16'h	7cb8;
14470	:douta	=	16'h	8519;
14471	:douta	=	16'h	7477;
14472	:douta	=	16'h	959b;
14473	:douta	=	16'h	7c97;
14474	:douta	=	16'h	6c36;
14475	:douta	=	16'h	6c36;
14476	:douta	=	16'h	7498;
14477	:douta	=	16'h	8d39;
14478	:douta	=	16'h	84d8;
14479	:douta	=	16'h	8519;
14480	:douta	=	16'h	8d39;
14481	:douta	=	16'h	8d39;
14482	:douta	=	16'h	8d39;
14483	:douta	=	16'h	8d39;
14484	:douta	=	16'h	a5fb;
14485	:douta	=	16'h	ae1c;
14486	:douta	=	16'h	957a;
14487	:douta	=	16'h	6c77;
14488	:douta	=	16'h	8d59;
14489	:douta	=	16'h	a5bb;
14490	:douta	=	16'h	959a;
14491	:douta	=	16'h	8d19;
14492	:douta	=	16'h	9d9a;
14493	:douta	=	16'h	8d5a;
14494	:douta	=	16'h	7cd8;
14495	:douta	=	16'h	7477;
14496	:douta	=	16'h	7cf9;
14497	:douta	=	16'h	7498;
14498	:douta	=	16'h	a5fc;
14499	:douta	=	16'h	8d59;
14500	:douta	=	16'h	6c56;
14501	:douta	=	16'h	7497;
14502	:douta	=	16'h	6416;
14503	:douta	=	16'h	6c77;
14504	:douta	=	16'h	7cb8;
14505	:douta	=	16'h	9ddc;
14506	:douta	=	16'h	8d39;
14507	:douta	=	16'h	8d3a;
14508	:douta	=	16'h	853a;
14509	:douta	=	16'h	53b5;
14510	:douta	=	16'h	5394;
14511	:douta	=	16'h	6cda;
14512	:douta	=	16'h	6cb9;
14513	:douta	=	16'h	7cfa;
14514	:douta	=	16'h	6457;
14515	:douta	=	16'h	6c98;
14516	:douta	=	16'h	7d3a;
14517	:douta	=	16'h	7d1a;
14518	:douta	=	16'h	74b8;
14519	:douta	=	16'h	74b8;
14520	:douta	=	16'h	6c77;
14521	:douta	=	16'h	7cd8;
14522	:douta	=	16'h	7cb8;
14523	:douta	=	16'h	6c15;
14524	:douta	=	16'h	7477;
14525	:douta	=	16'h	7497;
14526	:douta	=	16'h	84d8;
14527	:douta	=	16'h	7476;
14528	:douta	=	16'h	6c14;
14529	:douta	=	16'h	7477;
14530	:douta	=	16'h	84d9;
14531	:douta	=	16'h	5b73;
14532	:douta	=	16'h	5b73;
14533	:douta	=	16'h	6477;
14534	:douta	=	16'h	7cf8;
14535	:douta	=	16'h	7cb8;
14536	:douta	=	16'h	4b31;
14537	:douta	=	16'h	4b32;
14538	:douta	=	16'h	7cb8;
14539	:douta	=	16'h	6c56;
14540	:douta	=	16'h	7497;
14541	:douta	=	16'h	6c57;
14542	:douta	=	16'h	5bf5;
14543	:douta	=	16'h	4b94;
14544	:douta	=	16'h	6417;
14545	:douta	=	16'h	53d5;
14546	:douta	=	16'h	855b;
14547	:douta	=	16'h	7d1a;
14548	:douta	=	16'h	74fa;
14549	:douta	=	16'h	855b;
14550	:douta	=	16'h	857c;
14551	:douta	=	16'h	7d3b;
14552	:douta	=	16'h	7cfb;
14553	:douta	=	16'h	74da;
14554	:douta	=	16'h	7d3b;
14555	:douta	=	16'h	751b;
14556	:douta	=	16'h	7d1b;
14557	:douta	=	16'h	7d5b;
14558	:douta	=	16'h	7cfa;
14559	:douta	=	16'h	7d1a;
14560	:douta	=	16'h	6c98;
14561	:douta	=	16'h	7d3a;
14562	:douta	=	16'h	7d3a;
14563	:douta	=	16'h	857b;
14564	:douta	=	16'h	7cfa;
14565	:douta	=	16'h	7cda;
14566	:douta	=	16'h	74b9;
14567	:douta	=	16'h	7cfa;
14568	:douta	=	16'h	74d9;
14569	:douta	=	16'h	95dd;
14570	:douta	=	16'h	855b;
14571	:douta	=	16'h	74d9;
14572	:douta	=	16'h	7d1a;
14573	:douta	=	16'h	95bc;
14574	:douta	=	16'h	6437;
14575	:douta	=	16'h	7499;
14576	:douta	=	16'h	855b;
14577	:douta	=	16'h	8dbd;
14578	:douta	=	16'h	855b;
14579	:douta	=	16'h	7d5b;
14580	:douta	=	16'h	7d3b;
14581	:douta	=	16'h	7d1b;
14582	:douta	=	16'h	6c77;
14583	:douta	=	16'h	532f;
14584	:douta	=	16'h	7412;
14585	:douta	=	16'h	7c33;
14586	:douta	=	16'h	5330;
14587	:douta	=	16'h	6bd2;
14588	:douta	=	16'h	9493;
14589	:douta	=	16'h	8cb4;
14590	:douta	=	16'h	6391;
14591	:douta	=	16'h	7c53;
14592	:douta	=	16'h	19ed;
14593	:douta	=	16'h	3312;
14594	:douta	=	16'h	2ad0;
14595	:douta	=	16'h	2a50;
14596	:douta	=	16'h	4332;
14597	:douta	=	16'h	5bf6;
14598	:douta	=	16'h	53b4;
14599	:douta	=	16'h	7c97;
14600	:douta	=	16'h	6c36;
14601	:douta	=	16'h	7c97;
14602	:douta	=	16'h	5372;
14603	:douta	=	16'h	4acf;
14604	:douta	=	16'h	5311;
14605	:douta	=	16'h	5b92;
14606	:douta	=	16'h	7413;
14607	:douta	=	16'h	8454;
14608	:douta	=	16'h	b5b8;
14609	:douta	=	16'h	8c94;
14610	:douta	=	16'h	73f1;
14611	:douta	=	16'h	8c71;
14612	:douta	=	16'h	ad34;
14613	:douta	=	16'h	7bd0;
14614	:douta	=	16'h	cdb6;
14615	:douta	=	16'h	bd74;
14616	:douta	=	16'h	83ef;
14617	:douta	=	16'h	7b8e;
14618	:douta	=	16'h	bd73;
14619	:douta	=	16'h	d635;
14620	:douta	=	16'h	c593;
14621	:douta	=	16'h	7bce;
14622	:douta	=	16'h	a4b1;
14623	:douta	=	16'h	bd52;
14624	:douta	=	16'h	d614;
14625	:douta	=	16'h	738c;
14626	:douta	=	16'h	acaf;
14627	:douta	=	16'h	8c2d;
14628	:douta	=	16'h	bd72;
14629	:douta	=	16'h	9c90;
14630	:douta	=	16'h	7b6b;
14631	:douta	=	16'h	730a;
14632	:douta	=	16'h	834a;
14633	:douta	=	16'h	8bab;
14634	:douta	=	16'h	93cb;
14635	:douta	=	16'h	a40c;
14636	:douta	=	16'h	a42b;
14637	:douta	=	16'h	ac6c;
14638	:douta	=	16'h	b4ad;
14639	:douta	=	16'h	c50e;
14640	:douta	=	16'h	d570;
14641	:douta	=	16'h	ddd2;
14642	:douta	=	16'h	ddf2;
14643	:douta	=	16'h	de33;
14644	:douta	=	16'h	de33;
14645	:douta	=	16'h	e654;
14646	:douta	=	16'h	ddf2;
14647	:douta	=	16'h	ddd2;
14648	:douta	=	16'h	ddf2;
14649	:douta	=	16'h	ddf3;
14650	:douta	=	16'h	d591;
14651	:douta	=	16'h	bcce;
14652	:douta	=	16'h	ac6e;
14653	:douta	=	16'h	ac4d;
14654	:douta	=	16'h	9bec;
14655	:douta	=	16'h	a46e;
14656	:douta	=	16'h	940d;
14657	:douta	=	16'h	a46e;
14658	:douta	=	16'h	52aa;
14659	:douta	=	16'h	39ea;
14660	:douta	=	16'h	7b8d;
14661	:douta	=	16'h	734c;
14662	:douta	=	16'h	5aaa;
14663	:douta	=	16'h	39c9;
14664	:douta	=	16'h	31e9;
14665	:douta	=	16'h	2188;
14666	:douta	=	16'h	1126;
14667	:douta	=	16'h	2967;
14668	:douta	=	16'h	1905;
14669	:douta	=	16'h	0883;
14670	:douta	=	16'h	10c4;
14671	:douta	=	16'h	10e4;
14672	:douta	=	16'h	10e4;
14673	:douta	=	16'h	1905;
14674	:douta	=	16'h	0001;
14675	:douta	=	16'h	0042;
14676	:douta	=	16'h	0863;
14677	:douta	=	16'h	2168;
14678	:douta	=	16'h	1968;
14679	:douta	=	16'h	18e5;
14680	:douta	=	16'h	10e5;
14681	:douta	=	16'h	18e6;
14682	:douta	=	16'h	10a4;
14683	:douta	=	16'h	18e4;
14684	:douta	=	16'h	08a3;
14685	:douta	=	16'h	944e;
14686	:douta	=	16'h	52aa;
14687	:douta	=	16'h	9c8f;
14688	:douta	=	16'h	4a2a;
14689	:douta	=	16'h	5b0c;
14690	:douta	=	16'h	3a4c;
14691	:douta	=	16'h	320b;
14692	:douta	=	16'h	08c5;
14693	:douta	=	16'h	530d;
14694	:douta	=	16'h	424b;
14695	:douta	=	16'h	29ea;
14696	:douta	=	16'h	52cc;
14697	:douta	=	16'h	3a4c;
14698	:douta	=	16'h	634d;
14699	:douta	=	16'h	322a;
14700	:douta	=	16'h	39e9;
14701	:douta	=	16'h	1127;
14702	:douta	=	16'h	0885;
14703	:douta	=	16'h	1969;
14704	:douta	=	16'h	08c6;
14705	:douta	=	16'h	5b0c;
14706	:douta	=	16'h	4aab;
14707	:douta	=	16'h	39c8;
14708	:douta	=	16'h	31a8;
14709	:douta	=	16'h	ac6f;
14710	:douta	=	16'h	8434;
14711	:douta	=	16'h	8d7a;
14712	:douta	=	16'h	8d7a;
14713	:douta	=	16'h	6c56;
14714	:douta	=	16'h	63f5;
14715	:douta	=	16'h	5b93;
14716	:douta	=	16'h	3ad1;
14717	:douta	=	16'h	5353;
14718	:douta	=	16'h	8d19;
14719	:douta	=	16'h	8d19;
14720	:douta	=	16'h	7cb8;
14721	:douta	=	16'h	74b7;
14722	:douta	=	16'h	8518;
14723	:douta	=	16'h	9d7b;
14724	:douta	=	16'h	959b;
14725	:douta	=	16'h	7497;
14726	:douta	=	16'h	7cb8;
14727	:douta	=	16'h	9ddc;
14728	:douta	=	16'h	84f9;
14729	:douta	=	16'h	7cd9;
14730	:douta	=	16'h	6c77;
14731	:douta	=	16'h	955a;
14732	:douta	=	16'h	8d59;
14733	:douta	=	16'h	7478;
14734	:douta	=	16'h	7cb8;
14735	:douta	=	16'h	84f9;
14736	:douta	=	16'h	9dbb;
14737	:douta	=	16'h	8d5a;
14738	:douta	=	16'h	8d59;
14739	:douta	=	16'h	a5db;
14740	:douta	=	16'h	957a;
14741	:douta	=	16'h	9559;
14742	:douta	=	16'h	955a;
14743	:douta	=	16'h	a5fb;
14744	:douta	=	16'h	a5fc;
14745	:douta	=	16'h	6c77;
14746	:douta	=	16'h	7cf8;
14747	:douta	=	16'h	8d7a;
14748	:douta	=	16'h	957a;
14749	:douta	=	16'h	959a;
14750	:douta	=	16'h	9dbb;
14751	:douta	=	16'h	ae5d;
14752	:douta	=	16'h	7cf8;
14753	:douta	=	16'h	7cb7;
14754	:douta	=	16'h	63f4;
14755	:douta	=	16'h	5bf5;
14756	:douta	=	16'h	7c97;
14757	:douta	=	16'h	851a;
14758	:douta	=	16'h	7c98;
14759	:douta	=	16'h	7477;
14760	:douta	=	16'h	7cd8;
14761	:douta	=	16'h	4b74;
14762	:douta	=	16'h	4b73;
14763	:douta	=	16'h	7cd9;
14764	:douta	=	16'h	8d5a;
14765	:douta	=	16'h	857c;
14766	:douta	=	16'h	7d5b;
14767	:douta	=	16'h	6498;
14768	:douta	=	16'h	6c99;
14769	:douta	=	16'h	6437;
14770	:douta	=	16'h	6cb9;
14771	:douta	=	16'h	53d5;
14772	:douta	=	16'h	6457;
14773	:douta	=	16'h	7d1a;
14774	:douta	=	16'h	7d1a;
14775	:douta	=	16'h	7d1a;
14776	:douta	=	16'h	74b8;
14777	:douta	=	16'h	7497;
14778	:douta	=	16'h	7cb8;
14779	:douta	=	16'h	6c36;
14780	:douta	=	16'h	7497;
14781	:douta	=	16'h	7c97;
14782	:douta	=	16'h	63f4;
14783	:douta	=	16'h	63d4;
14784	:douta	=	16'h	6c35;
14785	:douta	=	16'h	63f4;
14786	:douta	=	16'h	63f4;
14787	:douta	=	16'h	7c96;
14788	:douta	=	16'h	7456;
14789	:douta	=	16'h	7496;
14790	:douta	=	16'h	7456;
14791	:douta	=	16'h	7456;
14792	:douta	=	16'h	6c56;
14793	:douta	=	16'h	7c97;
14794	:douta	=	16'h	6415;
14795	:douta	=	16'h	63f4;
14796	:douta	=	16'h	5bb3;
14797	:douta	=	16'h	7457;
14798	:douta	=	16'h	84d9;
14799	:douta	=	16'h	74d9;
14800	:douta	=	16'h	5bf6;
14801	:douta	=	16'h	5c16;
14802	:douta	=	16'h	4b74;
14803	:douta	=	16'h	6478;
14804	:douta	=	16'h	4b33;
14805	:douta	=	16'h	6498;
14806	:douta	=	16'h	6cb9;
14807	:douta	=	16'h	74fa;
14808	:douta	=	16'h	74da;
14809	:douta	=	16'h	859c;
14810	:douta	=	16'h	7d3b;
14811	:douta	=	16'h	6cba;
14812	:douta	=	16'h	853b;
14813	:douta	=	16'h	855b;
14814	:douta	=	16'h	6c98;
14815	:douta	=	16'h	74da;
14816	:douta	=	16'h	74d9;
14817	:douta	=	16'h	855b;
14818	:douta	=	16'h	7cfa;
14819	:douta	=	16'h	7d1a;
14820	:douta	=	16'h	8d5c;
14821	:douta	=	16'h	8d7c;
14822	:douta	=	16'h	855b;
14823	:douta	=	16'h	853a;
14824	:douta	=	16'h	853b;
14825	:douta	=	16'h	7d1a;
14826	:douta	=	16'h	7d3a;
14827	:douta	=	16'h	8d7b;
14828	:douta	=	16'h	95bc;
14829	:douta	=	16'h	7d3a;
14830	:douta	=	16'h	7d1a;
14831	:douta	=	16'h	855b;
14832	:douta	=	16'h	853b;
14833	:douta	=	16'h	74b8;
14834	:douta	=	16'h	7cb9;
14835	:douta	=	16'h	8d9c;
14836	:douta	=	16'h	8ddd;
14837	:douta	=	16'h	751a;
14838	:douta	=	16'h	74b9;
14839	:douta	=	16'h	2126;
14840	:douta	=	16'h	94d4;
14841	:douta	=	16'h	6370;
14842	:douta	=	16'h	bdd8;
14843	:douta	=	16'h	8c94;
14844	:douta	=	16'h	6351;
14845	:douta	=	16'h	532f;
14846	:douta	=	16'h	324d;
14847	:douta	=	16'h	6390;
14848	:douta	=	16'h	32b1;
14849	:douta	=	16'h	3af2;
14850	:douta	=	16'h	4b94;
14851	:douta	=	16'h	3b12;
14852	:douta	=	16'h	4b95;
14853	:douta	=	16'h	4b94;
14854	:douta	=	16'h	3ab0;
14855	:douta	=	16'h	5b73;
14856	:douta	=	16'h	63d4;
14857	:douta	=	16'h	6c15;
14858	:douta	=	16'h	6c35;
14859	:douta	=	16'h	73f4;
14860	:douta	=	16'h	7c76;
14861	:douta	=	16'h	6bf4;
14862	:douta	=	16'h	424b;
14863	:douta	=	16'h	6350;
14864	:douta	=	16'h	73f1;
14865	:douta	=	16'h	8432;
14866	:douta	=	16'h	9cb4;
14867	:douta	=	16'h	9cd4;
14868	:douta	=	16'h	bd96;
14869	:douta	=	16'h	7bd0;
14870	:douta	=	16'h	8410;
14871	:douta	=	16'h	a4b1;
14872	:douta	=	16'h	d615;
14873	:douta	=	16'h	ad11;
14874	:douta	=	16'h	b532;
14875	:douta	=	16'h	cdf5;
14876	:douta	=	16'h	b511;
14877	:douta	=	16'h	528b;
14878	:douta	=	16'h	6b2c;
14879	:douta	=	16'h	ad10;
14880	:douta	=	16'h	d5f5;
14881	:douta	=	16'h	bd72;
14882	:douta	=	16'h	de76;
14883	:douta	=	16'h	bdd4;
14884	:douta	=	16'h	a4d0;
14885	:douta	=	16'h	8bec;
14886	:douta	=	16'h	732a;
14887	:douta	=	16'h	7b2a;
14888	:douta	=	16'h	8b8b;
14889	:douta	=	16'h	93cb;
14890	:douta	=	16'h	8b6a;
14891	:douta	=	16'h	b48c;
14892	:douta	=	16'h	ac6c;
14893	:douta	=	16'h	ac6c;
14894	:douta	=	16'h	bccd;
14895	:douta	=	16'h	c50e;
14896	:douta	=	16'h	d5d2;
14897	:douta	=	16'h	de12;
14898	:douta	=	16'h	de33;
14899	:douta	=	16'h	e654;
14900	:douta	=	16'h	e634;
14901	:douta	=	16'h	e634;
14902	:douta	=	16'h	ddf2;
14903	:douta	=	16'h	d5b1;
14904	:douta	=	16'h	ddd1;
14905	:douta	=	16'h	d591;
14906	:douta	=	16'h	cd71;
14907	:douta	=	16'h	c50f;
14908	:douta	=	16'h	ac8f;
14909	:douta	=	16'h	8b4a;
14910	:douta	=	16'h	ac6e;
14911	:douta	=	16'h	b4cf;
14912	:douta	=	16'h	9c4d;
14913	:douta	=	16'h	9c4e;
14914	:douta	=	16'h	5acb;
14915	:douta	=	16'h	4a4a;
14916	:douta	=	16'h	8bed;
14917	:douta	=	16'h	734c;
14918	:douta	=	16'h	62eb;
14919	:douta	=	16'h	424b;
14920	:douta	=	16'h	31ea;
14921	:douta	=	16'h	2988;
14922	:douta	=	16'h	29c8;
14923	:douta	=	16'h	1947;
14924	:douta	=	16'h	31c8;
14925	:douta	=	16'h	10a4;
14926	:douta	=	16'h	10a4;
14927	:douta	=	16'h	18c4;
14928	:douta	=	16'h	10e4;
14929	:douta	=	16'h	10e4;
14930	:douta	=	16'h	10e4;
14931	:douta	=	16'h	0000;
14932	:douta	=	16'h	0042;
14933	:douta	=	16'h	0042;
14934	:douta	=	16'h	29ca;
14935	:douta	=	16'h	2168;
14936	:douta	=	16'h	10e5;
14937	:douta	=	16'h	1105;
14938	:douta	=	16'h	1906;
14939	:douta	=	16'h	5a89;
14940	:douta	=	16'h	2125;
14941	:douta	=	16'h	2146;
14942	:douta	=	16'h	39e7;
14943	:douta	=	16'h	6b2b;
14944	:douta	=	16'h	4a28;
14945	:douta	=	16'h	acf1;
14946	:douta	=	16'h	7bef;
14947	:douta	=	16'h	1969;
14948	:douta	=	16'h	29c9;
14949	:douta	=	16'h	29ec;
14950	:douta	=	16'h	00c7;
14951	:douta	=	16'h	1127;
14952	:douta	=	16'h	1127;
14953	:douta	=	16'h	3a6b;
14954	:douta	=	16'h	4a6a;
14955	:douta	=	16'h	29c9;
14956	:douta	=	16'h	73af;
14957	:douta	=	16'h	7bf0;
14958	:douta	=	16'h	428b;
14959	:douta	=	16'h	29eb;
14960	:douta	=	16'h	424b;
14961	:douta	=	16'h	31ea;
14962	:douta	=	16'h	29c9;
14963	:douta	=	16'h	1906;
14964	:douta	=	16'h	3146;
14965	:douta	=	16'h	9bed;
14966	:douta	=	16'h	8475;
14967	:douta	=	16'h	8d7a;
14968	:douta	=	16'h	8518;
14969	:douta	=	16'h	8539;
14970	:douta	=	16'h	8d59;
14971	:douta	=	16'h	8d59;
14972	:douta	=	16'h	7cd8;
14973	:douta	=	16'h	5392;
14974	:douta	=	16'h	3ab0;
14975	:douta	=	16'h	4b53;
14976	:douta	=	16'h	8519;
14977	:douta	=	16'h	8d5a;
14978	:douta	=	16'h	7456;
14979	:douta	=	16'h	9d9b;
14980	:douta	=	16'h	a5db;
14981	:douta	=	16'h	8d3a;
14982	:douta	=	16'h	7498;
14983	:douta	=	16'h	84f9;
14984	:douta	=	16'h	a5db;
14985	:douta	=	16'h	955a;
14986	:douta	=	16'h	7cb8;
14987	:douta	=	16'h	957a;
14988	:douta	=	16'h	7cd8;
14989	:douta	=	16'h	959a;
14990	:douta	=	16'h	8d7a;
14991	:douta	=	16'h	84f9;
14992	:douta	=	16'h	8d5a;
14993	:douta	=	16'h	9dbb;
14994	:douta	=	16'h	8d7a;
14995	:douta	=	16'h	7cd9;
14996	:douta	=	16'h	9d9a;
14997	:douta	=	16'h	957a;
14998	:douta	=	16'h	8d5a;
14999	:douta	=	16'h	8519;
15000	:douta	=	16'h	8539;
15001	:douta	=	16'h	955b;
15002	:douta	=	16'h	9ddc;
15003	:douta	=	16'h	a5db;
15004	:douta	=	16'h	84f9;
15005	:douta	=	16'h	84f9;
15006	:douta	=	16'h	63d5;
15007	:douta	=	16'h	7c98;
15008	:douta	=	16'h	8d7a;
15009	:douta	=	16'h	8d5a;
15010	:douta	=	16'h	7cd7;
15011	:douta	=	16'h	84f8;
15012	:douta	=	16'h	84b8;
15013	:douta	=	16'h	6c36;
15014	:douta	=	16'h	7497;
15015	:douta	=	16'h	6415;
15016	:douta	=	16'h	7cb8;
15017	:douta	=	16'h	8d5a;
15018	:douta	=	16'h	3af1;
15019	:douta	=	16'h	4b53;
15020	:douta	=	16'h	7d3b;
15021	:douta	=	16'h	74fb;
15022	:douta	=	16'h	751b;
15023	:douta	=	16'h	74d9;
15024	:douta	=	16'h	6457;
15025	:douta	=	16'h	74fa;
15026	:douta	=	16'h	5bd5;
15027	:douta	=	16'h	6416;
15028	:douta	=	16'h	3ab0;
15029	:douta	=	16'h	5373;
15030	:douta	=	16'h	7c98;
15031	:douta	=	16'h	74b8;
15032	:douta	=	16'h	6c56;
15033	:douta	=	16'h	7498;
15034	:douta	=	16'h	7497;
15035	:douta	=	16'h	7477;
15036	:douta	=	16'h	6c36;
15037	:douta	=	16'h	6c15;
15038	:douta	=	16'h	7476;
15039	:douta	=	16'h	7c97;
15040	:douta	=	16'h	63f4;
15041	:douta	=	16'h	6c14;
15042	:douta	=	16'h	6c14;
15043	:douta	=	16'h	63f4;
15044	:douta	=	16'h	7476;
15045	:douta	=	16'h	6c14;
15046	:douta	=	16'h	7477;
15047	:douta	=	16'h	7476;
15048	:douta	=	16'h	6c57;
15049	:douta	=	16'h	5bb3;
15050	:douta	=	16'h	63f5;
15051	:douta	=	16'h	6c35;
15052	:douta	=	16'h	5bd4;
15053	:douta	=	16'h	326e;
15054	:douta	=	16'h	5bd4;
15055	:douta	=	16'h	7d1b;
15056	:douta	=	16'h	6c99;
15057	:douta	=	16'h	5bf6;
15058	:douta	=	16'h	53f6;
15059	:douta	=	16'h	6499;
15060	:douta	=	16'h	4b94;
15061	:douta	=	16'h	6cb9;
15062	:douta	=	16'h	74fa;
15063	:douta	=	16'h	855b;
15064	:douta	=	16'h	855b;
15065	:douta	=	16'h	6cd9;
15066	:douta	=	16'h	8d9c;
15067	:douta	=	16'h	7d5b;
15068	:douta	=	16'h	7d1a;
15069	:douta	=	16'h	855b;
15070	:douta	=	16'h	6c98;
15071	:douta	=	16'h	853b;
15072	:douta	=	16'h	7d1a;
15073	:douta	=	16'h	74d9;
15074	:douta	=	16'h	857c;
15075	:douta	=	16'h	7d5b;
15076	:douta	=	16'h	7d1a;
15077	:douta	=	16'h	855b;
15078	:douta	=	16'h	8d7b;
15079	:douta	=	16'h	855b;
15080	:douta	=	16'h	857b;
15081	:douta	=	16'h	855b;
15082	:douta	=	16'h	8dbc;
15083	:douta	=	16'h	855b;
15084	:douta	=	16'h	857b;
15085	:douta	=	16'h	855b;
15086	:douta	=	16'h	855a;
15087	:douta	=	16'h	7d3b;
15088	:douta	=	16'h	7d3a;
15089	:douta	=	16'h	857c;
15090	:douta	=	16'h	7d1a;
15091	:douta	=	16'h	7cf9;
15092	:douta	=	16'h	74f9;
15093	:douta	=	16'h	855b;
15094	:douta	=	16'h	6c98;
15095	:douta	=	16'h	31a8;
15096	:douta	=	16'h	326d;
15097	:douta	=	16'h	6bf2;
15098	:douta	=	16'h	73f1;
15099	:douta	=	16'h	7c33;
15100	:douta	=	16'h	5b50;
15101	:douta	=	16'h	a557;
15102	:douta	=	16'h	7c33;
15103	:douta	=	16'h	42d0;
15104	:douta	=	16'h	32b0;
15105	:douta	=	16'h	4374;
15106	:douta	=	16'h	3312;
15107	:douta	=	16'h	2a90;
15108	:douta	=	16'h	222f;
15109	:douta	=	16'h	4353;
15110	:douta	=	16'h	3290;
15111	:douta	=	16'h	5352;
15112	:douta	=	16'h	63d4;
15113	:douta	=	16'h	84f8;
15114	:douta	=	16'h	63f5;
15115	:douta	=	16'h	3a4e;
15116	:douta	=	16'h	3a8e;
15117	:douta	=	16'h	6bf4;
15118	:douta	=	16'h	6350;
15119	:douta	=	16'h	7c33;
15120	:douta	=	16'h	73d2;
15121	:douta	=	16'h	8c93;
15122	:douta	=	16'h	8414;
15123	:douta	=	16'h	94d3;
15124	:douta	=	16'h	5b4f;
15125	:douta	=	16'h	7c31;
15126	:douta	=	16'h	ad55;
15127	:douta	=	16'h	bd74;
15128	:douta	=	16'h	de96;
15129	:douta	=	16'h	ad12;
15130	:douta	=	16'h	9c90;
15131	:douta	=	16'h	a4b1;
15132	:douta	=	16'h	e697;
15133	:douta	=	16'h	736d;
15134	:douta	=	16'h	7b6d;
15135	:douta	=	16'h	a4d1;
15136	:douta	=	16'h	cdf4;
15137	:douta	=	16'h	7bad;
15138	:douta	=	16'h	ce14;
15139	:douta	=	16'h	8c0e;
15140	:douta	=	16'h	838b;
15141	:douta	=	16'h	8b8c;
15142	:douta	=	16'h	7b2a;
15143	:douta	=	16'h	836a;
15144	:douta	=	16'h	93ec;
15145	:douta	=	16'h	93aa;
15146	:douta	=	16'h	8b8a;
15147	:douta	=	16'h	b4ad;
15148	:douta	=	16'h	b48b;
15149	:douta	=	16'h	bcac;
15150	:douta	=	16'h	c54f;
15151	:douta	=	16'h	cd90;
15152	:douta	=	16'h	ddf3;
15153	:douta	=	16'h	e654;
15154	:douta	=	16'h	e654;
15155	:douta	=	16'h	e654;
15156	:douta	=	16'h	de13;
15157	:douta	=	16'h	e654;
15158	:douta	=	16'h	ddf2;
15159	:douta	=	16'h	d5b1;
15160	:douta	=	16'h	cd50;
15161	:douta	=	16'h	c52f;
15162	:douta	=	16'h	bcef;
15163	:douta	=	16'h	b48e;
15164	:douta	=	16'h	8b69;
15165	:douta	=	16'h	c52f;
15166	:douta	=	16'h	c550;
15167	:douta	=	16'h	bd30;
15168	:douta	=	16'h	ac8f;
15169	:douta	=	16'h	acaf;
15170	:douta	=	16'h	734c;
15171	:douta	=	16'h	6aec;
15172	:douta	=	16'h	940e;
15173	:douta	=	16'h	83ae;
15174	:douta	=	16'h	7bae;
15175	:douta	=	16'h	422a;
15176	:douta	=	16'h	29a9;
15177	:douta	=	16'h	29a8;
15178	:douta	=	16'h	31c9;
15179	:douta	=	16'h	1926;
15180	:douta	=	16'h	10e5;
15181	:douta	=	16'h	2147;
15182	:douta	=	16'h	10c4;
15183	:douta	=	16'h	1905;
15184	:douta	=	16'h	10c4;
15185	:douta	=	16'h	10a3;
15186	:douta	=	16'h	10c3;
15187	:douta	=	16'h	10c4;
15188	:douta	=	16'h	0000;
15189	:douta	=	16'h	0000;
15190	:douta	=	16'h	0062;
15191	:douta	=	16'h	1106;
15192	:douta	=	16'h	2169;
15193	:douta	=	16'h	10a5;
15194	:douta	=	16'h	0063;
15195	:douta	=	16'h	29a7;
15196	:douta	=	16'h	0000;
15197	:douta	=	16'h	8bed;
15198	:douta	=	16'h	3186;
15199	:douta	=	16'h	734c;
15200	:douta	=	16'h	83ad;
15201	:douta	=	16'h	2966;
15202	:douta	=	16'h	630b;
15203	:douta	=	16'h	5aec;
15204	:douta	=	16'h	39e9;
15205	:douta	=	16'h	3a4b;
15206	:douta	=	16'h	4aac;
15207	:douta	=	16'h	1147;
15208	:douta	=	16'h	7bce;
15209	:douta	=	16'h	31ca;
15210	:douta	=	16'h	634e;
15211	:douta	=	16'h	426c;
15212	:douta	=	16'h	426b;
15213	:douta	=	16'h	1129;
15214	:douta	=	16'h	1128;
15215	:douta	=	16'h	0044;
15216	:douta	=	16'h	08e6;
15217	:douta	=	16'h	52ed;
15218	:douta	=	16'h	31c8;
15219	:douta	=	16'h	2167;
15220	:douta	=	16'h	a44e;
15221	:douta	=	16'h	836a;
15222	:douta	=	16'h	a5dc;
15223	:douta	=	16'h	8d39;
15224	:douta	=	16'h	8d59;
15225	:douta	=	16'h	9dba;
15226	:douta	=	16'h	957a;
15227	:douta	=	16'h	9d9a;
15228	:douta	=	16'h	9579;
15229	:douta	=	16'h	8d59;
15230	:douta	=	16'h	9dbb;
15231	:douta	=	16'h	adfc;
15232	:douta	=	16'h	6c14;
15233	:douta	=	16'h	5b93;
15234	:douta	=	16'h	53b4;
15235	:douta	=	16'h	6435;
15236	:douta	=	16'h	6cb7;
15237	:douta	=	16'h	8d7a;
15238	:douta	=	16'h	ae1c;
15239	:douta	=	16'h	957a;
15240	:douta	=	16'h	9d7a;
15241	:douta	=	16'h	8d3a;
15242	:douta	=	16'h	959b;
15243	:douta	=	16'h	957b;
15244	:douta	=	16'h	8d5a;
15245	:douta	=	16'h	853a;
15246	:douta	=	16'h	95bb;
15247	:douta	=	16'h	8d5a;
15248	:douta	=	16'h	955b;
15249	:douta	=	16'h	8d1a;
15250	:douta	=	16'h	957a;
15251	:douta	=	16'h	959b;
15252	:douta	=	16'h	74b8;
15253	:douta	=	16'h	8d3a;
15254	:douta	=	16'h	955a;
15255	:douta	=	16'h	7cd9;
15256	:douta	=	16'h	84f9;
15257	:douta	=	16'h	9dbb;
15258	:douta	=	16'h	8d5a;
15259	:douta	=	16'h	6c77;
15260	:douta	=	16'h	955a;
15261	:douta	=	16'h	957a;
15262	:douta	=	16'h	9ddb;
15263	:douta	=	16'h	be9e;
15264	:douta	=	16'h	7c76;
15265	:douta	=	16'h	5331;
15266	:douta	=	16'h	6c36;
15267	:douta	=	16'h	6c56;
15268	:douta	=	16'h	5bd5;
15269	:douta	=	16'h	6c56;
15270	:douta	=	16'h	6c76;
15271	:douta	=	16'h	6436;
15272	:douta	=	16'h	5393;
15273	:douta	=	16'h	5373;
15274	:douta	=	16'h	5394;
15275	:douta	=	16'h	6416;
15276	:douta	=	16'h	4b32;
15277	:douta	=	16'h	328f;
15278	:douta	=	16'h	42d0;
15279	:douta	=	16'h	6cb9;
15280	:douta	=	16'h	753b;
15281	:douta	=	16'h	5bd6;
15282	:douta	=	16'h	6458;
15283	:douta	=	16'h	6457;
15284	:douta	=	16'h	855b;
15285	:douta	=	16'h	6416;
15286	:douta	=	16'h	5393;
15287	:douta	=	16'h	4b53;
15288	:douta	=	16'h	5bd4;
15289	:douta	=	16'h	7cd8;
15290	:douta	=	16'h	7cd9;
15291	:douta	=	16'h	7497;
15292	:douta	=	16'h	7477;
15293	:douta	=	16'h	7436;
15294	:douta	=	16'h	84d8;
15295	:douta	=	16'h	7c77;
15296	:douta	=	16'h	63f5;
15297	:douta	=	16'h	7c97;
15298	:douta	=	16'h	7c97;
15299	:douta	=	16'h	7c96;
15300	:douta	=	16'h	84b7;
15301	:douta	=	16'h	7457;
15302	:douta	=	16'h	6bf4;
15303	:douta	=	16'h	6c35;
15304	:douta	=	16'h	7434;
15305	:douta	=	16'h	7455;
15306	:douta	=	16'h	5bf5;
15307	:douta	=	16'h	5373;
15308	:douta	=	16'h	4b93;
15309	:douta	=	16'h	4311;
15310	:douta	=	16'h	3a90;
15311	:douta	=	16'h	3b13;
15312	:douta	=	16'h	5c78;
15313	:douta	=	16'h	6cb9;
15314	:douta	=	16'h	5c38;
15315	:douta	=	16'h	5c58;
15316	:douta	=	16'h	751b;
15317	:douta	=	16'h	6c99;
15318	:douta	=	16'h	6458;
15319	:douta	=	16'h	6458;
15320	:douta	=	16'h	6478;
15321	:douta	=	16'h	74da;
15322	:douta	=	16'h	74fa;
15323	:douta	=	16'h	74da;
15324	:douta	=	16'h	7d1a;
15325	:douta	=	16'h	857c;
15326	:douta	=	16'h	855b;
15327	:douta	=	16'h	74d9;
15328	:douta	=	16'h	74fa;
15329	:douta	=	16'h	7d3a;
15330	:douta	=	16'h	7cfa;
15331	:douta	=	16'h	7d3a;
15332	:douta	=	16'h	7d3a;
15333	:douta	=	16'h	74fa;
15334	:douta	=	16'h	7d1a;
15335	:douta	=	16'h	7d3b;
15336	:douta	=	16'h	7d3a;
15337	:douta	=	16'h	8d9c;
15338	:douta	=	16'h	7d3a;
15339	:douta	=	16'h	7499;
15340	:douta	=	16'h	7cfa;
15341	:douta	=	16'h	8d9c;
15342	:douta	=	16'h	6cb9;
15343	:douta	=	16'h	7cd9;
15344	:douta	=	16'h	853b;
15345	:douta	=	16'h	8d7b;
15346	:douta	=	16'h	7d1a;
15347	:douta	=	16'h	7d1a;
15348	:douta	=	16'h	7d3b;
15349	:douta	=	16'h	6417;
15350	:douta	=	16'h	5bf5;
15351	:douta	=	16'h	1906;
15352	:douta	=	16'h	9d35;
15353	:douta	=	16'h	7c13;
15354	:douta	=	16'h	9518;
15355	:douta	=	16'h	63d3;
15356	:douta	=	16'h	8cf6;
15357	:douta	=	16'h	42cf;
15358	:douta	=	16'h	5b50;
15359	:douta	=	16'h	6bb1;
15360	:douta	=	16'h	4353;
15361	:douta	=	16'h	32d1;
15362	:douta	=	16'h	3b53;
15363	:douta	=	16'h	3291;
15364	:douta	=	16'h	3b12;
15365	:douta	=	16'h	4354;
15366	:douta	=	16'h	5bd4;
15367	:douta	=	16'h	5b93;
15368	:douta	=	16'h	5bb4;
15369	:douta	=	16'h	5392;
15370	:douta	=	16'h	5372;
15371	:douta	=	16'h	6392;
15372	:douta	=	16'h	6bf3;
15373	:douta	=	16'h	84b7;
15374	:douta	=	16'h	6370;
15375	:douta	=	16'h	7412;
15376	:douta	=	16'h	6bb1;
15377	:douta	=	16'h	94d4;
15378	:douta	=	16'h	634f;
15379	:douta	=	16'h	c5f7;
15380	:douta	=	16'h	a515;
15381	:douta	=	16'h	9d15;
15382	:douta	=	16'h	7390;
15383	:douta	=	16'h	b553;
15384	:douta	=	16'h	c5b4;
15385	:douta	=	16'h	a4f1;
15386	:douta	=	16'h	cdf4;
15387	:douta	=	16'h	c5d5;
15388	:douta	=	16'h	de76;
15389	:douta	=	16'h	734c;
15390	:douta	=	16'h	6aea;
15391	:douta	=	16'h	738c;
15392	:douta	=	16'h	acd1;
15393	:douta	=	16'h	9c8f;
15394	:douta	=	16'h	f77a;
15395	:douta	=	16'h	bd94;
15396	:douta	=	16'h	838a;
15397	:douta	=	16'h	8bac;
15398	:douta	=	16'h	8b6a;
15399	:douta	=	16'h	8b6a;
15400	:douta	=	16'h	93cb;
15401	:douta	=	16'h	9beb;
15402	:douta	=	16'h	93cb;
15403	:douta	=	16'h	b4ac;
15404	:douta	=	16'h	b4ac;
15405	:douta	=	16'h	c50e;
15406	:douta	=	16'h	cd6f;
15407	:douta	=	16'h	d5b1;
15408	:douta	=	16'h	e613;
15409	:douta	=	16'h	e655;
15410	:douta	=	16'h	e655;
15411	:douta	=	16'h	e654;
15412	:douta	=	16'h	ddf2;
15413	:douta	=	16'h	e633;
15414	:douta	=	16'h	ddf2;
15415	:douta	=	16'h	cd90;
15416	:douta	=	16'h	bcee;
15417	:douta	=	16'h	bcef;
15418	:douta	=	16'h	b48e;
15419	:douta	=	16'h	9bcb;
15420	:douta	=	16'h	8348;
15421	:douta	=	16'h	ac6d;
15422	:douta	=	16'h	ac8e;
15423	:douta	=	16'h	bd10;
15424	:douta	=	16'h	acaf;
15425	:douta	=	16'h	acaf;
15426	:douta	=	16'h	83cd;
15427	:douta	=	16'h	7b4c;
15428	:douta	=	16'h	9c4f;
15429	:douta	=	16'h	83ae;
15430	:douta	=	16'h	8bee;
15431	:douta	=	16'h	3a0a;
15432	:douta	=	16'h	2168;
15433	:douta	=	16'h	4229;
15434	:douta	=	16'h	31a9;
15435	:douta	=	16'h	2168;
15436	:douta	=	16'h	1905;
15437	:douta	=	16'h	1084;
15438	:douta	=	16'h	2966;
15439	:douta	=	16'h	18e5;
15440	:douta	=	16'h	18e5;
15441	:douta	=	16'h	10c3;
15442	:douta	=	16'h	10c4;
15443	:douta	=	16'h	1905;
15444	:douta	=	16'h	10c4;
15445	:douta	=	16'h	0042;
15446	:douta	=	16'h	0000;
15447	:douta	=	16'h	0062;
15448	:douta	=	16'h	21ca;
15449	:douta	=	16'h	1989;
15450	:douta	=	16'h	424a;
15451	:douta	=	16'h	2987;
15452	:douta	=	16'h	39c6;
15453	:douta	=	16'h	08c3;
15454	:douta	=	16'h	0883;
15455	:douta	=	16'h	5aaa;
15456	:douta	=	16'h	83cd;
15457	:douta	=	16'h	7bcd;
15458	:douta	=	16'h	736d;
15459	:douta	=	16'h	2967;
15460	:douta	=	16'h	83ce;
15461	:douta	=	16'h	29ca;
15462	:douta	=	16'h	1128;
15463	:douta	=	16'h	0064;
15464	:douta	=	16'h	29ca;
15465	:douta	=	16'h	08c5;
15466	:douta	=	16'h	320a;
15467	:douta	=	16'h	31c9;
15468	:douta	=	16'h	a4f1;
15469	:douta	=	16'h	4aad;
15470	:douta	=	16'h	73d0;
15471	:douta	=	16'h	426b;
15472	:douta	=	16'h	4a8b;
15473	:douta	=	16'h	3a2c;
15474	:douta	=	16'h	1968;
15475	:douta	=	16'h	08a5;
15476	:douta	=	16'h	6289;
15477	:douta	=	16'h	838c;
15478	:douta	=	16'h	9d9a;
15479	:douta	=	16'h	8d19;
15480	:douta	=	16'h	8d59;
15481	:douta	=	16'h	84f8;
15482	:douta	=	16'h	9559;
15483	:douta	=	16'h	9dba;
15484	:douta	=	16'h	a59a;
15485	:douta	=	16'h	9579;
15486	:douta	=	16'h	957a;
15487	:douta	=	16'h	9d9a;
15488	:douta	=	16'h	ae1c;
15489	:douta	=	16'h	a5fb;
15490	:douta	=	16'h	7476;
15491	:douta	=	16'h	5394;
15492	:douta	=	16'h	4b53;
15493	:douta	=	16'h	84d8;
15494	:douta	=	16'h	9dbb;
15495	:douta	=	16'h	959b;
15496	:douta	=	16'h	a5db;
15497	:douta	=	16'h	9d9b;
15498	:douta	=	16'h	959a;
15499	:douta	=	16'h	8d5a;
15500	:douta	=	16'h	9ddb;
15501	:douta	=	16'h	84f9;
15502	:douta	=	16'h	8d3a;
15503	:douta	=	16'h	9ddc;
15504	:douta	=	16'h	9ddc;
15505	:douta	=	16'h	9dbc;
15506	:douta	=	16'h	957b;
15507	:douta	=	16'h	957a;
15508	:douta	=	16'h	957a;
15509	:douta	=	16'h	8d5a;
15510	:douta	=	16'h	7cb8;
15511	:douta	=	16'h	7cf8;
15512	:douta	=	16'h	74b8;
15513	:douta	=	16'h	8519;
15514	:douta	=	16'h	8519;
15515	:douta	=	16'h	8d5a;
15516	:douta	=	16'h	959b;
15517	:douta	=	16'h	84d7;
15518	:douta	=	16'h	53b4;
15519	:douta	=	16'h	6c77;
15520	:douta	=	16'h	bebe;
15521	:douta	=	16'h	84b5;
15522	:douta	=	16'h	52ce;
15523	:douta	=	16'h	324c;
15524	:douta	=	16'h	21cb;
15525	:douta	=	16'h	4bb6;
15526	:douta	=	16'h	4bd4;
15527	:douta	=	16'h	4353;
15528	:douta	=	16'h	4b74;
15529	:douta	=	16'h	53d5;
15530	:douta	=	16'h	4b53;
15531	:douta	=	16'h	3af2;
15532	:douta	=	16'h	5373;
15533	:douta	=	16'h	5bb3;
15534	:douta	=	16'h	63d4;
15535	:douta	=	16'h	42b0;
15536	:douta	=	16'h	5b93;
15537	:douta	=	16'h	6c36;
15538	:douta	=	16'h	53d4;
15539	:douta	=	16'h	42f2;
15540	:douta	=	16'h	6c78;
15541	:douta	=	16'h	7498;
15542	:douta	=	16'h	6416;
15543	:douta	=	16'h	6416;
15544	:douta	=	16'h	5bd4;
15545	:douta	=	16'h	6415;
15546	:douta	=	16'h	7cf9;
15547	:douta	=	16'h	7d3a;
15548	:douta	=	16'h	8d5b;
15549	:douta	=	16'h	84d9;
15550	:douta	=	16'h	7497;
15551	:douta	=	16'h	7c97;
15552	:douta	=	16'h	7c97;
15553	:douta	=	16'h	7c97;
15554	:douta	=	16'h	84f8;
15555	:douta	=	16'h	7455;
15556	:douta	=	16'h	7434;
15557	:douta	=	16'h	7455;
15558	:douta	=	16'h	6bd3;
15559	:douta	=	16'h	73f4;
15560	:douta	=	16'h	4acd;
15561	:douta	=	16'h	324b;
15562	:douta	=	16'h	3aaf;
15563	:douta	=	16'h	4373;
15564	:douta	=	16'h	4bd6;
15565	:douta	=	16'h	5417;
15566	:douta	=	16'h	4bd5;
15567	:douta	=	16'h	4395;
15568	:douta	=	16'h	5c58;
15569	:douta	=	16'h	6458;
15570	:douta	=	16'h	6cb9;
15571	:douta	=	16'h	6478;
15572	:douta	=	16'h	5c58;
15573	:douta	=	16'h	74fb;
15574	:douta	=	16'h	751a;
15575	:douta	=	16'h	4395;
15576	:douta	=	16'h	5c16;
15577	:douta	=	16'h	6cba;
15578	:douta	=	16'h	74b9;
15579	:douta	=	16'h	7cfa;
15580	:douta	=	16'h	857b;
15581	:douta	=	16'h	74f9;
15582	:douta	=	16'h	857b;
15583	:douta	=	16'h	8d7c;
15584	:douta	=	16'h	7d3a;
15585	:douta	=	16'h	74fa;
15586	:douta	=	16'h	7d3a;
15587	:douta	=	16'h	857c;
15588	:douta	=	16'h	7d1a;
15589	:douta	=	16'h	6cb9;
15590	:douta	=	16'h	855b;
15591	:douta	=	16'h	855b;
15592	:douta	=	16'h	7d3a;
15593	:douta	=	16'h	7d3a;
15594	:douta	=	16'h	857b;
15595	:douta	=	16'h	7d3b;
15596	:douta	=	16'h	7cfa;
15597	:douta	=	16'h	7d3a;
15598	:douta	=	16'h	855b;
15599	:douta	=	16'h	6457;
15600	:douta	=	16'h	7cfa;
15601	:douta	=	16'h	855b;
15602	:douta	=	16'h	8d9c;
15603	:douta	=	16'h	7cf9;
15604	:douta	=	16'h	7d1a;
15605	:douta	=	16'h	7d1a;
15606	:douta	=	16'h	7cd9;
15607	:douta	=	16'h	2126;
15608	:douta	=	16'h	42ef;
15609	:douta	=	16'h	324d;
15610	:douta	=	16'h	4b30;
15611	:douta	=	16'h	6bb1;
15612	:douta	=	16'h	7c33;
15613	:douta	=	16'h	9517;
15614	:douta	=	16'h	42ce;
15615	:douta	=	16'h	5b71;
15616	:douta	=	16'h	32b1;
15617	:douta	=	16'h	4353;
15618	:douta	=	16'h	32d2;
15619	:douta	=	16'h	4bd6;
15620	:douta	=	16'h	2a6f;
15621	:douta	=	16'h	32d2;
15622	:douta	=	16'h	4b93;
15623	:douta	=	16'h	326e;
15624	:douta	=	16'h	5352;
15625	:douta	=	16'h	7456;
15626	:douta	=	16'h	7456;
15627	:douta	=	16'h	5330;
15628	:douta	=	16'h	42ce;
15629	:douta	=	16'h	7414;
15630	:douta	=	16'h	52cf;
15631	:douta	=	16'h	7c32;
15632	:douta	=	16'h	6bd2;
15633	:douta	=	16'h	a516;
15634	:douta	=	16'h	9495;
15635	:douta	=	16'h	8c93;
15636	:douta	=	16'h	9cb4;
15637	:douta	=	16'h	6bb0;
15638	:douta	=	16'h	7bd0;
15639	:douta	=	16'h	8c51;
15640	:douta	=	16'h	ce15;
15641	:douta	=	16'h	ce36;
15642	:douta	=	16'h	cdf6;
15643	:douta	=	16'h	d678;
15644	:douta	=	16'h	b554;
15645	:douta	=	16'h	a4b2;
15646	:douta	=	16'h	83cf;
15647	:douta	=	16'h	ad12;
15648	:douta	=	16'h	ad12;
15649	:douta	=	16'h	c5d4;
15650	:douta	=	16'h	836b;
15651	:douta	=	16'h	6aa9;
15652	:douta	=	16'h	8bab;
15653	:douta	=	16'h	9beb;
15654	:douta	=	16'h	93ab;
15655	:douta	=	16'h	93ec;
15656	:douta	=	16'h	93ab;
15657	:douta	=	16'h	b48c;
15658	:douta	=	16'h	ac4c;
15659	:douta	=	16'h	b4ad;
15660	:douta	=	16'h	c52e;
15661	:douta	=	16'h	cd2f;
15662	:douta	=	16'h	ddf2;
15663	:douta	=	16'h	e634;
15664	:douta	=	16'h	e676;
15665	:douta	=	16'h	e633;
15666	:douta	=	16'h	de34;
15667	:douta	=	16'h	ddd2;
15668	:douta	=	16'h	ddf2;
15669	:douta	=	16'h	c50f;
15670	:douta	=	16'h	ddd2;
15671	:douta	=	16'h	d590;
15672	:douta	=	16'h	b46d;
15673	:douta	=	16'h	b48e;
15674	:douta	=	16'h	9beb;
15675	:douta	=	16'h	9beb;
15676	:douta	=	16'h	a40c;
15677	:douta	=	16'h	b48e;
15678	:douta	=	16'h	bd0f;
15679	:douta	=	16'h	cd71;
15680	:douta	=	16'h	bcf0;
15681	:douta	=	16'h	b4cf;
15682	:douta	=	16'h	9c6e;
15683	:douta	=	16'h	940e;
15684	:douta	=	16'h	a46f;
15685	:douta	=	16'h	8bef;
15686	:douta	=	16'h	83ce;
15687	:douta	=	16'h	4a8b;
15688	:douta	=	16'h	424a;
15689	:douta	=	16'h	4a4a;
15690	:douta	=	16'h	3a0a;
15691	:douta	=	16'h	29ca;
15692	:douta	=	16'h	1947;
15693	:douta	=	16'h	2168;
15694	:douta	=	16'h	0883;
15695	:douta	=	16'h	422a;
15696	:douta	=	16'h	10a4;
15697	:douta	=	16'h	18e5;
15698	:douta	=	16'h	18c4;
15699	:douta	=	16'h	10e4;
15700	:douta	=	16'h	10c5;
15701	:douta	=	16'h	10a4;
15702	:douta	=	16'h	2126;
15703	:douta	=	16'h	10e5;
15704	:douta	=	16'h	0000;
15705	:douta	=	16'h	0000;
15706	:douta	=	16'h	52ee;
15707	:douta	=	16'h	4ace;
15708	:douta	=	16'h	424b;
15709	:douta	=	16'h	4a28;
15710	:douta	=	16'h	942e;
15711	:douta	=	16'h	39e8;
15712	:douta	=	16'h	8c2e;
15713	:douta	=	16'h	732c;
15714	:douta	=	16'h	2166;
15715	:douta	=	16'h	1063;
15716	:douta	=	16'h	3207;
15717	:douta	=	16'h	1105;
15718	:douta	=	16'h	4249;
15719	:douta	=	16'h	52aa;
15720	:douta	=	16'h	738d;
15721	:douta	=	16'h	9470;
15722	:douta	=	16'h	31ea;
15723	:douta	=	16'h	6b4d;
15724	:douta	=	16'h	116a;
15725	:douta	=	16'h	1128;
15726	:douta	=	16'h	00a5;
15727	:douta	=	16'h	320b;
15728	:douta	=	16'h	3a6b;
15729	:douta	=	16'h	52cc;
15730	:douta	=	16'h	4aac;
15731	:douta	=	16'h	2169;
15732	:douta	=	16'h	acaf;
15733	:douta	=	16'h	62ca;
15734	:douta	=	16'h	adfb;
15735	:douta	=	16'h	9d9a;
15736	:douta	=	16'h	957a;
15737	:douta	=	16'h	8d18;
15738	:douta	=	16'h	84f8;
15739	:douta	=	16'h	9d9a;
15740	:douta	=	16'h	9559;
15741	:douta	=	16'h	957a;
15742	:douta	=	16'h	9579;
15743	:douta	=	16'h	9559;
15744	:douta	=	16'h	8d39;
15745	:douta	=	16'h	9d9a;
15746	:douta	=	16'h	957a;
15747	:douta	=	16'h	9d9a;
15748	:douta	=	16'h	9dda;
15749	:douta	=	16'h	a5fb;
15750	:douta	=	16'h	8518;
15751	:douta	=	16'h	5bf6;
15752	:douta	=	16'h	7c97;
15753	:douta	=	16'h	8519;
15754	:douta	=	16'h	853a;
15755	:douta	=	16'h	7cd9;
15756	:douta	=	16'h	9ddb;
15757	:douta	=	16'h	957b;
15758	:douta	=	16'h	a5db;
15759	:douta	=	16'h	a5dc;
15760	:douta	=	16'h	959b;
15761	:douta	=	16'h	957b;
15762	:douta	=	16'h	8d5a;
15763	:douta	=	16'h	9dbc;
15764	:douta	=	16'h	851a;
15765	:douta	=	16'h	6457;
15766	:douta	=	16'h	9dbb;
15767	:douta	=	16'h	8d3a;
15768	:douta	=	16'h	8d3a;
15769	:douta	=	16'h	7497;
15770	:douta	=	16'h	8519;
15771	:douta	=	16'h	b65d;
15772	:douta	=	16'h	84d8;
15773	:douta	=	16'h	7477;
15774	:douta	=	16'h	8d19;
15775	:douta	=	16'h	8d59;
15776	:douta	=	16'h	7cb8;
15777	:douta	=	16'h	940f;
15778	:douta	=	16'h	7b4b;
15779	:douta	=	16'h	10e5;
15780	:douta	=	16'h	1905;
15781	:douta	=	16'h	1948;
15782	:douta	=	16'h	2af3;
15783	:douta	=	16'h	4bf6;
15784	:douta	=	16'h	3b33;
15785	:douta	=	16'h	4374;
15786	:douta	=	16'h	5bd5;
15787	:douta	=	16'h	5bf5;
15788	:douta	=	16'h	4312;
15789	:douta	=	16'h	5bd4;
15790	:douta	=	16'h	6c35;
15791	:douta	=	16'h	5bb3;
15792	:douta	=	16'h	5331;
15793	:douta	=	16'h	328e;
15794	:douta	=	16'h	5b93;
15795	:douta	=	16'h	7436;
15796	:douta	=	16'h	5bd4;
15797	:douta	=	16'h	6c97;
15798	:douta	=	16'h	5bd5;
15799	:douta	=	16'h	6c98;
15800	:douta	=	16'h	5c16;
15801	:douta	=	16'h	5c16;
15802	:douta	=	16'h	5bf6;
15803	:douta	=	16'h	6436;
15804	:douta	=	16'h	5bf5;
15805	:douta	=	16'h	5bb4;
15806	:douta	=	16'h	8d3a;
15807	:douta	=	16'h	955a;
15808	:douta	=	16'h	7cb7;
15809	:douta	=	16'h	7435;
15810	:douta	=	16'h	7455;
15811	:douta	=	16'h	6c14;
15812	:douta	=	16'h	6c35;
15813	:douta	=	16'h	7c75;
15814	:douta	=	16'h	73f2;
15815	:douta	=	16'h	4a6a;
15816	:douta	=	16'h	2106;
15817	:douta	=	16'h	2125;
15818	:douta	=	16'h	18c4;
15819	:douta	=	16'h	1a4f;
15820	:douta	=	16'h	3376;
15821	:douta	=	16'h	3b75;
15822	:douta	=	16'h	4395;
15823	:douta	=	16'h	4395;
15824	:douta	=	16'h	53f6;
15825	:douta	=	16'h	5c58;
15826	:douta	=	16'h	3b55;
15827	:douta	=	16'h	4395;
15828	:douta	=	16'h	5c38;
15829	:douta	=	16'h	6cba;
15830	:douta	=	16'h	751b;
15831	:douta	=	16'h	7d3b;
15832	:douta	=	16'h	857c;
15833	:douta	=	16'h	6c99;
15834	:douta	=	16'h	6c78;
15835	:douta	=	16'h	74fa;
15836	:douta	=	16'h	6437;
15837	:douta	=	16'h	5bf7;
15838	:douta	=	16'h	855b;
15839	:douta	=	16'h	7d1a;
15840	:douta	=	16'h	855b;
15841	:douta	=	16'h	7d3a;
15842	:douta	=	16'h	857b;
15843	:douta	=	16'h	7cfa;
15844	:douta	=	16'h	855b;
15845	:douta	=	16'h	857c;
15846	:douta	=	16'h	855b;
15847	:douta	=	16'h	7d1a;
15848	:douta	=	16'h	855b;
15849	:douta	=	16'h	855c;
15850	:douta	=	16'h	7d1a;
15851	:douta	=	16'h	7499;
15852	:douta	=	16'h	7cfa;
15853	:douta	=	16'h	8d7b;
15854	:douta	=	16'h	74fa;
15855	:douta	=	16'h	855b;
15856	:douta	=	16'h	855b;
15857	:douta	=	16'h	8d7b;
15858	:douta	=	16'h	7cd9;
15859	:douta	=	16'h	6478;
15860	:douta	=	16'h	7cf9;
15861	:douta	=	16'h	857b;
15862	:douta	=	16'h	74b9;
15863	:douta	=	16'h	1906;
15864	:douta	=	16'h	bdf9;
15865	:douta	=	16'h	84b6;
15866	:douta	=	16'h	b597;
15867	:douta	=	16'h	6bb1;
15868	:douta	=	16'h	6391;
15869	:douta	=	16'h	1149;
15870	:douta	=	16'h	5b71;
15871	:douta	=	16'h	7c74;
15872	:douta	=	16'h	32d1;
15873	:douta	=	16'h	32f2;
15874	:douta	=	16'h	3b53;
15875	:douta	=	16'h	4374;
15876	:douta	=	16'h	222f;
15877	:douta	=	16'h	3b12;
15878	:douta	=	16'h	6436;
15879	:douta	=	16'h	63f4;
15880	:douta	=	16'h	7456;
15881	:douta	=	16'h	4b31;
15882	:douta	=	16'h	42d0;
15883	:douta	=	16'h	6bd3;
15884	:douta	=	16'h	52f0;
15885	:douta	=	16'h	8cd7;
15886	:douta	=	16'h	6371;
15887	:douta	=	16'h	73f2;
15888	:douta	=	16'h	6391;
15889	:douta	=	16'h	8433;
15890	:douta	=	16'h	632f;
15891	:douta	=	16'h	a515;
15892	:douta	=	16'h	d638;
15893	:douta	=	16'h	94b3;
15894	:douta	=	16'h	8411;
15895	:douta	=	16'h	9c91;
15896	:douta	=	16'h	a4b1;
15897	:douta	=	16'h	73ef;
15898	:douta	=	16'h	bd94;
15899	:douta	=	16'h	d657;
15900	:douta	=	16'h	942f;
15901	:douta	=	16'h	bdb5;
15902	:douta	=	16'h	a4d3;
15903	:douta	=	16'h	b595;
15904	:douta	=	16'h	8bee;
15905	:douta	=	16'h	a511;
15906	:douta	=	16'h	7b2a;
15907	:douta	=	16'h	7b4a;
15908	:douta	=	16'h	93cb;
15909	:douta	=	16'h	a44c;
15910	:douta	=	16'h	8b6a;
15911	:douta	=	16'h	a42c;
15912	:douta	=	16'h	9beb;
15913	:douta	=	16'h	b44d;
15914	:douta	=	16'h	a40c;
15915	:douta	=	16'h	bcad;
15916	:douta	=	16'h	cd6f;
15917	:douta	=	16'h	cd70;
15918	:douta	=	16'h	ddf3;
15919	:douta	=	16'h	ee75;
15920	:douta	=	16'h	e655;
15921	:douta	=	16'h	de34;
15922	:douta	=	16'h	ddf2;
15923	:douta	=	16'h	e613;
15924	:douta	=	16'h	d571;
15925	:douta	=	16'h	bcae;
15926	:douta	=	16'h	d591;
15927	:douta	=	16'h	cd6f;
15928	:douta	=	16'h	a42d;
15929	:douta	=	16'h	9c0c;
15930	:douta	=	16'h	8308;
15931	:douta	=	16'h	b4ce;
15932	:douta	=	16'h	a40c;
15933	:douta	=	16'h	bcee;
15934	:douta	=	16'h	cd91;
15935	:douta	=	16'h	cdb2;
15936	:douta	=	16'h	c530;
15937	:douta	=	16'h	bcef;
15938	:douta	=	16'h	ac8f;
15939	:douta	=	16'h	9c4e;
15940	:douta	=	16'h	a48f;
15941	:douta	=	16'h	8c2f;
15942	:douta	=	16'h	8bef;
15943	:douta	=	16'h	52ac;
15944	:douta	=	16'h	5acc;
15945	:douta	=	16'h	52ac;
15946	:douta	=	16'h	424b;
15947	:douta	=	16'h	31ea;
15948	:douta	=	16'h	2188;
15949	:douta	=	16'h	2168;
15950	:douta	=	16'h	10e6;
15951	:douta	=	16'h	422a;
15952	:douta	=	16'h	4a4a;
15953	:douta	=	16'h	1084;
15954	:douta	=	16'h	10e4;
15955	:douta	=	16'h	10c4;
15956	:douta	=	16'h	10e5;
15957	:douta	=	16'h	10c4;
15958	:douta	=	16'h	10e5;
15959	:douta	=	16'h	2968;
15960	:douta	=	16'h	0000;
15961	:douta	=	16'h	0000;
15962	:douta	=	16'h	1107;
15963	:douta	=	16'h	5b0e;
15964	:douta	=	16'h	5b2f;
15965	:douta	=	16'h	4208;
15966	:douta	=	16'h	4a49;
15967	:douta	=	16'h	31a7;
15968	:douta	=	16'h	5269;
15969	:douta	=	16'h	6b2b;
15970	:douta	=	16'h	4a89;
15971	:douta	=	16'h	3966;
15972	:douta	=	16'h	7bcc;
15973	:douta	=	16'h	4a8a;
15974	:douta	=	16'h	29a9;
15975	:douta	=	16'h	29a9;
15976	:douta	=	16'h	10e6;
15977	:douta	=	16'h	738e;
15978	:douta	=	16'h	08e6;
15979	:douta	=	16'h	3a2a;
15980	:douta	=	16'h	5b0d;
15981	:douta	=	16'h	5b0d;
15982	:douta	=	16'h	21aa;
15983	:douta	=	16'h	4a8c;
15984	:douta	=	16'h	2a0c;
15985	:douta	=	16'h	2169;
15986	:douta	=	16'h	1148;
15987	:douta	=	16'h	0044;
15988	:douta	=	16'h	838c;
15989	:douta	=	16'h	6aca;
15990	:douta	=	16'h	9d79;
15991	:douta	=	16'h	8d18;
15992	:douta	=	16'h	8d39;
15993	:douta	=	16'h	8d59;
15994	:douta	=	16'h	959a;
15995	:douta	=	16'h	7cb7;
15996	:douta	=	16'h	8d39;
15997	:douta	=	16'h	9d9a;
15998	:douta	=	16'h	9559;
15999	:douta	=	16'h	9ddb;
16000	:douta	=	16'h	84f8;
16001	:douta	=	16'h	8d18;
16002	:douta	=	16'h	9579;
16003	:douta	=	16'h	9d9a;
16004	:douta	=	16'h	9559;
16005	:douta	=	16'h	9d9a;
16006	:douta	=	16'h	a5fb;
16007	:douta	=	16'h	a5db;
16008	:douta	=	16'h	7c76;
16009	:douta	=	16'h	7476;
16010	:douta	=	16'h	6416;
16011	:douta	=	16'h	7cd8;
16012	:douta	=	16'h	8519;
16013	:douta	=	16'h	a5db;
16014	:douta	=	16'h	957a;
16015	:douta	=	16'h	955a;
16016	:douta	=	16'h	9dbb;
16017	:douta	=	16'h	a5fc;
16018	:douta	=	16'h	8d5a;
16019	:douta	=	16'h	7cf9;
16020	:douta	=	16'h	959b;
16021	:douta	=	16'h	8519;
16022	:douta	=	16'h	8d5b;
16023	:douta	=	16'h	ae1b;
16024	:douta	=	16'h	ae1c;
16025	:douta	=	16'h	8d39;
16026	:douta	=	16'h	7cb8;
16027	:douta	=	16'h	8d39;
16028	:douta	=	16'h	b67d;
16029	:douta	=	16'h	9d9a;
16030	:douta	=	16'h	8497;
16031	:douta	=	16'h	7cb7;
16032	:douta	=	16'h	84d8;
16033	:douta	=	16'h	9471;
16034	:douta	=	16'h	834b;
16035	:douta	=	16'h	1105;
16036	:douta	=	16'h	18e5;
16037	:douta	=	16'h	1148;
16038	:douta	=	16'h	5373;
16039	:douta	=	16'h	53d5;
16040	:douta	=	16'h	5bf5;
16041	:douta	=	16'h	5c37;
16042	:douta	=	16'h	5bf5;
16043	:douta	=	16'h	6457;
16044	:douta	=	16'h	63f5;
16045	:douta	=	16'h	4b52;
16046	:douta	=	16'h	5b93;
16047	:douta	=	16'h	5b93;
16048	:douta	=	16'h	6bf5;
16049	:douta	=	16'h	42f0;
16050	:douta	=	16'h	42cf;
16051	:douta	=	16'h	63b3;
16052	:douta	=	16'h	5352;
16053	:douta	=	16'h	42f0;
16054	:douta	=	16'h	7d1a;
16055	:douta	=	16'h	5c37;
16056	:douta	=	16'h	6457;
16057	:douta	=	16'h	6437;
16058	:douta	=	16'h	5c16;
16059	:douta	=	16'h	6437;
16060	:douta	=	16'h	6436;
16061	:douta	=	16'h	6415;
16062	:douta	=	16'h	63f5;
16063	:douta	=	16'h	7cb7;
16064	:douta	=	16'h	84d7;
16065	:douta	=	16'h	7cb7;
16066	:douta	=	16'h	6c35;
16067	:douta	=	16'h	6c14;
16068	:douta	=	16'h	7413;
16069	:douta	=	16'h	7435;
16070	:douta	=	16'h	73f1;
16071	:douta	=	16'h	4208;
16072	:douta	=	16'h	2126;
16073	:douta	=	16'h	1905;
16074	:douta	=	16'h	10e5;
16075	:douta	=	16'h	3b34;
16076	:douta	=	16'h	4bb6;
16077	:douta	=	16'h	4396;
16078	:douta	=	16'h	4bd6;
16079	:douta	=	16'h	53f7;
16080	:douta	=	16'h	4bf6;
16081	:douta	=	16'h	5c78;
16082	:douta	=	16'h	6479;
16083	:douta	=	16'h	5c78;
16084	:douta	=	16'h	3b33;
16085	:douta	=	16'h	5c17;
16086	:douta	=	16'h	6458;
16087	:douta	=	16'h	74fa;
16088	:douta	=	16'h	7d5b;
16089	:douta	=	16'h	6478;
16090	:douta	=	16'h	751a;
16091	:douta	=	16'h	6cb9;
16092	:douta	=	16'h	857b;
16093	:douta	=	16'h	6cb9;
16094	:douta	=	16'h	6c58;
16095	:douta	=	16'h	6c78;
16096	:douta	=	16'h	6c98;
16097	:douta	=	16'h	7cf9;
16098	:douta	=	16'h	853a;
16099	:douta	=	16'h	8d9c;
16100	:douta	=	16'h	857b;
16101	:douta	=	16'h	855b;
16102	:douta	=	16'h	857c;
16103	:douta	=	16'h	8d9c;
16104	:douta	=	16'h	8d9c;
16105	:douta	=	16'h	7d3a;
16106	:douta	=	16'h	7d1a;
16107	:douta	=	16'h	7d3a;
16108	:douta	=	16'h	7d3a;
16109	:douta	=	16'h	853b;
16110	:douta	=	16'h	7d1a;
16111	:douta	=	16'h	855b;
16112	:douta	=	16'h	855b;
16113	:douta	=	16'h	853a;
16114	:douta	=	16'h	8d5b;
16115	:douta	=	16'h	7cf9;
16116	:douta	=	16'h	6478;
16117	:douta	=	16'h	7cd9;
16118	:douta	=	16'h	7cfa;
16119	:douta	=	16'h	2146;
16120	:douta	=	16'h	5b72;
16121	:douta	=	16'h	5330;
16122	:douta	=	16'h	9cd5;
16123	:douta	=	16'h	8cb4;
16124	:douta	=	16'h	a538;
16125	:douta	=	16'h	6392;
16126	:douta	=	16'h	63b3;
16127	:douta	=	16'h	5372;
16128	:douta	=	16'h	3b34;
16129	:douta	=	16'h	19cc;
16130	:douta	=	16'h	222f;
16131	:douta	=	16'h	3333;
16132	:douta	=	16'h	2a90;
16133	:douta	=	16'h	2a90;
16134	:douta	=	16'h	6cb9;
16135	:douta	=	16'h	53d4;
16136	:douta	=	16'h	7476;
16137	:douta	=	16'h	6c15;
16138	:douta	=	16'h	6c56;
16139	:douta	=	16'h	5331;
16140	:douta	=	16'h	6bd3;
16141	:douta	=	16'h	8cf8;
16142	:douta	=	16'h	7c34;
16143	:douta	=	16'h	8c54;
16144	:douta	=	16'h	7413;
16145	:douta	=	16'h	9cd6;
16146	:douta	=	16'h	7c12;
16147	:douta	=	16'h	ad56;
16148	:douta	=	16'h	8c93;
16149	:douta	=	16'h	a514;
16150	:douta	=	16'h	7bcf;
16151	:douta	=	16'h	8c50;
16152	:douta	=	16'h	c594;
16153	:douta	=	16'h	c5f6;
16154	:douta	=	16'h	d657;
16155	:douta	=	16'h	d657;
16156	:douta	=	16'h	deb7;
16157	:douta	=	16'h	8c50;
16158	:douta	=	16'h	6b2c;
16159	:douta	=	16'h	8c71;
16160	:douta	=	16'h	8c10;
16161	:douta	=	16'h	8bac;
16162	:douta	=	16'h	8b8b;
16163	:douta	=	16'h	8bab;
16164	:douta	=	16'h	8349;
16165	:douta	=	16'h	b48d;
16166	:douta	=	16'h	8b8b;
16167	:douta	=	16'h	ac6b;
16168	:douta	=	16'h	b4ad;
16169	:douta	=	16'h	ac8d;
16170	:douta	=	16'h	b48d;
16171	:douta	=	16'h	d56f;
16172	:douta	=	16'h	d5b1;
16173	:douta	=	16'h	de33;
16174	:douta	=	16'h	e675;
16175	:douta	=	16'h	e675;
16176	:douta	=	16'h	e675;
16177	:douta	=	16'h	de33;
16178	:douta	=	16'h	ddf3;
16179	:douta	=	16'h	ddf3;
16180	:douta	=	16'h	e613;
16181	:douta	=	16'h	9c0d;
16182	:douta	=	16'h	c52f;
16183	:douta	=	16'h	bcae;
16184	:douta	=	16'h	bcce;
16185	:douta	=	16'h	8b8a;
16186	:douta	=	16'h	9c0c;
16187	:douta	=	16'h	b4ae;
16188	:douta	=	16'h	acad;
16189	:douta	=	16'h	c54f;
16190	:douta	=	16'h	cd90;
16191	:douta	=	16'h	d5d2;
16192	:douta	=	16'h	cd70;
16193	:douta	=	16'h	c550;
16194	:douta	=	16'h	bcf0;
16195	:douta	=	16'h	b4d0;
16196	:douta	=	16'h	ac8f;
16197	:douta	=	16'h	a470;
16198	:douta	=	16'h	942f;
16199	:douta	=	16'h	736e;
16200	:douta	=	16'h	7b6f;
16201	:douta	=	16'h	630e;
16202	:douta	=	16'h	52ce;
16203	:douta	=	16'h	428c;
16204	:douta	=	16'h	3a2c;
16205	:douta	=	16'h	31eb;
16206	:douta	=	16'h	21a9;
16207	:douta	=	16'h	1906;
16208	:douta	=	16'h	08c5;
16209	:douta	=	16'h	526b;
16210	:douta	=	16'h	0063;
16211	:douta	=	16'h	18a4;
16212	:douta	=	16'h	10e4;
16213	:douta	=	16'h	10a4;
16214	:douta	=	16'h	1084;
16215	:douta	=	16'h	08a4;
16216	:douta	=	16'h	2146;
16217	:douta	=	16'h	18e5;
16218	:douta	=	16'h	0000;
16219	:douta	=	16'h	2988;
16220	:douta	=	16'h	5b50;
16221	:douta	=	16'h	4acd;
16222	:douta	=	16'h	6baf;
16223	:douta	=	16'h	0001;
16224	:douta	=	16'h	52ca;
16225	:douta	=	16'h	0842;
16226	:douta	=	16'h	08c3;
16227	:douta	=	16'h	62aa;
16228	:douta	=	16'h	2146;
16229	:douta	=	16'h	5289;
16230	:douta	=	16'h	3186;
16231	:douta	=	16'h	6b4c;
16232	:douta	=	16'h	5269;
16233	:douta	=	16'h	52ec;
16234	:douta	=	16'h	7b8d;
16235	:douta	=	16'h	b532;
16236	:douta	=	16'h	4a4b;
16237	:douta	=	16'h	6b2d;
16238	:douta	=	16'h	1948;
16239	:douta	=	16'h	636f;
16240	:douta	=	16'h	21a9;
16241	:douta	=	16'h	8430;
16242	:douta	=	16'h	426c;
16243	:douta	=	16'h	7bef;
16244	:douta	=	16'h	8c0f;
16245	:douta	=	16'h	732b;
16246	:douta	=	16'h	8d39;
16247	:douta	=	16'h	84b7;
16248	:douta	=	16'h	8d18;
16249	:douta	=	16'h	8d39;
16250	:douta	=	16'h	8d39;
16251	:douta	=	16'h	9579;
16252	:douta	=	16'h	a5ba;
16253	:douta	=	16'h	9579;
16254	:douta	=	16'h	8518;
16255	:douta	=	16'h	8d39;
16256	:douta	=	16'h	8d38;
16257	:douta	=	16'h	8d38;
16258	:douta	=	16'h	9579;
16259	:douta	=	16'h	a5ba;
16260	:douta	=	16'h	9579;
16261	:douta	=	16'h	957a;
16262	:douta	=	16'h	9d9a;
16263	:douta	=	16'h	9d9a;
16264	:douta	=	16'h	9dba;
16265	:douta	=	16'h	9dba;
16266	:douta	=	16'h	ae3c;
16267	:douta	=	16'h	8d39;
16268	:douta	=	16'h	9d59;
16269	:douta	=	16'h	5bf6;
16270	:douta	=	16'h	5bf6;
16271	:douta	=	16'h	9dbb;
16272	:douta	=	16'h	a5dc;
16273	:douta	=	16'h	955b;
16274	:douta	=	16'h	957a;
16275	:douta	=	16'h	95bb;
16276	:douta	=	16'h	a5fc;
16277	:douta	=	16'h	959b;
16278	:douta	=	16'h	853a;
16279	:douta	=	16'h	6c58;
16280	:douta	=	16'h	7cf9;
16281	:douta	=	16'h	7cf9;
16282	:douta	=	16'h	8519;
16283	:douta	=	16'h	a5fc;
16284	:douta	=	16'h	74b8;
16285	:douta	=	16'h	6c56;
16286	:douta	=	16'h	7c76;
16287	:douta	=	16'h	8518;
16288	:douta	=	16'h	a5db;
16289	:douta	=	16'h	94d6;
16290	:douta	=	16'h	8bad;
16291	:douta	=	16'h	1925;
16292	:douta	=	16'h	1905;
16293	:douta	=	16'h	0883;
16294	:douta	=	16'h	6c15;
16295	:douta	=	16'h	4b32;
16296	:douta	=	16'h	7497;
16297	:douta	=	16'h	7cd8;
16298	:douta	=	16'h	7cd9;
16299	:douta	=	16'h	7497;
16300	:douta	=	16'h	7cd8;
16301	:douta	=	16'h	7498;
16302	:douta	=	16'h	6c15;
16303	:douta	=	16'h	7cb7;
16304	:douta	=	16'h	6c35;
16305	:douta	=	16'h	7456;
16306	:douta	=	16'h	7476;
16307	:douta	=	16'h	6415;
16308	:douta	=	16'h	4311;
16309	:douta	=	16'h	5393;
16310	:douta	=	16'h	6415;
16311	:douta	=	16'h	5b73;
16312	:douta	=	16'h	5b94;
16313	:douta	=	16'h	6c77;
16314	:douta	=	16'h	6437;
16315	:douta	=	16'h	6c77;
16316	:douta	=	16'h	7cb8;
16317	:douta	=	16'h	5373;
16318	:douta	=	16'h	63d4;
16319	:douta	=	16'h	5bb3;
16320	:douta	=	16'h	7c56;
16321	:douta	=	16'h	5372;
16322	:douta	=	16'h	63d3;
16323	:douta	=	16'h	9d9a;
16324	:douta	=	16'h	84d7;
16325	:douta	=	16'h	7c34;
16326	:douta	=	16'h	6bd1;
16327	:douta	=	16'h	2967;
16328	:douta	=	16'h	1905;
16329	:douta	=	16'h	10e5;
16330	:douta	=	16'h	0884;
16331	:douta	=	16'h	7cd9;
16332	:douta	=	16'h	7477;
16333	:douta	=	16'h	6c57;
16334	:douta	=	16'h	6457;
16335	:douta	=	16'h	6cb9;
16336	:douta	=	16'h	5c37;
16337	:douta	=	16'h	53b6;
16338	:douta	=	16'h	5c58;
16339	:douta	=	16'h	6479;
16340	:douta	=	16'h	6499;
16341	:douta	=	16'h	74fa;
16342	:douta	=	16'h	74d9;
16343	:douta	=	16'h	5c37;
16344	:douta	=	16'h	53d5;
16345	:douta	=	16'h	53f6;
16346	:douta	=	16'h	6437;
16347	:douta	=	16'h	74f9;
16348	:douta	=	16'h	74d9;
16349	:douta	=	16'h	7d1a;
16350	:douta	=	16'h	74d9;
16351	:douta	=	16'h	7d3a;
16352	:douta	=	16'h	7d1a;
16353	:douta	=	16'h	7478;
16354	:douta	=	16'h	7477;
16355	:douta	=	16'h	6416;
16356	:douta	=	16'h	7d3a;
16357	:douta	=	16'h	855b;
16358	:douta	=	16'h	853b;
16359	:douta	=	16'h	8d9c;
16360	:douta	=	16'h	7d3a;
16361	:douta	=	16'h	7d3a;
16362	:douta	=	16'h	8d5b;
16363	:douta	=	16'h	7d1a;
16364	:douta	=	16'h	7d3a;
16365	:douta	=	16'h	8dbc;
16366	:douta	=	16'h	74b9;
16367	:douta	=	16'h	7cd9;
16368	:douta	=	16'h	7d1a;
16369	:douta	=	16'h	855b;
16370	:douta	=	16'h	8d9b;
16371	:douta	=	16'h	853a;
16372	:douta	=	16'h	7d1a;
16373	:douta	=	16'h	7d3a;
16374	:douta	=	16'h	7498;
16375	:douta	=	16'h	39ea;
16376	:douta	=	16'h	b5b8;
16377	:douta	=	16'h	9d57;
16378	:douta	=	16'h	b5b8;
16379	:douta	=	16'h	7413;
16380	:douta	=	16'h	42af;
16381	:douta	=	16'h	73f3;
16382	:douta	=	16'h	8c94;
16383	:douta	=	16'h	9517;
16384	:douta	=	16'h	3b13;
16385	:douta	=	16'h	2ab1;
16386	:douta	=	16'h	3b33;
16387	:douta	=	16'h	4b94;
16388	:douta	=	16'h	2a6f;
16389	:douta	=	16'h	222e;
16390	:douta	=	16'h	53d5;
16391	:douta	=	16'h	4b73;
16392	:douta	=	16'h	63d4;
16393	:douta	=	16'h	63f4;
16394	:douta	=	16'h	7477;
16395	:douta	=	16'h	5b72;
16396	:douta	=	16'h	4b10;
16397	:douta	=	16'h	7c55;
16398	:douta	=	16'h	5b91;
16399	:douta	=	16'h	7c13;
16400	:douta	=	16'h	8473;
16401	:douta	=	16'h	9d36;
16402	:douta	=	16'h	8c73;
16403	:douta	=	16'h	ad34;
16404	:douta	=	16'h	5b2f;
16405	:douta	=	16'h	a514;
16406	:douta	=	16'h	9c92;
16407	:douta	=	16'h	b574;
16408	:douta	=	16'h	9c90;
16409	:douta	=	16'h	7c0f;
16410	:douta	=	16'h	9c91;
16411	:douta	=	16'h	bd94;
16412	:douta	=	16'h	bd94;
16413	:douta	=	16'h	ce16;
16414	:douta	=	16'h	b574;
16415	:douta	=	16'h	be17;
16416	:douta	=	16'h	6b2b;
16417	:douta	=	16'h	8b8b;
16418	:douta	=	16'h	8bab;
16419	:douta	=	16'h	838a;
16420	:douta	=	16'h	8b8b;
16421	:douta	=	16'h	ac6c;
16422	:douta	=	16'h	9bca;
16423	:douta	=	16'h	ac8c;
16424	:douta	=	16'h	b4ad;
16425	:douta	=	16'h	b4ad;
16426	:douta	=	16'h	bcad;
16427	:douta	=	16'h	d5b0;
16428	:douta	=	16'h	de12;
16429	:douta	=	16'h	e633;
16430	:douta	=	16'h	ee96;
16431	:douta	=	16'h	e675;
16432	:douta	=	16'h	e634;
16433	:douta	=	16'h	de34;
16434	:douta	=	16'h	ddf2;
16435	:douta	=	16'h	d5d1;
16436	:douta	=	16'h	ddb2;
16437	:douta	=	16'h	a44e;
16438	:douta	=	16'h	9c0d;
16439	:douta	=	16'h	c50f;
16440	:douta	=	16'h	8b8a;
16441	:douta	=	16'h	8b8a;
16442	:douta	=	16'h	93aa;
16443	:douta	=	16'h	a44d;
16444	:douta	=	16'h	b4ad;
16445	:douta	=	16'h	cd70;
16446	:douta	=	16'h	cd91;
16447	:douta	=	16'h	d5d2;
16448	:douta	=	16'h	cd71;
16449	:douta	=	16'h	cd70;
16450	:douta	=	16'h	c530;
16451	:douta	=	16'h	bd10;
16452	:douta	=	16'h	ac8f;
16453	:douta	=	16'h	a450;
16454	:douta	=	16'h	9450;
16455	:douta	=	16'h	7b8f;
16456	:douta	=	16'h	7b8f;
16457	:douta	=	16'h	634e;
16458	:douta	=	16'h	52ce;
16459	:douta	=	16'h	4acd;
16460	:douta	=	16'h	428d;
16461	:douta	=	16'h	3a4c;
16462	:douta	=	16'h	29eb;
16463	:douta	=	16'h	29a9;
16464	:douta	=	16'h	1948;
16465	:douta	=	16'h	62ec;
16466	:douta	=	16'h	41e9;
16467	:douta	=	16'h	10a4;
16468	:douta	=	16'h	10c5;
16469	:douta	=	16'h	10a4;
16470	:douta	=	16'h	1084;
16471	:douta	=	16'h	1083;
16472	:douta	=	16'h	18e5;
16473	:douta	=	16'h	2146;
16474	:douta	=	16'h	0000;
16475	:douta	=	16'h	0000;
16476	:douta	=	16'h	29ca;
16477	:douta	=	16'h	5b2e;
16478	:douta	=	16'h	42ad;
16479	:douta	=	16'h	3166;
16480	:douta	=	16'h	0862;
16481	:douta	=	16'h	0842;
16482	:douta	=	16'h	0000;
16483	:douta	=	16'h	18c3;
16484	:douta	=	16'h	2125;
16485	:douta	=	16'h	52a9;
16486	:douta	=	16'h	2105;
16487	:douta	=	16'h	3a09;
16488	:douta	=	16'h	4208;
16489	:douta	=	16'h	3a29;
16490	:douta	=	16'h	2988;
16491	:douta	=	16'h	9c70;
16492	:douta	=	16'h	31a8;
16493	:douta	=	16'h	9471;
16494	:douta	=	16'h	5acd;
16495	:douta	=	16'h	4aad;
16496	:douta	=	16'h	424c;
16497	:douta	=	16'h	1127;
16498	:douta	=	16'h	29a9;
16499	:douta	=	16'h	3a6b;
16500	:douta	=	16'h	628a;
16501	:douta	=	16'h	730b;
16502	:douta	=	16'h	9d9a;
16503	:douta	=	16'h	9559;
16504	:douta	=	16'h	8d18;
16505	:douta	=	16'h	9559;
16506	:douta	=	16'h	8d38;
16507	:douta	=	16'h	9559;
16508	:douta	=	16'h	8d18;
16509	:douta	=	16'h	8d18;
16510	:douta	=	16'h	8d18;
16511	:douta	=	16'h	8d18;
16512	:douta	=	16'h	9579;
16513	:douta	=	16'h	9559;
16514	:douta	=	16'h	959a;
16515	:douta	=	16'h	959a;
16516	:douta	=	16'h	957a;
16517	:douta	=	16'h	84d7;
16518	:douta	=	16'h	84f8;
16519	:douta	=	16'h	a5ba;
16520	:douta	=	16'h	957a;
16521	:douta	=	16'h	957a;
16522	:douta	=	16'h	a5fa;
16523	:douta	=	16'h	b63b;
16524	:douta	=	16'h	be7c;
16525	:douta	=	16'h	a5ba;
16526	:douta	=	16'h	8cf8;
16527	:douta	=	16'h	6457;
16528	:douta	=	16'h	7478;
16529	:douta	=	16'h	8d3a;
16530	:douta	=	16'h	957b;
16531	:douta	=	16'h	7cf9;
16532	:douta	=	16'h	8539;
16533	:douta	=	16'h	8d3a;
16534	:douta	=	16'h	be9d;
16535	:douta	=	16'h	851a;
16536	:douta	=	16'h	8d7b;
16537	:douta	=	16'h	6457;
16538	:douta	=	16'h	7498;
16539	:douta	=	16'h	955b;
16540	:douta	=	16'h	8d5a;
16541	:douta	=	16'h	8518;
16542	:douta	=	16'h	63f5;
16543	:douta	=	16'h	5b93;
16544	:douta	=	16'h	8d19;
16545	:douta	=	16'h	8d18;
16546	:douta	=	16'h	93ef;
16547	:douta	=	16'h	2146;
16548	:douta	=	16'h	18e5;
16549	:douta	=	16'h	0042;
16550	:douta	=	16'h	a5bb;
16551	:douta	=	16'h	8d18;
16552	:douta	=	16'h	6415;
16553	:douta	=	16'h	9518;
16554	:douta	=	16'h	8539;
16555	:douta	=	16'h	8519;
16556	:douta	=	16'h	853a;
16557	:douta	=	16'h	7c98;
16558	:douta	=	16'h	7477;
16559	:douta	=	16'h	8d39;
16560	:douta	=	16'h	955a;
16561	:douta	=	16'h	6c36;
16562	:douta	=	16'h	7cd8;
16563	:douta	=	16'h	855b;
16564	:douta	=	16'h	7cd8;
16565	:douta	=	16'h	63f4;
16566	:douta	=	16'h	5373;
16567	:douta	=	16'h	6435;
16568	:douta	=	16'h	6c15;
16569	:douta	=	16'h	6416;
16570	:douta	=	16'h	7cd9;
16571	:douta	=	16'h	74b7;
16572	:douta	=	16'h	6c36;
16573	:douta	=	16'h	6c36;
16574	:douta	=	16'h	84b7;
16575	:douta	=	16'h	63f4;
16576	:douta	=	16'h	63d3;
16577	:douta	=	16'h	7435;
16578	:douta	=	16'h	63b3;
16579	:douta	=	16'h	6c35;
16580	:douta	=	16'h	957a;
16581	:douta	=	16'h	6bf3;
16582	:douta	=	16'h	6bb1;
16583	:douta	=	16'h	2105;
16584	:douta	=	16'h	18e5;
16585	:douta	=	16'h	10e5;
16586	:douta	=	16'h	10e5;
16587	:douta	=	16'h	7cb8;
16588	:douta	=	16'h	6c77;
16589	:douta	=	16'h	6c77;
16590	:douta	=	16'h	7498;
16591	:douta	=	16'h	6458;
16592	:douta	=	16'h	6c99;
16593	:douta	=	16'h	6c99;
16594	:douta	=	16'h	4bd6;
16595	:douta	=	16'h	53d6;
16596	:douta	=	16'h	5c17;
16597	:douta	=	16'h	6c99;
16598	:douta	=	16'h	6478;
16599	:douta	=	16'h	6cb9;
16600	:douta	=	16'h	74d9;
16601	:douta	=	16'h	6457;
16602	:douta	=	16'h	6457;
16603	:douta	=	16'h	6cb8;
16604	:douta	=	16'h	7d1a;
16605	:douta	=	16'h	74d9;
16606	:douta	=	16'h	6c98;
16607	:douta	=	16'h	7d1a;
16608	:douta	=	16'h	851a;
16609	:douta	=	16'h	7cd9;
16610	:douta	=	16'h	851a;
16611	:douta	=	16'h	6c37;
16612	:douta	=	16'h	7cb9;
16613	:douta	=	16'h	74b9;
16614	:douta	=	16'h	74b9;
16615	:douta	=	16'h	7cf9;
16616	:douta	=	16'h	8dbc;
16617	:douta	=	16'h	7d3b;
16618	:douta	=	16'h	7cda;
16619	:douta	=	16'h	8dbc;
16620	:douta	=	16'h	857b;
16621	:douta	=	16'h	7d3b;
16622	:douta	=	16'h	8d7c;
16623	:douta	=	16'h	7d3b;
16624	:douta	=	16'h	855b;
16625	:douta	=	16'h	7d1b;
16626	:douta	=	16'h	853a;
16627	:douta	=	16'h	7cd9;
16628	:douta	=	16'h	7d1a;
16629	:douta	=	16'h	7d1a;
16630	:douta	=	16'h	7477;
16631	:douta	=	16'h	2968;
16632	:douta	=	16'h	7433;
16633	:douta	=	16'h	63b3;
16634	:douta	=	16'h	b5d8;
16635	:douta	=	16'h	73f3;
16636	:douta	=	16'h	7434;
16637	:douta	=	16'h	8454;
16638	:douta	=	16'h	42d0;
16639	:douta	=	16'h	52ce;
16640	:douta	=	16'h	3b12;
16641	:douta	=	16'h	2a90;
16642	:douta	=	16'h	3b13;
16643	:douta	=	16'h	3313;
16644	:douta	=	16'h	2a70;
16645	:douta	=	16'h	2a90;
16646	:douta	=	16'h	6c98;
16647	:douta	=	16'h	6457;
16648	:douta	=	16'h	7c98;
16649	:douta	=	16'h	8519;
16650	:douta	=	16'h	6c56;
16651	:douta	=	16'h	5b93;
16652	:douta	=	16'h	5331;
16653	:douta	=	16'h	6392;
16654	:douta	=	16'h	6bf4;
16655	:douta	=	16'h	7c54;
16656	:douta	=	16'h	8434;
16657	:douta	=	16'h	94b5;
16658	:douta	=	16'h	73d2;
16659	:douta	=	16'h	b5b6;
16660	:douta	=	16'h	8452;
16661	:douta	=	16'h	a4f3;
16662	:douta	=	16'h	a4f3;
16663	:douta	=	16'h	b533;
16664	:douta	=	16'h	e6b9;
16665	:douta	=	16'h	ad54;
16666	:douta	=	16'h	b573;
16667	:douta	=	16'h	d677;
16668	:douta	=	16'h	de77;
16669	:douta	=	16'h	9491;
16670	:douta	=	16'h	9471;
16671	:douta	=	16'h	72c8;
16672	:douta	=	16'h	8b6a;
16673	:douta	=	16'h	8b8b;
16674	:douta	=	16'h	93aa;
16675	:douta	=	16'h	a42b;
16676	:douta	=	16'h	9beb;
16677	:douta	=	16'h	8b69;
16678	:douta	=	16'h	c52d;
16679	:douta	=	16'h	bccd;
16680	:douta	=	16'h	c52e;
16681	:douta	=	16'h	cd2e;
16682	:douta	=	16'h	cd4f;
16683	:douta	=	16'h	e634;
16684	:douta	=	16'h	ee96;
16685	:douta	=	16'h	ee96;
16686	:douta	=	16'h	e654;
16687	:douta	=	16'h	eeb6;
16688	:douta	=	16'h	de34;
16689	:douta	=	16'h	ddf4;
16690	:douta	=	16'h	e675;
16691	:douta	=	16'h	bd0f;
16692	:douta	=	16'h	cd71;
16693	:douta	=	16'h	ac4d;
16694	:douta	=	16'h	9c2d;
16695	:douta	=	16'h	7b07;
16696	:douta	=	16'h	d570;
16697	:douta	=	16'h	c52f;
16698	:douta	=	16'h	93eb;
16699	:douta	=	16'h	a42c;
16700	:douta	=	16'h	b4ad;
16701	:douta	=	16'h	d5b2;
16702	:douta	=	16'h	ddf3;
16703	:douta	=	16'h	d5b2;
16704	:douta	=	16'h	d5b2;
16705	:douta	=	16'h	cd71;
16706	:douta	=	16'h	c550;
16707	:douta	=	16'h	c530;
16708	:douta	=	16'h	acaf;
16709	:douta	=	16'h	9c70;
16710	:douta	=	16'h	9430;
16711	:douta	=	16'h	83ef;
16712	:douta	=	16'h	7baf;
16713	:douta	=	16'h	6b6f;
16714	:douta	=	16'h	634f;
16715	:douta	=	16'h	5b2e;
16716	:douta	=	16'h	52ce;
16717	:douta	=	16'h	428d;
16718	:douta	=	16'h	320b;
16719	:douta	=	16'h	29aa;
16720	:douta	=	16'h	29aa;
16721	:douta	=	16'h	08e6;
16722	:douta	=	16'h	31c8;
16723	:douta	=	16'h	08a4;
16724	:douta	=	16'h	10c3;
16725	:douta	=	16'h	10a4;
16726	:douta	=	16'h	10c4;
16727	:douta	=	16'h	10c4;
16728	:douta	=	16'h	18e4;
16729	:douta	=	16'h	10e4;
16730	:douta	=	16'h	18e5;
16731	:douta	=	16'h	2125;
16732	:douta	=	16'h	0000;
16733	:douta	=	16'h	2a2c;
16734	:douta	=	16'h	7475;
16735	:douta	=	16'h	5b0e;
16736	:douta	=	16'h	736d;
16737	:douta	=	16'h	8c50;
16738	:douta	=	16'h	7b8c;
16739	:douta	=	16'h	ad11;
16740	:douta	=	16'h	4207;
16741	:douta	=	16'h	5aaa;
16742	:douta	=	16'h	5a89;
16743	:douta	=	16'h	0000;
16744	:douta	=	16'h	0000;
16745	:douta	=	16'h	0042;
16746	:douta	=	16'h	41e7;
16747	:douta	=	16'h	83ee;
16748	:douta	=	16'h	8c70;
16749	:douta	=	16'h	73ef;
16750	:douta	=	16'h	39c8;
16751	:douta	=	16'h	39ea;
16752	:douta	=	16'h	3a09;
16753	:douta	=	16'h	29a8;
16754	:douta	=	16'h	3a2b;
16755	:douta	=	16'h	5b0d;
16756	:douta	=	16'h	b512;
16757	:douta	=	16'h	7b6c;
16758	:douta	=	16'h	9dba;
16759	:douta	=	16'h	8517;
16760	:douta	=	16'h	8d38;
16761	:douta	=	16'h	8d18;
16762	:douta	=	16'h	84d7;
16763	:douta	=	16'h	84f8;
16764	:douta	=	16'h	84f8;
16765	:douta	=	16'h	8d18;
16766	:douta	=	16'h	9599;
16767	:douta	=	16'h	8d38;
16768	:douta	=	16'h	9559;
16769	:douta	=	16'h	9559;
16770	:douta	=	16'h	9559;
16771	:douta	=	16'h	8d59;
16772	:douta	=	16'h	9599;
16773	:douta	=	16'h	9dba;
16774	:douta	=	16'h	9d9a;
16775	:douta	=	16'h	9559;
16776	:douta	=	16'h	8d59;
16777	:douta	=	16'h	9559;
16778	:douta	=	16'h	a5da;
16779	:douta	=	16'h	957a;
16780	:douta	=	16'h	9d9a;
16781	:douta	=	16'h	a5ba;
16782	:douta	=	16'h	adfb;
16783	:douta	=	16'h	9dda;
16784	:douta	=	16'h	9dda;
16785	:douta	=	16'h	9d9a;
16786	:douta	=	16'h	84f9;
16787	:douta	=	16'h	7498;
16788	:douta	=	16'h	8519;
16789	:douta	=	16'h	8d5a;
16790	:douta	=	16'h	8d7b;
16791	:douta	=	16'h	95bb;
16792	:douta	=	16'h	959b;
16793	:douta	=	16'h	a5fc;
16794	:douta	=	16'h	9ddc;
16795	:douta	=	16'h	8d3a;
16796	:douta	=	16'h	7cd8;
16797	:douta	=	16'h	7c77;
16798	:douta	=	16'h	7c97;
16799	:douta	=	16'h	7cb7;
16800	:douta	=	16'h	7cb7;
16801	:douta	=	16'h	84f9;
16802	:douta	=	16'h	9493;
16803	:douta	=	16'h	4a09;
16804	:douta	=	16'h	10e5;
16805	:douta	=	16'h	10c4;
16806	:douta	=	16'h	7c76;
16807	:douta	=	16'h	9539;
16808	:douta	=	16'h	7c96;
16809	:douta	=	16'h	7c97;
16810	:douta	=	16'h	957a;
16811	:douta	=	16'h	84d8;
16812	:douta	=	16'h	7c98;
16813	:douta	=	16'h	9d9b;
16814	:douta	=	16'h	a5fc;
16815	:douta	=	16'h	84d8;
16816	:douta	=	16'h	7cb7;
16817	:douta	=	16'h	63f4;
16818	:douta	=	16'h	84f9;
16819	:douta	=	16'h	959b;
16820	:douta	=	16'h	8d9b;
16821	:douta	=	16'h	853a;
16822	:douta	=	16'h	7477;
16823	:douta	=	16'h	8d19;
16824	:douta	=	16'h	7cd8;
16825	:douta	=	16'h	63b4;
16826	:douta	=	16'h	6c15;
16827	:douta	=	16'h	63d4;
16828	:douta	=	16'h	7c97;
16829	:douta	=	16'h	84f8;
16830	:douta	=	16'h	7476;
16831	:douta	=	16'h	7456;
16832	:douta	=	16'h	6c36;
16833	:douta	=	16'h	7cd8;
16834	:douta	=	16'h	7456;
16835	:douta	=	16'h	6bf5;
16836	:douta	=	16'h	5351;
16837	:douta	=	16'h	6c35;
16838	:douta	=	16'h	39ea;
16839	:douta	=	16'h	2125;
16840	:douta	=	16'h	1905;
16841	:douta	=	16'h	10e4;
16842	:douta	=	16'h	320b;
16843	:douta	=	16'h	6456;
16844	:douta	=	16'h	6c36;
16845	:douta	=	16'h	6436;
16846	:douta	=	16'h	6416;
16847	:douta	=	16'h	74d9;
16848	:douta	=	16'h	74d9;
16849	:douta	=	16'h	74d9;
16850	:douta	=	16'h	751b;
16851	:douta	=	16'h	6cda;
16852	:douta	=	16'h	751a;
16853	:douta	=	16'h	6c78;
16854	:douta	=	16'h	6457;
16855	:douta	=	16'h	6457;
16856	:douta	=	16'h	6478;
16857	:douta	=	16'h	6c98;
16858	:douta	=	16'h	6457;
16859	:douta	=	16'h	7498;
16860	:douta	=	16'h	63f5;
16861	:douta	=	16'h	6c36;
16862	:douta	=	16'h	7cf9;
16863	:douta	=	16'h	7cd9;
16864	:douta	=	16'h	74b8;
16865	:douta	=	16'h	74b8;
16866	:douta	=	16'h	8d7b;
16867	:douta	=	16'h	7cd9;
16868	:douta	=	16'h	74b8;
16869	:douta	=	16'h	855b;
16870	:douta	=	16'h	7498;
16871	:douta	=	16'h	7cb8;
16872	:douta	=	16'h	7498;
16873	:douta	=	16'h	74d9;
16874	:douta	=	16'h	74b9;
16875	:douta	=	16'h	7cf9;
16876	:douta	=	16'h	7cfa;
16877	:douta	=	16'h	855b;
16878	:douta	=	16'h	7d1a;
16879	:douta	=	16'h	74d9;
16880	:douta	=	16'h	7d1a;
16881	:douta	=	16'h	8d7b;
16882	:douta	=	16'h	851a;
16883	:douta	=	16'h	7cb9;
16884	:douta	=	16'h	7cfa;
16885	:douta	=	16'h	7d3a;
16886	:douta	=	16'h	6c15;
16887	:douta	=	16'h	7c53;
16888	:douta	=	16'h	ad98;
16889	:douta	=	16'h	84b6;
16890	:douta	=	16'h	8494;
16891	:douta	=	16'h	6391;
16892	:douta	=	16'h	7c33;
16893	:douta	=	16'h	6391;
16894	:douta	=	16'h	7434;
16895	:douta	=	16'h	20e3;
16896	:douta	=	16'h	2a0d;
16897	:douta	=	16'h	32d2;
16898	:douta	=	16'h	4374;
16899	:douta	=	16'h	5c58;
16900	:douta	=	16'h	4bd6;
16901	:douta	=	16'h	32d2;
16902	:douta	=	16'h	3b33;
16903	:douta	=	16'h	53f6;
16904	:douta	=	16'h	63f5;
16905	:douta	=	16'h	63f5;
16906	:douta	=	16'h	7478;
16907	:douta	=	16'h	7436;
16908	:douta	=	16'h	63b2;
16909	:douta	=	16'h	8476;
16910	:douta	=	16'h	5b93;
16911	:douta	=	16'h	4aef;
16912	:douta	=	16'h	73d2;
16913	:douta	=	16'h	7c33;
16914	:douta	=	16'h	8cb4;
16915	:douta	=	16'h	bdd8;
16916	:douta	=	16'h	8433;
16917	:douta	=	16'h	bd74;
16918	:douta	=	16'h	8411;
16919	:douta	=	16'h	cdf6;
16920	:douta	=	16'h	c5f5;
16921	:douta	=	16'h	b575;
16922	:douta	=	16'h	d616;
16923	:douta	=	16'h	d657;
16924	:douta	=	16'h	b574;
16925	:douta	=	16'h	c5f6;
16926	:douta	=	16'h	946f;
16927	:douta	=	16'h	938b;
16928	:douta	=	16'h	8b8b;
16929	:douta	=	16'h	93ab;
16930	:douta	=	16'h	9bcb;
16931	:douta	=	16'h	ac4b;
16932	:douta	=	16'h	ac6c;
16933	:douta	=	16'h	9389;
16934	:douta	=	16'h	cd4e;
16935	:douta	=	16'h	bced;
16936	:douta	=	16'h	cd4e;
16937	:douta	=	16'h	cd70;
16938	:douta	=	16'h	d590;
16939	:douta	=	16'h	e654;
16940	:douta	=	16'h	ee96;
16941	:douta	=	16'h	ee95;
16942	:douta	=	16'h	e654;
16943	:douta	=	16'h	e654;
16944	:douta	=	16'h	e654;
16945	:douta	=	16'h	d591;
16946	:douta	=	16'h	de34;
16947	:douta	=	16'h	b4cf;
16948	:douta	=	16'h	bcd0;
16949	:douta	=	16'h	a44d;
16950	:douta	=	16'h	7b29;
16951	:douta	=	16'h	834a;
16952	:douta	=	16'h	d570;
16953	:douta	=	16'h	ddd2;
16954	:douta	=	16'h	bd0e;
16955	:douta	=	16'h	bd2f;
16956	:douta	=	16'h	c52f;
16957	:douta	=	16'h	d5f2;
16958	:douta	=	16'h	ddf3;
16959	:douta	=	16'h	d5d2;
16960	:douta	=	16'h	d591;
16961	:douta	=	16'h	cd71;
16962	:douta	=	16'h	cd71;
16963	:douta	=	16'h	cd71;
16964	:douta	=	16'h	b4d0;
16965	:douta	=	16'h	a470;
16966	:douta	=	16'h	9c50;
16967	:douta	=	16'h	8c10;
16968	:douta	=	16'h	7bcf;
16969	:douta	=	16'h	738f;
16970	:douta	=	16'h	636f;
16971	:douta	=	16'h	5b2e;
16972	:douta	=	16'h	52cf;
16973	:douta	=	16'h	426d;
16974	:douta	=	16'h	29eb;
16975	:douta	=	16'h	31eb;
16976	:douta	=	16'h	29ca;
16977	:douta	=	16'h	29c9;
16978	:douta	=	16'h	10e6;
16979	:douta	=	16'h	424a;
16980	:douta	=	16'h	10a4;
16981	:douta	=	16'h	10c4;
16982	:douta	=	16'h	10a4;
16983	:douta	=	16'h	10e4;
16984	:douta	=	16'h	1904;
16985	:douta	=	16'h	10e4;
16986	:douta	=	16'h	10c4;
16987	:douta	=	16'h	1906;
16988	:douta	=	16'h	2146;
16989	:douta	=	16'h	0000;
16990	:douta	=	16'h	29eb;
16991	:douta	=	16'h	5b0e;
16992	:douta	=	16'h	3a6b;
16993	:douta	=	16'h	08a4;
16994	:douta	=	16'h	5a49;
16995	:douta	=	16'h	944d;
16996	:douta	=	16'h	3165;
16997	:douta	=	16'h	630a;
16998	:douta	=	16'h	8bed;
16999	:douta	=	16'h	736c;
17000	:douta	=	16'h	5aa9;
17001	:douta	=	16'h	39a7;
17002	:douta	=	16'h	2146;
17003	:douta	=	16'h	0885;
17004	:douta	=	16'h	21a9;
17005	:douta	=	16'h	29c8;
17006	:douta	=	16'h	8c2f;
17007	:douta	=	16'h	5aab;
17008	:douta	=	16'h	a4d1;
17009	:douta	=	16'h	31e9;
17010	:douta	=	16'h	632d;
17011	:douta	=	16'h	426c;
17012	:douta	=	16'h	736e;
17013	:douta	=	16'h	6aec;
17014	:douta	=	16'h	b65c;
17015	:douta	=	16'h	9579;
17016	:douta	=	16'h	8d38;
17017	:douta	=	16'h	84f8;
17018	:douta	=	16'h	84f7;
17019	:douta	=	16'h	8d58;
17020	:douta	=	16'h	8d58;
17021	:douta	=	16'h	84f8;
17022	:douta	=	16'h	7cb7;
17023	:douta	=	16'h	84f8;
17024	:douta	=	16'h	8d38;
17025	:douta	=	16'h	9579;
17026	:douta	=	16'h	8d39;
17027	:douta	=	16'h	9559;
17028	:douta	=	16'h	9579;
17029	:douta	=	16'h	9559;
17030	:douta	=	16'h	8d39;
17031	:douta	=	16'h	8d39;
17032	:douta	=	16'h	9d9a;
17033	:douta	=	16'h	9579;
17034	:douta	=	16'h	9559;
17035	:douta	=	16'h	9559;
17036	:douta	=	16'h	9dba;
17037	:douta	=	16'h	9559;
17038	:douta	=	16'h	957a;
17039	:douta	=	16'h	adfa;
17040	:douta	=	16'h	9d9a;
17041	:douta	=	16'h	adfb;
17042	:douta	=	16'h	a5fb;
17043	:douta	=	16'h	9d9a;
17044	:douta	=	16'h	7cd9;
17045	:douta	=	16'h	74b8;
17046	:douta	=	16'h	7c97;
17047	:douta	=	16'h	957a;
17048	:douta	=	16'h	ae3c;
17049	:douta	=	16'h	95bb;
17050	:douta	=	16'h	84f9;
17051	:douta	=	16'h	a5dc;
17052	:douta	=	16'h	957a;
17053	:douta	=	16'h	8d19;
17054	:douta	=	16'h	7435;
17055	:douta	=	16'h	84d7;
17056	:douta	=	16'h	7cb7;
17057	:douta	=	16'h	7477;
17058	:douta	=	16'h	8474;
17059	:douta	=	16'h	5249;
17060	:douta	=	16'h	1905;
17061	:douta	=	16'h	10e5;
17062	:douta	=	16'h	5b91;
17063	:douta	=	16'h	9559;
17064	:douta	=	16'h	8d18;
17065	:douta	=	16'h	84f8;
17066	:douta	=	16'h	9579;
17067	:douta	=	16'h	9d9a;
17068	:douta	=	16'h	9dbb;
17069	:douta	=	16'h	7cb8;
17070	:douta	=	16'h	8d3a;
17071	:douta	=	16'h	8d18;
17072	:douta	=	16'h	8d39;
17073	:douta	=	16'h	8519;
17074	:douta	=	16'h	7cb8;
17075	:douta	=	16'h	7cf9;
17076	:douta	=	16'h	9ddc;
17077	:douta	=	16'h	a63e;
17078	:douta	=	16'h	84f9;
17079	:douta	=	16'h	7cb7;
17080	:douta	=	16'h	84d9;
17081	:douta	=	16'h	7c97;
17082	:douta	=	16'h	7cb7;
17083	:douta	=	16'h	6c35;
17084	:douta	=	16'h	6c14;
17085	:douta	=	16'h	7435;
17086	:douta	=	16'h	84d7;
17087	:douta	=	16'h	9559;
17088	:douta	=	16'h	84d8;
17089	:douta	=	16'h	6c35;
17090	:douta	=	16'h	63d4;
17091	:douta	=	16'h	6bf4;
17092	:douta	=	16'h	6c35;
17093	:douta	=	16'h	6c15;
17094	:douta	=	16'h	39a8;
17095	:douta	=	16'h	2126;
17096	:douta	=	16'h	1905;
17097	:douta	=	16'h	10e4;
17098	:douta	=	16'h	4ad0;
17099	:douta	=	16'h	6436;
17100	:douta	=	16'h	5bf5;
17101	:douta	=	16'h	6415;
17102	:douta	=	16'h	7498;
17103	:douta	=	16'h	6457;
17104	:douta	=	16'h	6cb9;
17105	:douta	=	16'h	6478;
17106	:douta	=	16'h	6cda;
17107	:douta	=	16'h	751b;
17108	:douta	=	16'h	5c16;
17109	:douta	=	16'h	74b9;
17110	:douta	=	16'h	74f9;
17111	:douta	=	16'h	5c37;
17112	:douta	=	16'h	6c78;
17113	:douta	=	16'h	6c98;
17114	:douta	=	16'h	74b9;
17115	:douta	=	16'h	7cd9;
17116	:douta	=	16'h	7cf9;
17117	:douta	=	16'h	7cb8;
17118	:douta	=	16'h	7498;
17119	:douta	=	16'h	74b8;
17120	:douta	=	16'h	7cd9;
17121	:douta	=	16'h	7498;
17122	:douta	=	16'h	74b8;
17123	:douta	=	16'h	74b8;
17124	:douta	=	16'h	7cf9;
17125	:douta	=	16'h	6c57;
17126	:douta	=	16'h	8d5b;
17127	:douta	=	16'h	7cf9;
17128	:douta	=	16'h	851a;
17129	:douta	=	16'h	74f9;
17130	:douta	=	16'h	7d1a;
17131	:douta	=	16'h	6457;
17132	:douta	=	16'h	7cd9;
17133	:douta	=	16'h	74d9;
17134	:douta	=	16'h	7d1a;
17135	:douta	=	16'h	7d1a;
17136	:douta	=	16'h	7cd9;
17137	:douta	=	16'h	7499;
17138	:douta	=	16'h	8d7b;
17139	:douta	=	16'h	7cf9;
17140	:douta	=	16'h	74b8;
17141	:douta	=	16'h	7cf9;
17142	:douta	=	16'h	5b73;
17143	:douta	=	16'h	84d6;
17144	:douta	=	16'h	a598;
17145	:douta	=	16'h	6bf3;
17146	:douta	=	16'h	bdf9;
17147	:douta	=	16'h	94d5;
17148	:douta	=	16'h	94b6;
17149	:douta	=	16'h	42cf;
17150	:douta	=	16'h	4aee;
17151	:douta	=	16'h	0800;
17152	:douta	=	16'h	222e;
17153	:douta	=	16'h	4375;
17154	:douta	=	16'h	32f2;
17155	:douta	=	16'h	4b54;
17156	:douta	=	16'h	4375;
17157	:douta	=	16'h	32d1;
17158	:douta	=	16'h	4333;
17159	:douta	=	16'h	6458;
17160	:douta	=	16'h	5332;
17161	:douta	=	16'h	84f9;
17162	:douta	=	16'h	7cb9;
17163	:douta	=	16'h	63d4;
17164	:douta	=	16'h	4af0;
17165	:douta	=	16'h	73f3;
17166	:douta	=	16'h	7475;
17167	:douta	=	16'h	5b92;
17168	:douta	=	16'h	7c54;
17169	:douta	=	16'h	9cf5;
17170	:douta	=	16'h	73f4;
17171	:douta	=	16'h	b576;
17172	:douta	=	16'h	a536;
17173	:douta	=	16'h	ad35;
17174	:douta	=	16'h	8c94;
17175	:douta	=	16'h	b534;
17176	:douta	=	16'h	eef9;
17177	:douta	=	16'h	bdb5;
17178	:douta	=	16'h	bd74;
17179	:douta	=	16'h	ce36;
17180	:douta	=	16'h	c5f6;
17181	:douta	=	16'h	7b09;
17182	:douta	=	16'h	8369;
17183	:douta	=	16'h	93cb;
17184	:douta	=	16'h	938a;
17185	:douta	=	16'h	ac4c;
17186	:douta	=	16'h	ac4c;
17187	:douta	=	16'h	bc8b;
17188	:douta	=	16'h	bcad;
17189	:douta	=	16'h	b48c;
17190	:douta	=	16'h	c52e;
17191	:douta	=	16'h	d5b0;
17192	:douta	=	16'h	ddf2;
17193	:douta	=	16'h	de12;
17194	:douta	=	16'h	e654;
17195	:douta	=	16'h	ee75;
17196	:douta	=	16'h	e674;
17197	:douta	=	16'h	e634;
17198	:douta	=	16'h	e654;
17199	:douta	=	16'h	e674;
17200	:douta	=	16'h	de13;
17201	:douta	=	16'h	c550;
17202	:douta	=	16'h	bcef;
17203	:douta	=	16'h	c551;
17204	:douta	=	16'h	9c2c;
17205	:douta	=	16'h	72e8;
17206	:douta	=	16'h	b4ae;
17207	:douta	=	16'h	93ec;
17208	:douta	=	16'h	838b;
17209	:douta	=	16'h	9c0d;
17210	:douta	=	16'h	c550;
17211	:douta	=	16'h	de13;
17212	:douta	=	16'h	d5f3;
17213	:douta	=	16'h	d5f3;
17214	:douta	=	16'h	de13;
17215	:douta	=	16'h	ddf3;
17216	:douta	=	16'h	d5b2;
17217	:douta	=	16'h	d591;
17218	:douta	=	16'h	cd71;
17219	:douta	=	16'h	cd50;
17220	:douta	=	16'h	c530;
17221	:douta	=	16'h	acb0;
17222	:douta	=	16'h	9c50;
17223	:douta	=	16'h	8c10;
17224	:douta	=	16'h	83d0;
17225	:douta	=	16'h	6b6f;
17226	:douta	=	16'h	6b6f;
17227	:douta	=	16'h	6b70;
17228	:douta	=	16'h	634f;
17229	:douta	=	16'h	5b50;
17230	:douta	=	16'h	5330;
17231	:douta	=	16'h	42af;
17232	:douta	=	16'h	3a8e;
17233	:douta	=	16'h	324d;
17234	:douta	=	16'h	29eb;
17235	:douta	=	16'h	2988;
17236	:douta	=	16'h	2126;
17237	:douta	=	16'h	0063;
17238	:douta	=	16'h	10e4;
17239	:douta	=	16'h	10e4;
17240	:douta	=	16'h	10c3;
17241	:douta	=	16'h	10e4;
17242	:douta	=	16'h	10c3;
17243	:douta	=	16'h	10a4;
17244	:douta	=	16'h	10a4;
17245	:douta	=	16'h	2967;
17246	:douta	=	16'h	10e5;
17247	:douta	=	16'h	3acf;
17248	:douta	=	16'h	10c6;
17249	:douta	=	16'h	1926;
17250	:douta	=	16'h	08c5;
17251	:douta	=	16'h	2167;
17252	:douta	=	16'h	6b4b;
17253	:douta	=	16'h	6b0a;
17254	:douta	=	16'h	ad11;
17255	:douta	=	16'h	39a6;
17256	:douta	=	16'h	39c6;
17257	:douta	=	16'h	3145;
17258	:douta	=	16'h	5aca;
17259	:douta	=	16'h	4228;
17260	:douta	=	16'h	528a;
17261	:douta	=	16'h	528a;
17262	:douta	=	16'h	8c50;
17263	:douta	=	16'h	942f;
17264	:douta	=	16'h	31c9;
17265	:douta	=	16'h	0064;
17266	:douta	=	16'h	0085;
17267	:douta	=	16'h	1105;
17268	:douta	=	16'h	524a;
17269	:douta	=	16'h	72eb;
17270	:douta	=	16'h	7cd7;
17271	:douta	=	16'h	5bb4;
17272	:douta	=	16'h	9558;
17273	:douta	=	16'h	8d37;
17274	:douta	=	16'h	9559;
17275	:douta	=	16'h	9579;
17276	:douta	=	16'h	adfb;
17277	:douta	=	16'h	9539;
17278	:douta	=	16'h	8d39;
17279	:douta	=	16'h	8d18;
17280	:douta	=	16'h	8d18;
17281	:douta	=	16'h	84f8;
17282	:douta	=	16'h	84d7;
17283	:douta	=	16'h	8d18;
17284	:douta	=	16'h	84f8;
17285	:douta	=	16'h	8d18;
17286	:douta	=	16'h	7cd7;
17287	:douta	=	16'h	957a;
17288	:douta	=	16'h	8d39;
17289	:douta	=	16'h	9559;
17290	:douta	=	16'h	9579;
17291	:douta	=	16'h	9d9a;
17292	:douta	=	16'h	9559;
17293	:douta	=	16'h	8d39;
17294	:douta	=	16'h	9559;
17295	:douta	=	16'h	9559;
17296	:douta	=	16'h	a5db;
17297	:douta	=	16'h	a5db;
17298	:douta	=	16'h	9dbb;
17299	:douta	=	16'h	a5db;
17300	:douta	=	16'h	9dbb;
17301	:douta	=	16'h	959a;
17302	:douta	=	16'h	a5db;
17303	:douta	=	16'h	9d9a;
17304	:douta	=	16'h	6c15;
17305	:douta	=	16'h	7497;
17306	:douta	=	16'h	7cd9;
17307	:douta	=	16'h	9ddc;
17308	:douta	=	16'h	8d3a;
17309	:douta	=	16'h	8d39;
17310	:douta	=	16'h	8d18;
17311	:douta	=	16'h	84f8;
17312	:douta	=	16'h	8518;
17313	:douta	=	16'h	6c14;
17314	:douta	=	16'h	7435;
17315	:douta	=	16'h	838b;
17316	:douta	=	16'h	31a7;
17317	:douta	=	16'h	1905;
17318	:douta	=	16'h	31c9;
17319	:douta	=	16'h	8cf8;
17320	:douta	=	16'h	84f8;
17321	:douta	=	16'h	8d18;
17322	:douta	=	16'h	8d39;
17323	:douta	=	16'h	9d7a;
17324	:douta	=	16'h	a5fb;
17325	:douta	=	16'h	9dba;
17326	:douta	=	16'h	957a;
17327	:douta	=	16'h	8d39;
17328	:douta	=	16'h	955a;
17329	:douta	=	16'h	7cb7;
17330	:douta	=	16'h	8519;
17331	:douta	=	16'h	8d39;
17332	:douta	=	16'h	957b;
17333	:douta	=	16'h	84f8;
17334	:douta	=	16'h	7cb9;
17335	:douta	=	16'h	8539;
17336	:douta	=	16'h	8d5a;
17337	:douta	=	16'h	8d7a;
17338	:douta	=	16'h	8d5a;
17339	:douta	=	16'h	957a;
17340	:douta	=	16'h	957a;
17341	:douta	=	16'h	9559;
17342	:douta	=	16'h	6bf4;
17343	:douta	=	16'h	63d3;
17344	:douta	=	16'h	7435;
17345	:douta	=	16'h	9539;
17346	:douta	=	16'h	9559;
17347	:douta	=	16'h	8518;
17348	:douta	=	16'h	7c55;
17349	:douta	=	16'h	6c15;
17350	:douta	=	16'h	2905;
17351	:douta	=	16'h	2146;
17352	:douta	=	16'h	10c5;
17353	:douta	=	16'h	1905;
17354	:douta	=	16'h	5c15;
17355	:douta	=	16'h	5c16;
17356	:douta	=	16'h	7d5a;
17357	:douta	=	16'h	751a;
17358	:douta	=	16'h	74d9;
17359	:douta	=	16'h	6cb9;
17360	:douta	=	16'h	6c79;
17361	:douta	=	16'h	6cb8;
17362	:douta	=	16'h	6c98;
17363	:douta	=	16'h	74da;
17364	:douta	=	16'h	6cb9;
17365	:douta	=	16'h	6cb9;
17366	:douta	=	16'h	6c98;
17367	:douta	=	16'h	74d9;
17368	:douta	=	16'h	74d9;
17369	:douta	=	16'h	7cf9;
17370	:douta	=	16'h	74d9;
17371	:douta	=	16'h	74b9;
17372	:douta	=	16'h	6c56;
17373	:douta	=	16'h	7457;
17374	:douta	=	16'h	74d9;
17375	:douta	=	16'h	7d1a;
17376	:douta	=	16'h	7498;
17377	:douta	=	16'h	5bd5;
17378	:douta	=	16'h	63f6;
17379	:douta	=	16'h	8d5b;
17380	:douta	=	16'h	6c77;
17381	:douta	=	16'h	7498;
17382	:douta	=	16'h	7cd9;
17383	:douta	=	16'h	851a;
17384	:douta	=	16'h	7478;
17385	:douta	=	16'h	853a;
17386	:douta	=	16'h	7cf9;
17387	:douta	=	16'h	853b;
17388	:douta	=	16'h	7d1a;
17389	:douta	=	16'h	855a;
17390	:douta	=	16'h	853a;
17391	:douta	=	16'h	8519;
17392	:douta	=	16'h	7cfa;
17393	:douta	=	16'h	853a;
17394	:douta	=	16'h	853a;
17395	:douta	=	16'h	851a;
17396	:douta	=	16'h	853a;
17397	:douta	=	16'h	6c77;
17398	:douta	=	16'h	29cb;
17399	:douta	=	16'h	defd;
17400	:douta	=	16'h	6c15;
17401	:douta	=	16'h	8496;
17402	:douta	=	16'h	8cb6;
17403	:douta	=	16'h	a558;
17404	:douta	=	16'h	42ae;
17405	:douta	=	16'h	8cd4;
17406	:douta	=	16'h	73b0;
17407	:douta	=	16'h	3a2a;
17408	:douta	=	16'h	3ad1;
17409	:douta	=	16'h	2a4f;
17410	:douta	=	16'h	2a4f;
17411	:douta	=	16'h	4374;
17412	:douta	=	16'h	32b1;
17413	:douta	=	16'h	3312;
17414	:douta	=	16'h	4374;
17415	:douta	=	16'h	53d5;
17416	:douta	=	16'h	3290;
17417	:douta	=	16'h	6c36;
17418	:douta	=	16'h	6415;
17419	:douta	=	16'h	5373;
17420	:douta	=	16'h	63b4;
17421	:douta	=	16'h	7435;
17422	:douta	=	16'h	9559;
17423	:douta	=	16'h	7414;
17424	:douta	=	16'h	73f3;
17425	:douta	=	16'h	7c33;
17426	:douta	=	16'h	6bd2;
17427	:douta	=	16'h	ad36;
17428	:douta	=	16'h	a537;
17429	:douta	=	16'h	eefb;
17430	:douta	=	16'h	9d15;
17431	:douta	=	16'h	ad34;
17432	:douta	=	16'h	bd94;
17433	:douta	=	16'h	b594;
17434	:douta	=	16'h	bd95;
17435	:douta	=	16'h	e6f9;
17436	:douta	=	16'h	9cd3;
17437	:douta	=	16'h	8329;
17438	:douta	=	16'h	93cb;
17439	:douta	=	16'h	93aa;
17440	:douta	=	16'h	93aa;
17441	:douta	=	16'h	b44b;
17442	:douta	=	16'h	b48c;
17443	:douta	=	16'h	c4cd;
17444	:douta	=	16'h	bccd;
17445	:douta	=	16'h	c4ed;
17446	:douta	=	16'h	cd6f;
17447	:douta	=	16'h	ddd1;
17448	:douta	=	16'h	de33;
17449	:douta	=	16'h	de33;
17450	:douta	=	16'h	ee75;
17451	:douta	=	16'h	e675;
17452	:douta	=	16'h	ee96;
17453	:douta	=	16'h	de13;
17454	:douta	=	16'h	e633;
17455	:douta	=	16'h	de34;
17456	:douta	=	16'h	ddd2;
17457	:douta	=	16'h	cd91;
17458	:douta	=	16'h	bcef;
17459	:douta	=	16'h	c50f;
17460	:douta	=	16'h	b4ae;
17461	:douta	=	16'h	72e7;
17462	:douta	=	16'h	b4ce;
17463	:douta	=	16'h	a42d;
17464	:douta	=	16'h	838b;
17465	:douta	=	16'h	8bab;
17466	:douta	=	16'h	a48c;
17467	:douta	=	16'h	cd91;
17468	:douta	=	16'h	d5d2;
17469	:douta	=	16'h	de34;
17470	:douta	=	16'h	de14;
17471	:douta	=	16'h	de13;
17472	:douta	=	16'h	d5b2;
17473	:douta	=	16'h	d5b2;
17474	:douta	=	16'h	cd71;
17475	:douta	=	16'h	cd71;
17476	:douta	=	16'h	c551;
17477	:douta	=	16'h	b4d0;
17478	:douta	=	16'h	9c50;
17479	:douta	=	16'h	9410;
17480	:douta	=	16'h	83cf;
17481	:douta	=	16'h	73b0;
17482	:douta	=	16'h	6b6f;
17483	:douta	=	16'h	634f;
17484	:douta	=	16'h	5b2f;
17485	:douta	=	16'h	5b0f;
17486	:douta	=	16'h	52ef;
17487	:douta	=	16'h	42ef;
17488	:douta	=	16'h	42ae;
17489	:douta	=	16'h	3a6d;
17490	:douta	=	16'h	3a6d;
17491	:douta	=	16'h	2189;
17492	:douta	=	16'h	6b4e;
17493	:douta	=	16'h	18e5;
17494	:douta	=	16'h	10e4;
17495	:douta	=	16'h	0883;
17496	:douta	=	16'h	10c4;
17497	:douta	=	16'h	10c4;
17498	:douta	=	16'h	10e4;
17499	:douta	=	16'h	10c4;
17500	:douta	=	16'h	10c5;
17501	:douta	=	16'h	10e5;
17502	:douta	=	16'h	2146;
17503	:douta	=	16'h	0000;
17504	:douta	=	16'h	2988;
17505	:douta	=	16'h	2189;
17506	:douta	=	16'h	1947;
17507	:douta	=	16'h	10e5;
17508	:douta	=	16'h	10c5;
17509	:douta	=	16'h	18e4;
17510	:douta	=	16'h	738c;
17511	:douta	=	16'h	62ea;
17512	:douta	=	16'h	5289;
17513	:douta	=	16'h	736c;
17514	:douta	=	16'h	528a;
17515	:douta	=	16'h	10c4;
17516	:douta	=	16'h	0043;
17517	:douta	=	16'h	0000;
17518	:douta	=	16'h	6b8e;
17519	:douta	=	16'h	b551;
17520	:douta	=	16'h	944f;
17521	:douta	=	16'h	8c0f;
17522	:douta	=	16'h	6b4d;
17523	:douta	=	16'h	29c9;
17524	:douta	=	16'h	0884;
17525	:douta	=	16'h	628a;
17526	:douta	=	16'h	9539;
17527	:douta	=	16'h	7cf7;
17528	:douta	=	16'h	7455;
17529	:douta	=	16'h	7476;
17530	:douta	=	16'h	7cb7;
17531	:douta	=	16'h	7c96;
17532	:douta	=	16'h	7cb7;
17533	:douta	=	16'h	957a;
17534	:douta	=	16'h	9559;
17535	:douta	=	16'h	9579;
17536	:douta	=	16'h	9579;
17537	:douta	=	16'h	9d9a;
17538	:douta	=	16'h	8d18;
17539	:douta	=	16'h	84d7;
17540	:douta	=	16'h	9d9a;
17541	:douta	=	16'h	9579;
17542	:douta	=	16'h	8518;
17543	:douta	=	16'h	8d38;
17544	:douta	=	16'h	7cb7;
17545	:douta	=	16'h	8d18;
17546	:douta	=	16'h	8d18;
17547	:douta	=	16'h	9599;
17548	:douta	=	16'h	84d7;
17549	:douta	=	16'h	9d9a;
17550	:douta	=	16'h	8d18;
17551	:douta	=	16'h	9d9a;
17552	:douta	=	16'h	9d9a;
17553	:douta	=	16'h	a5da;
17554	:douta	=	16'h	a5ba;
17555	:douta	=	16'h	a5ba;
17556	:douta	=	16'h	a5db;
17557	:douta	=	16'h	adfb;
17558	:douta	=	16'h	8d5a;
17559	:douta	=	16'h	ae3c;
17560	:douta	=	16'h	b67d;
17561	:douta	=	16'h	9d9a;
17562	:douta	=	16'h	8d39;
17563	:douta	=	16'h	7cd9;
17564	:douta	=	16'h	7cf9;
17565	:douta	=	16'h	95bb;
17566	:douta	=	16'h	8d39;
17567	:douta	=	16'h	84d8;
17568	:douta	=	16'h	84f8;
17569	:douta	=	16'h	8cf9;
17570	:douta	=	16'h	84d7;
17571	:douta	=	16'h	93ed;
17572	:douta	=	16'h	4a08;
17573	:douta	=	16'h	1905;
17574	:douta	=	16'h	10a5;
17575	:douta	=	16'h	6c15;
17576	:douta	=	16'h	8d19;
17577	:douta	=	16'h	8cd8;
17578	:douta	=	16'h	8d39;
17579	:douta	=	16'h	8d39;
17580	:douta	=	16'h	84b7;
17581	:douta	=	16'h	a5db;
17582	:douta	=	16'h	a5ba;
17583	:douta	=	16'h	9d9a;
17584	:douta	=	16'h	9dbb;
17585	:douta	=	16'h	a5fb;
17586	:douta	=	16'h	8d5a;
17587	:douta	=	16'h	8d59;
17588	:douta	=	16'h	8519;
17589	:douta	=	16'h	957b;
17590	:douta	=	16'h	955a;
17591	:douta	=	16'h	7456;
17592	:douta	=	16'h	6c15;
17593	:douta	=	16'h	84f8;
17594	:douta	=	16'h	9559;
17595	:douta	=	16'h	9dbb;
17596	:douta	=	16'h	8d39;
17597	:douta	=	16'h	8d18;
17598	:douta	=	16'h	8cd8;
17599	:douta	=	16'h	7c55;
17600	:douta	=	16'h	7435;
17601	:douta	=	16'h	7414;
17602	:douta	=	16'h	7c75;
17603	:douta	=	16'h	84f8;
17604	:douta	=	16'h	8d18;
17605	:douta	=	16'h	8519;
17606	:douta	=	16'h	2105;
17607	:douta	=	16'h	2126;
17608	:douta	=	16'h	10e5;
17609	:douta	=	16'h	10c5;
17610	:douta	=	16'h	5c17;
17611	:douta	=	16'h	6437;
17612	:douta	=	16'h	6437;
17613	:douta	=	16'h	6458;
17614	:douta	=	16'h	6458;
17615	:douta	=	16'h	6cba;
17616	:douta	=	16'h	74fa;
17617	:douta	=	16'h	6cd9;
17618	:douta	=	16'h	74da;
17619	:douta	=	16'h	751a;
17620	:douta	=	16'h	74fa;
17621	:douta	=	16'h	74d9;
17622	:douta	=	16'h	855b;
17623	:douta	=	16'h	74b8;
17624	:douta	=	16'h	7498;
17625	:douta	=	16'h	855a;
17626	:douta	=	16'h	74b8;
17627	:douta	=	16'h	7498;
17628	:douta	=	16'h	7cf9;
17629	:douta	=	16'h	74b8;
17630	:douta	=	16'h	74b8;
17631	:douta	=	16'h	7cd9;
17632	:douta	=	16'h	7498;
17633	:douta	=	16'h	7cf9;
17634	:douta	=	16'h	7498;
17635	:douta	=	16'h	7cd8;
17636	:douta	=	16'h	8d9b;
17637	:douta	=	16'h	853a;
17638	:douta	=	16'h	7478;
17639	:douta	=	16'h	7cd9;
17640	:douta	=	16'h	7cd9;
17641	:douta	=	16'h	74d9;
17642	:douta	=	16'h	7cd9;
17643	:douta	=	16'h	8d5b;
17644	:douta	=	16'h	7d1a;
17645	:douta	=	16'h	74d9;
17646	:douta	=	16'h	7d3a;
17647	:douta	=	16'h	7cda;
17648	:douta	=	16'h	8d3a;
17649	:douta	=	16'h	7cd9;
17650	:douta	=	16'h	8d7b;
17651	:douta	=	16'h	855a;
17652	:douta	=	16'h	7d3a;
17653	:douta	=	16'h	6415;
17654	:douta	=	16'h	31a9;
17655	:douta	=	16'h	b61a;
17656	:douta	=	16'h	5bb3;
17657	:douta	=	16'h	8cb6;
17658	:douta	=	16'h	d69b;
17659	:douta	=	16'h	9d37;
17660	:douta	=	16'h	532f;
17661	:douta	=	16'h	5331;
17662	:douta	=	16'h	39e8;
17663	:douta	=	16'h	4aad;
17664	:douta	=	16'h	2a0c;
17665	:douta	=	16'h	2a6f;
17666	:douta	=	16'h	2a90;
17667	:douta	=	16'h	3b33;
17668	:douta	=	16'h	64da;
17669	:douta	=	16'h	2ab0;
17670	:douta	=	16'h	32b1;
17671	:douta	=	16'h	4b75;
17672	:douta	=	16'h	3ad1;
17673	:douta	=	16'h	63d4;
17674	:douta	=	16'h	5bb4;
17675	:douta	=	16'h	7477;
17676	:douta	=	16'h	6c35;
17677	:douta	=	16'h	6bf3;
17678	:douta	=	16'h	63f4;
17679	:douta	=	16'h	5b72;
17680	:douta	=	16'h	73f3;
17681	:douta	=	16'h	8c74;
17682	:douta	=	16'h	94d5;
17683	:douta	=	16'h	b5b7;
17684	:douta	=	16'h	b597;
17685	:douta	=	16'h	a515;
17686	:douta	=	16'h	94b4;
17687	:douta	=	16'h	9cb3;
17688	:douta	=	16'h	b574;
17689	:douta	=	16'h	bdb6;
17690	:douta	=	16'h	c5f6;
17691	:douta	=	16'h	bdb6;
17692	:douta	=	16'h	72a8;
17693	:douta	=	16'h	8b8a;
17694	:douta	=	16'h	a42a;
17695	:douta	=	16'h	93ca;
17696	:douta	=	16'h	ac4c;
17697	:douta	=	16'h	b46c;
17698	:douta	=	16'h	c4cd;
17699	:douta	=	16'h	cd0d;
17700	:douta	=	16'h	cd4f;
17701	:douta	=	16'h	cd2e;
17702	:douta	=	16'h	ddd1;
17703	:douta	=	16'h	ddd1;
17704	:douta	=	16'h	e675;
17705	:douta	=	16'h	ee75;
17706	:douta	=	16'h	ee75;
17707	:douta	=	16'h	ee95;
17708	:douta	=	16'h	ee75;
17709	:douta	=	16'h	e634;
17710	:douta	=	16'h	c52f;
17711	:douta	=	16'h	ddd1;
17712	:douta	=	16'h	d5b1;
17713	:douta	=	16'h	b4ad;
17714	:douta	=	16'h	a44d;
17715	:douta	=	16'h	9c0b;
17716	:douta	=	16'h	8327;
17717	:douta	=	16'h	9c2c;
17718	:douta	=	16'h	ac8e;
17719	:douta	=	16'h	bcef;
17720	:douta	=	16'h	b4ae;
17721	:douta	=	16'h	b4ae;
17722	:douta	=	16'h	b4ae;
17723	:douta	=	16'h	cd70;
17724	:douta	=	16'h	d5d2;
17725	:douta	=	16'h	de13;
17726	:douta	=	16'h	de34;
17727	:douta	=	16'h	de13;
17728	:douta	=	16'h	d5b1;
17729	:douta	=	16'h	d591;
17730	:douta	=	16'h	d5b2;
17731	:douta	=	16'h	cd71;
17732	:douta	=	16'h	c531;
17733	:douta	=	16'h	bd11;
17734	:douta	=	16'h	a491;
17735	:douta	=	16'h	9430;
17736	:douta	=	16'h	8c10;
17737	:douta	=	16'h	73b0;
17738	:douta	=	16'h	7390;
17739	:douta	=	16'h	7390;
17740	:douta	=	16'h	6b91;
17741	:douta	=	16'h	6b71;
17742	:douta	=	16'h	5b30;
17743	:douta	=	16'h	4aef;
17744	:douta	=	16'h	4acf;
17745	:douta	=	16'h	3a4d;
17746	:douta	=	16'h	322c;
17747	:douta	=	16'h	3a0b;
17748	:douta	=	16'h	1127;
17749	:douta	=	16'h	528d;
17750	:douta	=	16'h	18e5;
17751	:douta	=	16'h	0883;
17752	:douta	=	16'h	10a4;
17753	:douta	=	16'h	10c4;
17754	:douta	=	16'h	10c4;
17755	:douta	=	16'h	10e4;
17756	:douta	=	16'h	10e4;
17757	:douta	=	16'h	10a4;
17758	:douta	=	16'h	10e4;
17759	:douta	=	16'h	1906;
17760	:douta	=	16'h	0063;
17761	:douta	=	16'h	0884;
17762	:douta	=	16'h	21a9;
17763	:douta	=	16'h	1947;
17764	:douta	=	16'h	1106;
17765	:douta	=	16'h	62ea;
17766	:douta	=	16'h	7bcd;
17767	:douta	=	16'h	62e9;
17768	:douta	=	16'h	2126;
17769	:douta	=	16'h	732b;
17770	:douta	=	16'h	0042;
17771	:douta	=	16'h	5248;
17772	:douta	=	16'h	18e5;
17773	:douta	=	16'h	2966;
17774	:douta	=	16'h	7bcc;
17775	:douta	=	16'h	6b6e;
17776	:douta	=	16'h	31a8;
17777	:douta	=	16'h	3a29;
17778	:douta	=	16'h	4aab;
17779	:douta	=	16'h	632e;
17780	:douta	=	16'h	7b8d;
17781	:douta	=	16'h	b532;
17782	:douta	=	16'h	84d6;
17783	:douta	=	16'h	9559;
17784	:douta	=	16'h	6c14;
17785	:douta	=	16'h	7455;
17786	:douta	=	16'h	7455;
17787	:douta	=	16'h	957a;
17788	:douta	=	16'h	b63c;
17789	:douta	=	16'h	8d18;
17790	:douta	=	16'h	6c36;
17791	:douta	=	16'h	63f4;
17792	:douta	=	16'h	8d18;
17793	:douta	=	16'h	84f7;
17794	:douta	=	16'h	9d9a;
17795	:douta	=	16'h	9d7a;
17796	:douta	=	16'h	9539;
17797	:douta	=	16'h	9599;
17798	:douta	=	16'h	9579;
17799	:douta	=	16'h	8518;
17800	:douta	=	16'h	9579;
17801	:douta	=	16'h	8d39;
17802	:douta	=	16'h	957a;
17803	:douta	=	16'h	9d9a;
17804	:douta	=	16'h	957a;
17805	:douta	=	16'h	8d39;
17806	:douta	=	16'h	957a;
17807	:douta	=	16'h	9d9a;
17808	:douta	=	16'h	9d9a;
17809	:douta	=	16'h	9d9a;
17810	:douta	=	16'h	8d39;
17811	:douta	=	16'h	959a;
17812	:douta	=	16'h	9dba;
17813	:douta	=	16'h	9dbb;
17814	:douta	=	16'h	a5db;
17815	:douta	=	16'h	957a;
17816	:douta	=	16'h	957a;
17817	:douta	=	16'h	9dbb;
17818	:douta	=	16'h	95bb;
17819	:douta	=	16'h	9ddb;
17820	:douta	=	16'h	a5fb;
17821	:douta	=	16'h	9d9a;
17822	:douta	=	16'h	7cb8;
17823	:douta	=	16'h	6c36;
17824	:douta	=	16'h	8d19;
17825	:douta	=	16'h	957a;
17826	:douta	=	16'h	7c98;
17827	:douta	=	16'h	a46f;
17828	:douta	=	16'h	6b0a;
17829	:douta	=	16'h	10e5;
17830	:douta	=	16'h	0862;
17831	:douta	=	16'h	322c;
17832	:douta	=	16'h	84d8;
17833	:douta	=	16'h	84f8;
17834	:douta	=	16'h	9559;
17835	:douta	=	16'h	9539;
17836	:douta	=	16'h	9dba;
17837	:douta	=	16'h	9d7a;
17838	:douta	=	16'h	9d79;
17839	:douta	=	16'h	9518;
17840	:douta	=	16'h	7c95;
17841	:douta	=	16'h	9559;
17842	:douta	=	16'h	9559;
17843	:douta	=	16'h	957a;
17844	:douta	=	16'h	a5dc;
17845	:douta	=	16'h	9dfc;
17846	:douta	=	16'h	9dbb;
17847	:douta	=	16'h	9d9a;
17848	:douta	=	16'h	84f8;
17849	:douta	=	16'h	84b6;
17850	:douta	=	16'h	8475;
17851	:douta	=	16'h	7c13;
17852	:douta	=	16'h	7c33;
17853	:douta	=	16'h	8d17;
17854	:douta	=	16'h	84d7;
17855	:douta	=	16'h	84d7;
17856	:douta	=	16'h	84b7;
17857	:douta	=	16'h	84d7;
17858	:douta	=	16'h	84f8;
17859	:douta	=	16'h	7456;
17860	:douta	=	16'h	6c35;
17861	:douta	=	16'h	6392;
17862	:douta	=	16'h	2146;
17863	:douta	=	16'h	1925;
17864	:douta	=	16'h	10e5;
17865	:douta	=	16'h	2106;
17866	:douta	=	16'h	53d6;
17867	:douta	=	16'h	4313;
17868	:douta	=	16'h	5bf6;
17869	:douta	=	16'h	5c78;
17870	:douta	=	16'h	4bf6;
17871	:douta	=	16'h	6458;
17872	:douta	=	16'h	6457;
17873	:douta	=	16'h	5bf6;
17874	:douta	=	16'h	6c98;
17875	:douta	=	16'h	74d9;
17876	:douta	=	16'h	74d9;
17877	:douta	=	16'h	74f9;
17878	:douta	=	16'h	7d19;
17879	:douta	=	16'h	7cf9;
17880	:douta	=	16'h	6c78;
17881	:douta	=	16'h	6c77;
17882	:douta	=	16'h	74b8;
17883	:douta	=	16'h	7cf9;
17884	:douta	=	16'h	853a;
17885	:douta	=	16'h	7d19;
17886	:douta	=	16'h	851a;
17887	:douta	=	16'h	7cf9;
17888	:douta	=	16'h	7cf9;
17889	:douta	=	16'h	74b8;
17890	:douta	=	16'h	7cd9;
17891	:douta	=	16'h	851a;
17892	:douta	=	16'h	7497;
17893	:douta	=	16'h	6436;
17894	:douta	=	16'h	8519;
17895	:douta	=	16'h	8d9b;
17896	:douta	=	16'h	7cf9;
17897	:douta	=	16'h	6c77;
17898	:douta	=	16'h	853a;
17899	:douta	=	16'h	8d5b;
17900	:douta	=	16'h	7d1a;
17901	:douta	=	16'h	8d7b;
17902	:douta	=	16'h	8d7a;
17903	:douta	=	16'h	7d1a;
17904	:douta	=	16'h	8d7b;
17905	:douta	=	16'h	8d7b;
17906	:douta	=	16'h	851a;
17907	:douta	=	16'h	7cf9;
17908	:douta	=	16'h	7cd9;
17909	:douta	=	16'h	428d;
17910	:douta	=	16'h	73d0;
17911	:douta	=	16'h	63b1;
17912	:douta	=	16'h	8cb6;
17913	:douta	=	16'h	b5d9;
17914	:douta	=	16'h	328e;
17915	:douta	=	16'h	5b71;
17916	:douta	=	16'h	7c33;
17917	:douta	=	16'h	5aee;
17918	:douta	=	16'h	0000;
17919	:douta	=	16'h	a557;
17920	:douta	=	16'h	328f;
17921	:douta	=	16'h	2a6f;
17922	:douta	=	16'h	2a4f;
17923	:douta	=	16'h	3af3;
17924	:douta	=	16'h	3b33;
17925	:douta	=	16'h	2250;
17926	:douta	=	16'h	4374;
17927	:douta	=	16'h	6457;
17928	:douta	=	16'h	4312;
17929	:douta	=	16'h	5b93;
17930	:douta	=	16'h	5373;
17931	:douta	=	16'h	5bf5;
17932	:douta	=	16'h	6415;
17933	:douta	=	16'h	4acf;
17934	:douta	=	16'h	84d7;
17935	:douta	=	16'h	7c96;
17936	:douta	=	16'h	8c94;
17937	:douta	=	16'h	73f3;
17938	:douta	=	16'h	a536;
17939	:douta	=	16'h	9cb4;
17940	:douta	=	16'h	bdd7;
17941	:douta	=	16'h	bdd7;
17942	:douta	=	16'h	b5b6;
17943	:douta	=	16'h	ad34;
17944	:douta	=	16'h	8c31;
17945	:douta	=	16'h	a4f3;
17946	:douta	=	16'h	ad76;
17947	:douta	=	16'h	ad13;
17948	:douta	=	16'h	832a;
17949	:douta	=	16'h	9beb;
17950	:douta	=	16'h	ac4b;
17951	:douta	=	16'h	a40b;
17952	:douta	=	16'h	ac4c;
17953	:douta	=	16'h	b46b;
17954	:douta	=	16'h	cd4e;
17955	:douta	=	16'h	cd0d;
17956	:douta	=	16'h	d58f;
17957	:douta	=	16'h	cd6e;
17958	:douta	=	16'h	de13;
17959	:douta	=	16'h	cd90;
17960	:douta	=	16'h	e654;
17961	:douta	=	16'h	eeb7;
17962	:douta	=	16'h	eeb6;
17963	:douta	=	16'h	e675;
17964	:douta	=	16'h	e654;
17965	:douta	=	16'h	e654;
17966	:douta	=	16'h	ac6c;
17967	:douta	=	16'h	b4ae;
17968	:douta	=	16'h	ddd1;
17969	:douta	=	16'h	ac4c;
17970	:douta	=	16'h	a42d;
17971	:douta	=	16'h	72a6;
17972	:douta	=	16'h	9c2b;
17973	:douta	=	16'h	9c2d;
17974	:douta	=	16'h	ac6d;
17975	:douta	=	16'h	ac8d;
17976	:douta	=	16'h	c50f;
17977	:douta	=	16'h	bd0f;
17978	:douta	=	16'h	cd71;
17979	:douta	=	16'h	d5b2;
17980	:douta	=	16'h	ddf3;
17981	:douta	=	16'h	de14;
17982	:douta	=	16'h	de34;
17983	:douta	=	16'h	de13;
17984	:douta	=	16'h	d5b2;
17985	:douta	=	16'h	d5b2;
17986	:douta	=	16'h	d591;
17987	:douta	=	16'h	d591;
17988	:douta	=	16'h	c530;
17989	:douta	=	16'h	bd11;
17990	:douta	=	16'h	acb1;
17991	:douta	=	16'h	9c51;
17992	:douta	=	16'h	9430;
17993	:douta	=	16'h	83d0;
17994	:douta	=	16'h	7bd1;
17995	:douta	=	16'h	73b1;
17996	:douta	=	16'h	6b70;
17997	:douta	=	16'h	6b71;
17998	:douta	=	16'h	6371;
17999	:douta	=	16'h	5b50;
18000	:douta	=	16'h	530f;
18001	:douta	=	16'h	4aae;
18002	:douta	=	16'h	428d;
18003	:douta	=	16'h	3a2c;
18004	:douta	=	16'h	320c;
18005	:douta	=	16'h	2169;
18006	:douta	=	16'h	6b2c;
18007	:douta	=	16'h	1906;
18008	:douta	=	16'h	18e4;
18009	:douta	=	16'h	10c4;
18010	:douta	=	16'h	10c4;
18011	:douta	=	16'h	10c3;
18012	:douta	=	16'h	10e4;
18013	:douta	=	16'h	10a3;
18014	:douta	=	16'h	10c4;
18015	:douta	=	16'h	10e5;
18016	:douta	=	16'h	1906;
18017	:douta	=	16'h	0863;
18018	:douta	=	16'h	2167;
18019	:douta	=	16'h	2189;
18020	:douta	=	16'h	1946;
18021	:douta	=	16'h	08a5;
18022	:douta	=	16'h	0884;
18023	:douta	=	16'h	3a07;
18024	:douta	=	16'h	08a4;
18025	:douta	=	16'h	c592;
18026	:douta	=	16'h	2947;
18027	:douta	=	16'h	944f;
18028	:douta	=	16'h	2124;
18029	:douta	=	16'h	5249;
18030	:douta	=	16'h	18a3;
18031	:douta	=	16'h	630c;
18032	:douta	=	16'h	2146;
18033	:douta	=	16'h	ad12;
18034	:douta	=	16'h	8c30;
18035	:douta	=	16'h	52cc;
18036	:douta	=	16'h	83ed;
18037	:douta	=	16'h	7b8d;
18038	:douta	=	16'h	6bd2;
18039	:douta	=	16'h	ae3c;
18040	:douta	=	16'h	a5db;
18041	:douta	=	16'h	84b6;
18042	:douta	=	16'h	7415;
18043	:douta	=	16'h	7cb6;
18044	:douta	=	16'h	8cf8;
18045	:douta	=	16'h	a5fb;
18046	:douta	=	16'h	a5db;
18047	:douta	=	16'h	7cb7;
18048	:douta	=	16'h	9559;
18049	:douta	=	16'h	8d39;
18050	:douta	=	16'h	84f8;
18051	:douta	=	16'h	b65b;
18052	:douta	=	16'h	b63b;
18053	:douta	=	16'h	a5da;
18054	:douta	=	16'h	a5ba;
18055	:douta	=	16'h	8d59;
18056	:douta	=	16'h	9559;
18057	:douta	=	16'h	a5ba;
18058	:douta	=	16'h	8d39;
18059	:douta	=	16'h	8d18;
18060	:douta	=	16'h	9559;
18061	:douta	=	16'h	a5ba;
18062	:douta	=	16'h	a5ba;
18063	:douta	=	16'h	957a;
18064	:douta	=	16'h	9559;
18065	:douta	=	16'h	a5ba;
18066	:douta	=	16'h	9d9a;
18067	:douta	=	16'h	957a;
18068	:douta	=	16'h	9559;
18069	:douta	=	16'h	9559;
18070	:douta	=	16'h	9dba;
18071	:douta	=	16'h	a5ba;
18072	:douta	=	16'h	9dba;
18073	:douta	=	16'h	957a;
18074	:douta	=	16'h	9dba;
18075	:douta	=	16'h	a5db;
18076	:douta	=	16'h	8d5a;
18077	:douta	=	16'h	9dbb;
18078	:douta	=	16'h	adfb;
18079	:douta	=	16'h	8d39;
18080	:douta	=	16'h	7c77;
18081	:douta	=	16'h	8d39;
18082	:douta	=	16'h	84d8;
18083	:douta	=	16'h	a4f2;
18084	:douta	=	16'h	8b8b;
18085	:douta	=	16'h	10e5;
18086	:douta	=	16'h	10c4;
18087	:douta	=	16'h	2167;
18088	:douta	=	16'h	7cb8;
18089	:douta	=	16'h	6415;
18090	:douta	=	16'h	9559;
18091	:douta	=	16'h	a5db;
18092	:douta	=	16'h	84f8;
18093	:douta	=	16'h	9d79;
18094	:douta	=	16'h	a5ba;
18095	:douta	=	16'h	9d58;
18096	:douta	=	16'h	9d79;
18097	:douta	=	16'h	84d6;
18098	:douta	=	16'h	84b6;
18099	:douta	=	16'h	8d39;
18100	:douta	=	16'h	9dbb;
18101	:douta	=	16'h	9dbb;
18102	:douta	=	16'h	a61c;
18103	:douta	=	16'h	9d9a;
18104	:douta	=	16'h	9518;
18105	:douta	=	16'h	8495;
18106	:douta	=	16'h	8495;
18107	:douta	=	16'h	8cb4;
18108	:douta	=	16'h	7c12;
18109	:douta	=	16'h	8495;
18110	:douta	=	16'h	8cd7;
18111	:douta	=	16'h	84b7;
18112	:douta	=	16'h	8cf8;
18113	:douta	=	16'h	8d19;
18114	:douta	=	16'h	84d8;
18115	:douta	=	16'h	84d7;
18116	:douta	=	16'h	7476;
18117	:douta	=	16'h	4a8d;
18118	:douta	=	16'h	2146;
18119	:douta	=	16'h	1905;
18120	:douta	=	16'h	18e5;
18121	:douta	=	16'h	2107;
18122	:douta	=	16'h	8ddf;
18123	:douta	=	16'h	4333;
18124	:douta	=	16'h	3b12;
18125	:douta	=	16'h	5417;
18126	:douta	=	16'h	6499;
18127	:douta	=	16'h	5c58;
18128	:douta	=	16'h	6cda;
18129	:douta	=	16'h	5c37;
18130	:douta	=	16'h	4b94;
18131	:douta	=	16'h	5394;
18132	:douta	=	16'h	5c16;
18133	:douta	=	16'h	7d3a;
18134	:douta	=	16'h	7519;
18135	:douta	=	16'h	74d9;
18136	:douta	=	16'h	7cd9;
18137	:douta	=	16'h	7498;
18138	:douta	=	16'h	7d19;
18139	:douta	=	16'h	7498;
18140	:douta	=	16'h	851a;
18141	:douta	=	16'h	84f9;
18142	:douta	=	16'h	851a;
18143	:douta	=	16'h	853a;
18144	:douta	=	16'h	7cd9;
18145	:douta	=	16'h	7cd9;
18146	:douta	=	16'h	7cd9;
18147	:douta	=	16'h	7cd9;
18148	:douta	=	16'h	8d5a;
18149	:douta	=	16'h	8d5b;
18150	:douta	=	16'h	7498;
18151	:douta	=	16'h	7498;
18152	:douta	=	16'h	8d5a;
18153	:douta	=	16'h	7d19;
18154	:douta	=	16'h	6c57;
18155	:douta	=	16'h	853a;
18156	:douta	=	16'h	853a;
18157	:douta	=	16'h	7cf9;
18158	:douta	=	16'h	959b;
18159	:douta	=	16'h	853a;
18160	:douta	=	16'h	8519;
18161	:douta	=	16'h	8d5a;
18162	:douta	=	16'h	8d7b;
18163	:douta	=	16'h	7cf9;
18164	:douta	=	16'h	7cf9;
18165	:douta	=	16'h	3a0a;
18166	:douta	=	16'h	52ac;
18167	:douta	=	16'h	8434;
18168	:douta	=	16'h	adb9;
18169	:douta	=	16'h	be3a;
18170	:douta	=	16'h	7c33;
18171	:douta	=	16'h	8495;
18172	:douta	=	16'h	3a8f;
18173	:douta	=	16'h	41c8;
18174	:douta	=	16'h	0041;
18175	:douta	=	16'h	a577;
18176	:douta	=	16'h	2106;
18177	:douta	=	16'h	32f2;
18178	:douta	=	16'h	2a90;
18179	:douta	=	16'h	3af2;
18180	:douta	=	16'h	751c;
18181	:douta	=	16'h	5416;
18182	:douta	=	16'h	2a4f;
18183	:douta	=	16'h	3b12;
18184	:douta	=	16'h	53b4;
18185	:douta	=	16'h	63f5;
18186	:douta	=	16'h	63f5;
18187	:douta	=	16'h	5bb4;
18188	:douta	=	16'h	6c35;
18189	:douta	=	16'h	6392;
18190	:douta	=	16'h	7cb7;
18191	:douta	=	16'h	6392;
18192	:douta	=	16'h	4ace;
18193	:douta	=	16'h	7bf2;
18194	:douta	=	16'h	8433;
18195	:douta	=	16'h	a536;
18196	:douta	=	16'h	bdb7;
18197	:douta	=	16'h	c618;
18198	:douta	=	16'h	c618;
18199	:douta	=	16'h	8411;
18200	:douta	=	16'h	9493;
18201	:douta	=	16'h	c5f6;
18202	:douta	=	16'h	834b;
18203	:douta	=	16'h	834a;
18204	:douta	=	16'h	8b8b;
18205	:douta	=	16'h	b44b;
18206	:douta	=	16'h	ac2a;
18207	:douta	=	16'h	b4ac;
18208	:douta	=	16'h	c4ed;
18209	:douta	=	16'h	c4ed;
18210	:douta	=	16'h	d58f;
18211	:douta	=	16'h	d5b0;
18212	:douta	=	16'h	ddd1;
18213	:douta	=	16'h	d5b0;
18214	:douta	=	16'h	de13;
18215	:douta	=	16'h	ee75;
18216	:douta	=	16'h	de13;
18217	:douta	=	16'h	de13;
18218	:douta	=	16'h	ee95;
18219	:douta	=	16'h	e634;
18220	:douta	=	16'h	de12;
18221	:douta	=	16'h	d5b1;
18222	:douta	=	16'h	cd71;
18223	:douta	=	16'h	bcf0;
18224	:douta	=	16'h	9beb;
18225	:douta	=	16'h	ac8d;
18226	:douta	=	16'h	7285;
18227	:douta	=	16'h	b4ce;
18228	:douta	=	16'h	bd30;
18229	:douta	=	16'h	acae;
18230	:douta	=	16'h	bd2f;
18231	:douta	=	16'h	c54f;
18232	:douta	=	16'h	c550;
18233	:douta	=	16'h	cd71;
18234	:douta	=	16'h	d5b1;
18235	:douta	=	16'h	e634;
18236	:douta	=	16'h	e634;
18237	:douta	=	16'h	ee75;
18238	:douta	=	16'h	e655;
18239	:douta	=	16'h	de13;
18240	:douta	=	16'h	ddf3;
18241	:douta	=	16'h	d5d2;
18242	:douta	=	16'h	cd71;
18243	:douta	=	16'h	cd50;
18244	:douta	=	16'h	c531;
18245	:douta	=	16'h	bd11;
18246	:douta	=	16'h	acb1;
18247	:douta	=	16'h	a471;
18248	:douta	=	16'h	9c51;
18249	:douta	=	16'h	8c31;
18250	:douta	=	16'h	8411;
18251	:douta	=	16'h	8411;
18252	:douta	=	16'h	73d1;
18253	:douta	=	16'h	73d1;
18254	:douta	=	16'h	6370;
18255	:douta	=	16'h	5b50;
18256	:douta	=	16'h	6350;
18257	:douta	=	16'h	5b30;
18258	:douta	=	16'h	5330;
18259	:douta	=	16'h	6372;
18260	:douta	=	16'h	29a9;
18261	:douta	=	16'h	18e5;
18262	:douta	=	16'h	10e6;
18263	:douta	=	16'h	2146;
18264	:douta	=	16'h	39ea;
18265	:douta	=	16'h	0862;
18266	:douta	=	16'h	10a4;
18267	:douta	=	16'h	10e4;
18268	:douta	=	16'h	10c4;
18269	:douta	=	16'h	10c4;
18270	:douta	=	16'h	10c4;
18271	:douta	=	16'h	10a3;
18272	:douta	=	16'h	10c5;
18273	:douta	=	16'h	1905;
18274	:douta	=	16'h	1084;
18275	:douta	=	16'h	0042;
18276	:douta	=	16'h	2188;
18277	:douta	=	16'h	08a5;
18278	:douta	=	16'h	18c5;
18279	:douta	=	16'h	840d;
18280	:douta	=	16'h	39a6;
18281	:douta	=	16'h	bd72;
18282	:douta	=	16'h	5ac9;
18283	:douta	=	16'h	39a7;
18284	:douta	=	16'h	3186;
18285	:douta	=	16'h	5269;
18286	:douta	=	16'h	b510;
18287	:douta	=	16'h	630c;
18288	:douta	=	16'h	2967;
18289	:douta	=	16'h	632d;
18290	:douta	=	16'h	29a9;
18291	:douta	=	16'h	2187;
18292	:douta	=	16'h	5acb;
18293	:douta	=	16'h	2146;
18294	:douta	=	16'h	6b4d;
18295	:douta	=	16'h	7c95;
18296	:douta	=	16'h	84d7;
18297	:douta	=	16'h	8d38;
18298	:douta	=	16'h	8d38;
18299	:douta	=	16'h	84f8;
18300	:douta	=	16'h	957a;
18301	:douta	=	16'h	9559;
18302	:douta	=	16'h	7476;
18303	:douta	=	16'h	7c97;
18304	:douta	=	16'h	84b8;
18305	:douta	=	16'h	9559;
18306	:douta	=	16'h	9dba;
18307	:douta	=	16'h	7456;
18308	:douta	=	16'h	5352;
18309	:douta	=	16'h	5bb2;
18310	:douta	=	16'h	84f7;
18311	:douta	=	16'h	a5ba;
18312	:douta	=	16'h	8d18;
18313	:douta	=	16'h	9579;
18314	:douta	=	16'h	a5ba;
18315	:douta	=	16'h	9579;
18316	:douta	=	16'h	9579;
18317	:douta	=	16'h	959a;
18318	:douta	=	16'h	9d9a;
18319	:douta	=	16'h	a5da;
18320	:douta	=	16'h	a5da;
18321	:douta	=	16'h	9579;
18322	:douta	=	16'h	8d59;
18323	:douta	=	16'h	9d9a;
18324	:douta	=	16'h	9d9a;
18325	:douta	=	16'h	9559;
18326	:douta	=	16'h	adfa;
18327	:douta	=	16'h	a5db;
18328	:douta	=	16'h	9559;
18329	:douta	=	16'h	a5db;
18330	:douta	=	16'h	9d9a;
18331	:douta	=	16'h	a5fb;
18332	:douta	=	16'h	8d59;
18333	:douta	=	16'h	7cd8;
18334	:douta	=	16'h	8539;
18335	:douta	=	16'h	959a;
18336	:douta	=	16'h	957a;
18337	:douta	=	16'h	8d39;
18338	:douta	=	16'h	9dbb;
18339	:douta	=	16'h	94f6;
18340	:douta	=	16'h	bccf;
18341	:douta	=	16'h	2126;
18342	:douta	=	16'h	18e5;
18343	:douta	=	16'h	0042;
18344	:douta	=	16'h	9ddc;
18345	:douta	=	16'h	957a;
18346	:douta	=	16'h	8d39;
18347	:douta	=	16'h	8d39;
18348	:douta	=	16'h	84b8;
18349	:douta	=	16'h	84d8;
18350	:douta	=	16'h	84d8;
18351	:douta	=	16'h	957a;
18352	:douta	=	16'h	7c76;
18353	:douta	=	16'h	84b7;
18354	:douta	=	16'h	9539;
18355	:douta	=	16'h	9d9a;
18356	:douta	=	16'h	9559;
18357	:douta	=	16'h	8518;
18358	:douta	=	16'h	8cf8;
18359	:douta	=	16'h	9d99;
18360	:douta	=	16'h	9d58;
18361	:douta	=	16'h	8cd6;
18362	:douta	=	16'h	94f6;
18363	:douta	=	16'h	8c75;
18364	:douta	=	16'h	8d18;
18365	:douta	=	16'h	9539;
18366	:douta	=	16'h	7455;
18367	:douta	=	16'h	7455;
18368	:douta	=	16'h	84b7;
18369	:douta	=	16'h	84b8;
18370	:douta	=	16'h	84f8;
18371	:douta	=	16'h	7cd8;
18372	:douta	=	16'h	8d7b;
18373	:douta	=	16'h	31a7;
18374	:douta	=	16'h	2126;
18375	:douta	=	16'h	10e5;
18376	:douta	=	16'h	2104;
18377	:douta	=	16'h	426d;
18378	:douta	=	16'h	5c16;
18379	:douta	=	16'h	6478;
18380	:douta	=	16'h	751a;
18381	:douta	=	16'h	7d3b;
18382	:douta	=	16'h	5c36;
18383	:douta	=	16'h	3b34;
18384	:douta	=	16'h	5417;
18385	:douta	=	16'h	7d5c;
18386	:douta	=	16'h	6cb9;
18387	:douta	=	16'h	53f6;
18388	:douta	=	16'h	5c16;
18389	:douta	=	16'h	5bf6;
18390	:douta	=	16'h	6c77;
18391	:douta	=	16'h	857b;
18392	:douta	=	16'h	8d9c;
18393	:douta	=	16'h	855b;
18394	:douta	=	16'h	6c77;
18395	:douta	=	16'h	7498;
18396	:douta	=	16'h	7cd9;
18397	:douta	=	16'h	74b8;
18398	:douta	=	16'h	7cd9;
18399	:douta	=	16'h	7cf9;
18400	:douta	=	16'h	853a;
18401	:douta	=	16'h	7cd9;
18402	:douta	=	16'h	853a;
18403	:douta	=	16'h	7cd9;
18404	:douta	=	16'h	7cd9;
18405	:douta	=	16'h	7cf9;
18406	:douta	=	16'h	7cd9;
18407	:douta	=	16'h	8d5a;
18408	:douta	=	16'h	959b;
18409	:douta	=	16'h	6c77;
18410	:douta	=	16'h	74b8;
18411	:douta	=	16'h	853a;
18412	:douta	=	16'h	8d5a;
18413	:douta	=	16'h	7478;
18414	:douta	=	16'h	7cf9;
18415	:douta	=	16'h	853a;
18416	:douta	=	16'h	8dbc;
18417	:douta	=	16'h	855b;
18418	:douta	=	16'h	6477;
18419	:douta	=	16'h	8d7b;
18420	:douta	=	16'h	8d5b;
18421	:douta	=	16'h	39ca;
18422	:douta	=	16'h	7c95;
18423	:douta	=	16'h	be3a;
18424	:douta	=	16'h	63f4;
18425	:douta	=	16'h	5330;
18426	:douta	=	16'h	7c33;
18427	:douta	=	16'h	9d16;
18428	:douta	=	16'h	94f6;
18429	:douta	=	16'h	0000;
18430	:douta	=	16'h	7c33;
18431	:douta	=	16'h	5310;
18432	:douta	=	16'h	2106;
18433	:douta	=	16'h	32f2;
18434	:douta	=	16'h	53f7;
18435	:douta	=	16'h	32b0;
18436	:douta	=	16'h	4bb5;
18437	:douta	=	16'h	32b1;
18438	:douta	=	16'h	3ad1;
18439	:douta	=	16'h	5394;
18440	:douta	=	16'h	6457;
18441	:douta	=	16'h	7cb8;
18442	:douta	=	16'h	7c98;
18443	:douta	=	16'h	7478;
18444	:douta	=	16'h	63f5;
18445	:douta	=	16'h	3a6d;
18446	:douta	=	16'h	63b3;
18447	:douta	=	16'h	5b92;
18448	:douta	=	16'h	9493;
18449	:douta	=	16'h	a536;
18450	:douta	=	16'h	94f6;
18451	:douta	=	16'h	7bd2;
18452	:douta	=	16'h	9493;
18453	:douta	=	16'h	8c93;
18454	:douta	=	16'h	73f1;
18455	:douta	=	16'h	bd96;
18456	:douta	=	16'h	b596;
18457	:douta	=	16'h	ad54;
18458	:douta	=	16'h	8329;
18459	:douta	=	16'h	93ab;
18460	:douta	=	16'h	93cb;
18461	:douta	=	16'h	b46b;
18462	:douta	=	16'h	bcab;
18463	:douta	=	16'h	c50d;
18464	:douta	=	16'h	cd2e;
18465	:douta	=	16'h	cd2e;
18466	:douta	=	16'h	d5b0;
18467	:douta	=	16'h	d5b0;
18468	:douta	=	16'h	ddf3;
18469	:douta	=	16'h	ddd2;
18470	:douta	=	16'h	de13;
18471	:douta	=	16'h	eeb6;
18472	:douta	=	16'h	eeb6;
18473	:douta	=	16'h	ddd1;
18474	:douta	=	16'h	ddf3;
18475	:douta	=	16'h	e655;
18476	:douta	=	16'h	d5d2;
18477	:douta	=	16'h	cd70;
18478	:douta	=	16'h	bd10;
18479	:douta	=	16'h	c510;
18480	:douta	=	16'h	a44c;
18481	:douta	=	16'h	8349;
18482	:douta	=	16'h	8b69;
18483	:douta	=	16'h	a44d;
18484	:douta	=	16'h	b4ee;
18485	:douta	=	16'h	bd0f;
18486	:douta	=	16'h	c550;
18487	:douta	=	16'h	c570;
18488	:douta	=	16'h	ddd1;
18489	:douta	=	16'h	d5b2;
18490	:douta	=	16'h	ddf3;
18491	:douta	=	16'h	de13;
18492	:douta	=	16'h	de13;
18493	:douta	=	16'h	e634;
18494	:douta	=	16'h	e634;
18495	:douta	=	16'h	de34;
18496	:douta	=	16'h	de14;
18497	:douta	=	16'h	ddf3;
18498	:douta	=	16'h	d591;
18499	:douta	=	16'h	cd50;
18500	:douta	=	16'h	c511;
18501	:douta	=	16'h	bcf1;
18502	:douta	=	16'h	b4d1;
18503	:douta	=	16'h	a491;
18504	:douta	=	16'h	9c72;
18505	:douta	=	16'h	9452;
18506	:douta	=	16'h	8c32;
18507	:douta	=	16'h	8412;
18508	:douta	=	16'h	7bf2;
18509	:douta	=	16'h	73f2;
18510	:douta	=	16'h	6bb1;
18511	:douta	=	16'h	6391;
18512	:douta	=	16'h	6bb1;
18513	:douta	=	16'h	6bd3;
18514	:douta	=	16'h	5b72;
18515	:douta	=	16'h	4acf;
18516	:douta	=	16'h	31a8;
18517	:douta	=	16'h	2168;
18518	:douta	=	16'h	39ca;
18519	:douta	=	16'h	10e5;
18520	:douta	=	16'h	3a2b;
18521	:douta	=	16'h	3a2c;
18522	:douta	=	16'h	1083;
18523	:douta	=	16'h	10a4;
18524	:douta	=	16'h	10e4;
18525	:douta	=	16'h	10c4;
18526	:douta	=	16'h	10c3;
18527	:douta	=	16'h	18c4;
18528	:douta	=	16'h	18e5;
18529	:douta	=	16'h	18e5;
18530	:douta	=	16'h	1905;
18531	:douta	=	16'h	10c4;
18532	:douta	=	16'h	08c5;
18533	:douta	=	16'h	0884;
18534	:douta	=	16'h	4a8b;
18535	:douta	=	16'h	4aaa;
18536	:douta	=	16'h	5228;
18537	:douta	=	16'h	73cd;
18538	:douta	=	16'h	840e;
18539	:douta	=	16'h	840f;
18540	:douta	=	16'h	b4f1;
18541	:douta	=	16'h	83ce;
18542	:douta	=	16'h	83ac;
18543	:douta	=	16'h	5aca;
18544	:douta	=	16'h	18e4;
18545	:douta	=	16'h	7bae;
18546	:douta	=	16'h	736d;
18547	:douta	=	16'h	2967;
18548	:douta	=	16'h	630c;
18549	:douta	=	16'h	4a29;
18550	:douta	=	16'h	5a6a;
18551	:douta	=	16'h	63d2;
18552	:douta	=	16'h	9559;
18553	:douta	=	16'h	8d18;
18554	:douta	=	16'h	9539;
18555	:douta	=	16'h	84d7;
18556	:douta	=	16'h	7c96;
18557	:douta	=	16'h	84f8;
18558	:douta	=	16'h	8d18;
18559	:douta	=	16'h	84d8;
18560	:douta	=	16'h	6415;
18561	:douta	=	16'h	7456;
18562	:douta	=	16'h	7476;
18563	:douta	=	16'h	ae1c;
18564	:douta	=	16'h	9d9a;
18565	:douta	=	16'h	6414;
18566	:douta	=	16'h	5372;
18567	:douta	=	16'h	7c75;
18568	:douta	=	16'h	8d18;
18569	:douta	=	16'h	a5da;
18570	:douta	=	16'h	be5c;
18571	:douta	=	16'h	adfb;
18572	:douta	=	16'h	a5fa;
18573	:douta	=	16'h	9559;
18574	:douta	=	16'h	957a;
18575	:douta	=	16'h	9dba;
18576	:douta	=	16'h	9d7a;
18577	:douta	=	16'h	9d9a;
18578	:douta	=	16'h	9d9a;
18579	:douta	=	16'h	9dba;
18580	:douta	=	16'h	a5da;
18581	:douta	=	16'h	9dba;
18582	:douta	=	16'h	9d99;
18583	:douta	=	16'h	b63b;
18584	:douta	=	16'h	ae1b;
18585	:douta	=	16'h	957a;
18586	:douta	=	16'h	9579;
18587	:douta	=	16'h	9559;
18588	:douta	=	16'h	9d9a;
18589	:douta	=	16'h	9579;
18590	:douta	=	16'h	8d18;
18591	:douta	=	16'h	8539;
18592	:douta	=	16'h	9579;
18593	:douta	=	16'h	953a;
18594	:douta	=	16'h	8d18;
18595	:douta	=	16'h	94f7;
18596	:douta	=	16'h	b4d0;
18597	:douta	=	16'h	39a7;
18598	:douta	=	16'h	1105;
18599	:douta	=	16'h	1083;
18600	:douta	=	16'h	8519;
18601	:douta	=	16'h	9559;
18602	:douta	=	16'h	84f8;
18603	:douta	=	16'h	957a;
18604	:douta	=	16'h	957a;
18605	:douta	=	16'h	84d8;
18606	:douta	=	16'h	84b8;
18607	:douta	=	16'h	84d7;
18608	:douta	=	16'h	9559;
18609	:douta	=	16'h	8d18;
18610	:douta	=	16'h	7c76;
18611	:douta	=	16'h	84d7;
18612	:douta	=	16'h	a5ba;
18613	:douta	=	16'h	957a;
18614	:douta	=	16'h	9539;
18615	:douta	=	16'h	9558;
18616	:douta	=	16'h	8495;
18617	:douta	=	16'h	8cd6;
18618	:douta	=	16'h	9517;
18619	:douta	=	16'h	9516;
18620	:douta	=	16'h	9518;
18621	:douta	=	16'h	8d18;
18622	:douta	=	16'h	9559;
18623	:douta	=	16'h	84d8;
18624	:douta	=	16'h	6c55;
18625	:douta	=	16'h	84d8;
18626	:douta	=	16'h	84f8;
18627	:douta	=	16'h	7cd8;
18628	:douta	=	16'h	8d9b;
18629	:douta	=	16'h	1905;
18630	:douta	=	16'h	1906;
18631	:douta	=	16'h	08c4;
18632	:douta	=	16'h	2125;
18633	:douta	=	16'h	4b10;
18634	:douta	=	16'h	6478;
18635	:douta	=	16'h	5c37;
18636	:douta	=	16'h	74b9;
18637	:douta	=	16'h	6cd9;
18638	:douta	=	16'h	6cb9;
18639	:douta	=	16'h	53f7;
18640	:douta	=	16'h	4353;
18641	:douta	=	16'h	4b74;
18642	:douta	=	16'h	74fa;
18643	:douta	=	16'h	855b;
18644	:douta	=	16'h	32f2;
18645	:douta	=	16'h	5c37;
18646	:douta	=	16'h	6cb9;
18647	:douta	=	16'h	5bd5;
18648	:douta	=	16'h	6c57;
18649	:douta	=	16'h	8ddd;
18650	:douta	=	16'h	74d9;
18651	:douta	=	16'h	7cf9;
18652	:douta	=	16'h	74d9;
18653	:douta	=	16'h	7d1a;
18654	:douta	=	16'h	8d5b;
18655	:douta	=	16'h	6c77;
18656	:douta	=	16'h	7cf9;
18657	:douta	=	16'h	6c77;
18658	:douta	=	16'h	7497;
18659	:douta	=	16'h	8d3a;
18660	:douta	=	16'h	7cf9;
18661	:douta	=	16'h	7cd9;
18662	:douta	=	16'h	84f9;
18663	:douta	=	16'h	7498;
18664	:douta	=	16'h	8519;
18665	:douta	=	16'h	959b;
18666	:douta	=	16'h	7cd9;
18667	:douta	=	16'h	7498;
18668	:douta	=	16'h	7cb8;
18669	:douta	=	16'h	8d9b;
18670	:douta	=	16'h	7497;
18671	:douta	=	16'h	6c36;
18672	:douta	=	16'h	74b8;
18673	:douta	=	16'h	7cf9;
18674	:douta	=	16'h	7cd9;
18675	:douta	=	16'h	6c77;
18676	:douta	=	16'h	63f3;
18677	:douta	=	16'h	42ad;
18678	:douta	=	16'h	6bf3;
18679	:douta	=	16'h	a5b9;
18680	:douta	=	16'h	6c34;
18681	:douta	=	16'h	a598;
18682	:douta	=	16'h	7c33;
18683	:douta	=	16'h	63b1;
18684	:douta	=	16'h	8432;
18685	:douta	=	16'h	2127;
18686	:douta	=	16'h	9d58;
18687	:douta	=	16'h	8c95;
18688	:douta	=	16'h	1884;
18689	:douta	=	16'h	2a4f;
18690	:douta	=	16'h	3ad2;
18691	:douta	=	16'h	21ec;
18692	:douta	=	16'h	53d5;
18693	:douta	=	16'h	53d6;
18694	:douta	=	16'h	3ad2;
18695	:douta	=	16'h	32f2;
18696	:douta	=	16'h	6457;
18697	:douta	=	16'h	4b31;
18698	:douta	=	16'h	5b73;
18699	:douta	=	16'h	6416;
18700	:douta	=	16'h	5b93;
18701	:douta	=	16'h	4acf;
18702	:douta	=	16'h	7c76;
18703	:douta	=	16'h	8cd7;
18704	:douta	=	16'h	6bb1;
18705	:douta	=	16'h	8453;
18706	:douta	=	16'h	6bb1;
18707	:douta	=	16'h	8433;
18708	:douta	=	16'h	9cd4;
18709	:douta	=	16'h	bdd7;
18710	:douta	=	16'h	a535;
18711	:douta	=	16'h	9c93;
18712	:douta	=	16'h	7b6c;
18713	:douta	=	16'h	7b0a;
18714	:douta	=	16'h	8bab;
18715	:douta	=	16'h	9c0b;
18716	:douta	=	16'h	a40b;
18717	:douta	=	16'h	c50e;
18718	:douta	=	16'h	cd6e;
18719	:douta	=	16'h	c52e;
18720	:douta	=	16'h	cd6e;
18721	:douta	=	16'h	d590;
18722	:douta	=	16'h	de13;
18723	:douta	=	16'h	e634;
18724	:douta	=	16'h	e695;
18725	:douta	=	16'h	e655;
18726	:douta	=	16'h	ee75;
18727	:douta	=	16'h	e654;
18728	:douta	=	16'h	ee75;
18729	:douta	=	16'h	ee96;
18730	:douta	=	16'h	e654;
18731	:douta	=	16'h	d5d3;
18732	:douta	=	16'h	cd71;
18733	:douta	=	16'h	b4ad;
18734	:douta	=	16'h	ac6d;
18735	:douta	=	16'h	b4ae;
18736	:douta	=	16'h	7b09;
18737	:douta	=	16'h	9c0c;
18738	:douta	=	16'h	9c0c;
18739	:douta	=	16'h	a42d;
18740	:douta	=	16'h	ac8e;
18741	:douta	=	16'h	bd0f;
18742	:douta	=	16'h	cd70;
18743	:douta	=	16'h	cd91;
18744	:douta	=	16'h	d5f2;
18745	:douta	=	16'h	de13;
18746	:douta	=	16'h	de34;
18747	:douta	=	16'h	e654;
18748	:douta	=	16'h	e654;
18749	:douta	=	16'h	e654;
18750	:douta	=	16'h	e634;
18751	:douta	=	16'h	de13;
18752	:douta	=	16'h	ddf3;
18753	:douta	=	16'h	d5b3;
18754	:douta	=	16'h	cd71;
18755	:douta	=	16'h	c551;
18756	:douta	=	16'h	bcf1;
18757	:douta	=	16'h	bd11;
18758	:douta	=	16'h	acb0;
18759	:douta	=	16'h	9451;
18760	:douta	=	16'h	8c31;
18761	:douta	=	16'h	9c72;
18762	:douta	=	16'h	9472;
18763	:douta	=	16'h	8c73;
18764	:douta	=	16'h	8433;
18765	:douta	=	16'h	8433;
18766	:douta	=	16'h	8c74;
18767	:douta	=	16'h	8c74;
18768	:douta	=	16'h	7c13;
18769	:douta	=	16'h	5352;
18770	:douta	=	16'h	1948;
18771	:douta	=	16'h	9bca;
18772	:douta	=	16'h	320b;
18773	:douta	=	16'h	39ea;
18774	:douta	=	16'h	420a;
18775	:douta	=	16'h	2167;
18776	:douta	=	16'h	10c5;
18777	:douta	=	16'h	0042;
18778	:douta	=	16'h	428d;
18779	:douta	=	16'h	1083;
18780	:douta	=	16'h	18e4;
18781	:douta	=	16'h	10c5;
18782	:douta	=	16'h	18e5;
18783	:douta	=	16'h	18e4;
18784	:douta	=	16'h	10c4;
18785	:douta	=	16'h	10e4;
18786	:douta	=	16'h	10e4;
18787	:douta	=	16'h	18e5;
18788	:douta	=	16'h	2126;
18789	:douta	=	16'h	21a8;
18790	:douta	=	16'h	855a;
18791	:douta	=	16'h	52cd;
18792	:douta	=	16'h	73f1;
18793	:douta	=	16'h	4a28;
18794	:douta	=	16'h	7bce;
18795	:douta	=	16'h	2946;
18796	:douta	=	16'h	6b2b;
18797	:douta	=	16'h	3145;
18798	:douta	=	16'h	31c8;
18799	:douta	=	16'h	2945;
18800	:douta	=	16'h	62ca;
18801	:douta	=	16'h	7b6d;
18802	:douta	=	16'h	bd72;
18803	:douta	=	16'h	944f;
18804	:douta	=	16'h	4167;
18805	:douta	=	16'h	630c;
18806	:douta	=	16'h	4a08;
18807	:douta	=	16'h	62ec;
18808	:douta	=	16'h	8d59;
18809	:douta	=	16'h	9559;
18810	:douta	=	16'h	9539;
18811	:douta	=	16'h	7c96;
18812	:douta	=	16'h	7c96;
18813	:douta	=	16'h	84d7;
18814	:douta	=	16'h	8d39;
18815	:douta	=	16'h	8d39;
18816	:douta	=	16'h	84f8;
18817	:douta	=	16'h	7cb7;
18818	:douta	=	16'h	84b7;
18819	:douta	=	16'h	84d7;
18820	:douta	=	16'h	84d7;
18821	:douta	=	16'h	84d7;
18822	:douta	=	16'h	84f8;
18823	:douta	=	16'h	9579;
18824	:douta	=	16'h	8518;
18825	:douta	=	16'h	7c96;
18826	:douta	=	16'h	7cb6;
18827	:douta	=	16'h	84b6;
18828	:douta	=	16'h	7cb6;
18829	:douta	=	16'h	9d9a;
18830	:douta	=	16'h	ae3c;
18831	:douta	=	16'h	9d99;
18832	:douta	=	16'h	8d18;
18833	:douta	=	16'h	a5da;
18834	:douta	=	16'h	8d38;
18835	:douta	=	16'h	a5ba;
18836	:douta	=	16'h	9d9a;
18837	:douta	=	16'h	9579;
18838	:douta	=	16'h	9dba;
18839	:douta	=	16'h	a5da;
18840	:douta	=	16'h	a5ba;
18841	:douta	=	16'h	ae1b;
18842	:douta	=	16'h	ae1b;
18843	:douta	=	16'h	9d9a;
18844	:douta	=	16'h	9dba;
18845	:douta	=	16'h	9d9a;
18846	:douta	=	16'h	adfa;
18847	:douta	=	16'h	a5da;
18848	:douta	=	16'h	a5da;
18849	:douta	=	16'h	8d39;
18850	:douta	=	16'h	8d38;
18851	:douta	=	16'h	8d39;
18852	:douta	=	16'h	9d16;
18853	:douta	=	16'h	ac6d;
18854	:douta	=	16'h	0063;
18855	:douta	=	16'h	10c4;
18856	:douta	=	16'h	5392;
18857	:douta	=	16'h	a5fc;
18858	:douta	=	16'h	9d7a;
18859	:douta	=	16'h	84d8;
18860	:douta	=	16'h	7cb8;
18861	:douta	=	16'h	8d5a;
18862	:douta	=	16'h	8d5a;
18863	:douta	=	16'h	8d39;
18864	:douta	=	16'h	8d38;
18865	:douta	=	16'h	9d59;
18866	:douta	=	16'h	7c76;
18867	:douta	=	16'h	7c76;
18868	:douta	=	16'h	84b7;
18869	:douta	=	16'h	7c55;
18870	:douta	=	16'h	9d58;
18871	:douta	=	16'h	9d58;
18872	:douta	=	16'h	8cf7;
18873	:douta	=	16'h	a578;
18874	:douta	=	16'h	9d58;
18875	:douta	=	16'h	9d37;
18876	:douta	=	16'h	9558;
18877	:douta	=	16'h	8d18;
18878	:douta	=	16'h	955a;
18879	:douta	=	16'h	8d7a;
18880	:douta	=	16'h	8d5a;
18881	:douta	=	16'h	959b;
18882	:douta	=	16'h	8d39;
18883	:douta	=	16'h	851a;
18884	:douta	=	16'h	8519;
18885	:douta	=	16'h	3167;
18886	:douta	=	16'h	0884;
18887	:douta	=	16'h	10a4;
18888	:douta	=	16'h	39c9;
18889	:douta	=	16'h	6457;
18890	:douta	=	16'h	7d3a;
18891	:douta	=	16'h	74b9;
18892	:douta	=	16'h	6c99;
18893	:douta	=	16'h	6cb9;
18894	:douta	=	16'h	751a;
18895	:douta	=	16'h	855b;
18896	:douta	=	16'h	74fa;
18897	:douta	=	16'h	7d1b;
18898	:douta	=	16'h	7d3a;
18899	:douta	=	16'h	53d5;
18900	:douta	=	16'h	4354;
18901	:douta	=	16'h	855b;
18902	:douta	=	16'h	7d3a;
18903	:douta	=	16'h	6437;
18904	:douta	=	16'h	5bf6;
18905	:douta	=	16'h	53d4;
18906	:douta	=	16'h	6c98;
18907	:douta	=	16'h	6c98;
18908	:douta	=	16'h	855b;
18909	:douta	=	16'h	853a;
18910	:douta	=	16'h	7477;
18911	:douta	=	16'h	7478;
18912	:douta	=	16'h	7cf9;
18913	:douta	=	16'h	8d7b;
18914	:douta	=	16'h	853a;
18915	:douta	=	16'h	8d5b;
18916	:douta	=	16'h	853a;
18917	:douta	=	16'h	84f9;
18918	:douta	=	16'h	7cf9;
18919	:douta	=	16'h	851a;
18920	:douta	=	16'h	8519;
18921	:douta	=	16'h	855a;
18922	:douta	=	16'h	7cd9;
18923	:douta	=	16'h	851a;
18924	:douta	=	16'h	95dc;
18925	:douta	=	16'h	851a;
18926	:douta	=	16'h	6436;
18927	:douta	=	16'h	7457;
18928	:douta	=	16'h	95bc;
18929	:douta	=	16'h	95bc;
18930	:douta	=	16'h	7cf9;
18931	:douta	=	16'h	6bf3;
18932	:douta	=	16'h	39a8;
18933	:douta	=	16'h	84d6;
18934	:douta	=	16'h	9538;
18935	:douta	=	16'h	8cf7;
18936	:douta	=	16'h	6c14;
18937	:douta	=	16'h	4b11;
18938	:douta	=	16'h	63d2;
18939	:douta	=	16'h	7413;
18940	:douta	=	16'h	28e3;
18941	:douta	=	16'h	7454;
18942	:douta	=	16'h	9515;
18943	:douta	=	16'h	8c95;
18944	:douta	=	16'h	10c2;
18945	:douta	=	16'h	2a0c;
18946	:douta	=	16'h	4354;
18947	:douta	=	16'h	2a6f;
18948	:douta	=	16'h	3b12;
18949	:douta	=	16'h	53f6;
18950	:douta	=	16'h	116b;
18951	:douta	=	16'h	226f;
18952	:douta	=	16'h	6436;
18953	:douta	=	16'h	5bd4;
18954	:douta	=	16'h	7456;
18955	:douta	=	16'h	7d1a;
18956	:douta	=	16'h	74b9;
18957	:douta	=	16'h	322c;
18958	:douta	=	16'h	63f4;
18959	:douta	=	16'h	5331;
18960	:douta	=	16'h	7413;
18961	:douta	=	16'h	8c95;
18962	:douta	=	16'h	9d16;
18963	:douta	=	16'h	7c13;
18964	:douta	=	16'h	9cd4;
18965	:douta	=	16'h	636f;
18966	:douta	=	16'h	8411;
18967	:douta	=	16'h	b556;
18968	:douta	=	16'h	7b2b;
18969	:douta	=	16'h	8bcb;
18970	:douta	=	16'h	93cb;
18971	:douta	=	16'h	ac4b;
18972	:douta	=	16'h	ac4b;
18973	:douta	=	16'h	cd4e;
18974	:douta	=	16'h	cd6f;
18975	:douta	=	16'h	cd6f;
18976	:douta	=	16'h	d5b0;
18977	:douta	=	16'h	ddd1;
18978	:douta	=	16'h	de34;
18979	:douta	=	16'h	e655;
18980	:douta	=	16'h	e674;
18981	:douta	=	16'h	e634;
18982	:douta	=	16'h	eeb6;
18983	:douta	=	16'h	e634;
18984	:douta	=	16'h	e675;
18985	:douta	=	16'h	e654;
18986	:douta	=	16'h	e634;
18987	:douta	=	16'h	cd92;
18988	:douta	=	16'h	d5d2;
18989	:douta	=	16'h	c530;
18990	:douta	=	16'h	a42c;
18991	:douta	=	16'h	a42c;
18992	:douta	=	16'h	8b8a;
18993	:douta	=	16'h	9beb;
18994	:douta	=	16'h	a42c;
18995	:douta	=	16'h	a44d;
18996	:douta	=	16'h	ac8d;
18997	:douta	=	16'h	bcee;
18998	:douta	=	16'h	d591;
18999	:douta	=	16'h	d5b1;
19000	:douta	=	16'h	ddf2;
19001	:douta	=	16'h	de13;
19002	:douta	=	16'h	e654;
19003	:douta	=	16'h	e654;
19004	:douta	=	16'h	e654;
19005	:douta	=	16'h	e654;
19006	:douta	=	16'h	e654;
19007	:douta	=	16'h	ddf3;
19008	:douta	=	16'h	ddf3;
19009	:douta	=	16'h	d5b3;
19010	:douta	=	16'h	c531;
19011	:douta	=	16'h	c531;
19012	:douta	=	16'h	bd11;
19013	:douta	=	16'h	bcf1;
19014	:douta	=	16'h	acb0;
19015	:douta	=	16'h	8c31;
19016	:douta	=	16'h	9431;
19017	:douta	=	16'h	9452;
19018	:douta	=	16'h	8c72;
19019	:douta	=	16'h	8c53;
19020	:douta	=	16'h	8c53;
19021	:douta	=	16'h	7c12;
19022	:douta	=	16'h	8c74;
19023	:douta	=	16'h	7c33;
19024	:douta	=	16'h	a556;
19025	:douta	=	16'h	31a8;
19026	:douta	=	16'h	69e3;
19027	:douta	=	16'h	b50f;
19028	:douta	=	16'h	3a0b;
19029	:douta	=	16'h	424a;
19030	:douta	=	16'h	4209;
19031	:douta	=	16'h	2987;
19032	:douta	=	16'h	1906;
19033	:douta	=	16'h	18e4;
19034	:douta	=	16'h	2147;
19035	:douta	=	16'h	2147;
19036	:douta	=	16'h	0863;
19037	:douta	=	16'h	10c4;
19038	:douta	=	16'h	10a4;
19039	:douta	=	16'h	10c4;
19040	:douta	=	16'h	10a4;
19041	:douta	=	16'h	10a4;
19042	:douta	=	16'h	18e5;
19043	:douta	=	16'h	18c4;
19044	:douta	=	16'h	1906;
19045	:douta	=	16'h	0001;
19046	:douta	=	16'h	08e5;
19047	:douta	=	16'h	84f7;
19048	:douta	=	16'h	4aac;
19049	:douta	=	16'h	31a8;
19050	:douta	=	16'h	6bce;
19051	:douta	=	16'h	08a3;
19052	:douta	=	16'h	8c0f;
19053	:douta	=	16'h	83cd;
19054	:douta	=	16'h	5aca;
19055	:douta	=	16'h	736c;
19056	:douta	=	16'h	5a8a;
19057	:douta	=	16'h	2146;
19058	:douta	=	16'h	5269;
19059	:douta	=	16'h	39a6;
19060	:douta	=	16'h	bd92;
19061	:douta	=	16'h	634b;
19062	:douta	=	16'h	9c70;
19063	:douta	=	16'h	6aca;
19064	:douta	=	16'h	a61c;
19065	:douta	=	16'h	84f8;
19066	:douta	=	16'h	9d7a;
19067	:douta	=	16'h	8d39;
19068	:douta	=	16'h	8d59;
19069	:douta	=	16'h	84d7;
19070	:douta	=	16'h	8d39;
19071	:douta	=	16'h	8d39;
19072	:douta	=	16'h	8d18;
19073	:douta	=	16'h	8d18;
19074	:douta	=	16'h	7c96;
19075	:douta	=	16'h	84f8;
19076	:douta	=	16'h	84d7;
19077	:douta	=	16'h	8d18;
19078	:douta	=	16'h	84f8;
19079	:douta	=	16'h	84d7;
19080	:douta	=	16'h	9579;
19081	:douta	=	16'h	8d18;
19082	:douta	=	16'h	8d39;
19083	:douta	=	16'h	9559;
19084	:douta	=	16'h	8518;
19085	:douta	=	16'h	6c35;
19086	:douta	=	16'h	6c15;
19087	:douta	=	16'h	addb;
19088	:douta	=	16'h	adfb;
19089	:douta	=	16'h	8d39;
19090	:douta	=	16'h	adda;
19091	:douta	=	16'h	b63b;
19092	:douta	=	16'h	9d9a;
19093	:douta	=	16'h	9d7a;
19094	:douta	=	16'h	8d18;
19095	:douta	=	16'h	9579;
19096	:douta	=	16'h	9599;
19097	:douta	=	16'h	8d59;
19098	:douta	=	16'h	9599;
19099	:douta	=	16'h	adfa;
19100	:douta	=	16'h	a5ba;
19101	:douta	=	16'h	adda;
19102	:douta	=	16'h	a5da;
19103	:douta	=	16'h	9d9a;
19104	:douta	=	16'h	a5ba;
19105	:douta	=	16'h	8d39;
19106	:douta	=	16'h	8518;
19107	:douta	=	16'h	9dba;
19108	:douta	=	16'h	9538;
19109	:douta	=	16'h	cd2f;
19110	:douta	=	16'h	1083;
19111	:douta	=	16'h	0063;
19112	:douta	=	16'h	29e9;
19113	:douta	=	16'h	8d5a;
19114	:douta	=	16'h	9538;
19115	:douta	=	16'h	8d39;
19116	:douta	=	16'h	6c35;
19117	:douta	=	16'h	7497;
19118	:douta	=	16'h	8539;
19119	:douta	=	16'h	8d39;
19120	:douta	=	16'h	84f8;
19121	:douta	=	16'h	9539;
19122	:douta	=	16'h	9d79;
19123	:douta	=	16'h	8496;
19124	:douta	=	16'h	84b6;
19125	:douta	=	16'h	7c54;
19126	:douta	=	16'h	7c55;
19127	:douta	=	16'h	8cb6;
19128	:douta	=	16'h	8496;
19129	:douta	=	16'h	9517;
19130	:douta	=	16'h	8cd6;
19131	:douta	=	16'h	8cb6;
19132	:douta	=	16'h	9538;
19133	:douta	=	16'h	8d39;
19134	:douta	=	16'h	9dbb;
19135	:douta	=	16'h	9dbb;
19136	:douta	=	16'h	8d39;
19137	:douta	=	16'h	8d5a;
19138	:douta	=	16'h	959b;
19139	:douta	=	16'h	8d9b;
19140	:douta	=	16'h	63d3;
19141	:douta	=	16'h	2987;
19142	:douta	=	16'h	1083;
19143	:douta	=	16'h	2146;
19144	:douta	=	16'h	426c;
19145	:douta	=	16'h	7d5c;
19146	:douta	=	16'h	7d1a;
19147	:douta	=	16'h	7d3b;
19148	:douta	=	16'h	7d1a;
19149	:douta	=	16'h	6c98;
19150	:douta	=	16'h	6c98;
19151	:douta	=	16'h	857b;
19152	:douta	=	16'h	857b;
19153	:douta	=	16'h	7d1a;
19154	:douta	=	16'h	857b;
19155	:douta	=	16'h	9ddd;
19156	:douta	=	16'h	5c17;
19157	:douta	=	16'h	5c16;
19158	:douta	=	16'h	5c16;
19159	:douta	=	16'h	7d3b;
19160	:douta	=	16'h	74b9;
19161	:douta	=	16'h	5c16;
19162	:douta	=	16'h	6437;
19163	:douta	=	16'h	6437;
19164	:douta	=	16'h	74b8;
19165	:douta	=	16'h	7498;
19166	:douta	=	16'h	7d1a;
19167	:douta	=	16'h	6c36;
19168	:douta	=	16'h	7477;
19169	:douta	=	16'h	8519;
19170	:douta	=	16'h	7477;
19171	:douta	=	16'h	855a;
19172	:douta	=	16'h	959b;
19173	:douta	=	16'h	8d9b;
19174	:douta	=	16'h	853a;
19175	:douta	=	16'h	7cfa;
19176	:douta	=	16'h	84f9;
19177	:douta	=	16'h	8d7b;
19178	:douta	=	16'h	8d9b;
19179	:douta	=	16'h	851a;
19180	:douta	=	16'h	74b8;
19181	:douta	=	16'h	8d7b;
19182	:douta	=	16'h	95dc;
19183	:douta	=	16'h	7cd8;
19184	:douta	=	16'h	6416;
19185	:douta	=	16'h	74b8;
19186	:douta	=	16'h	853a;
19187	:douta	=	16'h	41ea;
19188	:douta	=	16'h	52cd;
19189	:douta	=	16'h	7434;
19190	:douta	=	16'h	6c13;
19191	:douta	=	16'h	6392;
19192	:douta	=	16'h	9d58;
19193	:douta	=	16'h	8d17;
19194	:douta	=	16'h	9d79;
19195	:douta	=	16'h	9559;
19196	:douta	=	16'h	0800;
19197	:douta	=	16'h	63f4;
19198	:douta	=	16'h	8474;
19199	:douta	=	16'h	8474;
19200	:douta	=	16'h	1082;
19201	:douta	=	16'h	324d;
19202	:douta	=	16'h	53f7;
19203	:douta	=	16'h	21ed;
19204	:douta	=	16'h	2a4e;
19205	:douta	=	16'h	19cc;
19206	:douta	=	16'h	4354;
19207	:douta	=	16'h	32f2;
19208	:douta	=	16'h	74d9;
19209	:douta	=	16'h	5352;
19210	:douta	=	16'h	7477;
19211	:douta	=	16'h	74b8;
19212	:douta	=	16'h	6c36;
19213	:douta	=	16'h	6392;
19214	:douta	=	16'h	7435;
19215	:douta	=	16'h	8497;
19216	:douta	=	16'h	8cb6;
19217	:douta	=	16'h	8c95;
19218	:douta	=	16'h	9d16;
19219	:douta	=	16'h	5b30;
19220	:douta	=	16'h	6b90;
19221	:douta	=	16'h	8c52;
19222	:douta	=	16'h	8c72;
19223	:douta	=	16'h	8bcb;
19224	:douta	=	16'h	93ac;
19225	:douta	=	16'h	938b;
19226	:douta	=	16'h	a42b;
19227	:douta	=	16'h	bcad;
19228	:douta	=	16'h	bccd;
19229	:douta	=	16'h	cd4f;
19230	:douta	=	16'h	d5b1;
19231	:douta	=	16'h	cd6f;
19232	:douta	=	16'h	d5b0;
19233	:douta	=	16'h	e633;
19234	:douta	=	16'h	ee95;
19235	:douta	=	16'h	ee96;
19236	:douta	=	16'h	ee96;
19237	:douta	=	16'h	e634;
19238	:douta	=	16'h	ddf3;
19239	:douta	=	16'h	eeb6;
19240	:douta	=	16'h	e654;
19241	:douta	=	16'h	ddf2;
19242	:douta	=	16'h	d5d1;
19243	:douta	=	16'h	c50e;
19244	:douta	=	16'h	bd0f;
19245	:douta	=	16'h	b4ce;
19246	:douta	=	16'h	8349;
19247	:douta	=	16'h	8b8a;
19248	:douta	=	16'h	93eb;
19249	:douta	=	16'h	a42d;
19250	:douta	=	16'h	ac4c;
19251	:douta	=	16'h	c54f;
19252	:douta	=	16'h	c54f;
19253	:douta	=	16'h	d5b0;
19254	:douta	=	16'h	d5d2;
19255	:douta	=	16'h	de13;
19256	:douta	=	16'h	e675;
19257	:douta	=	16'h	ee75;
19258	:douta	=	16'h	e654;
19259	:douta	=	16'h	de14;
19260	:douta	=	16'h	e634;
19261	:douta	=	16'h	de33;
19262	:douta	=	16'h	de13;
19263	:douta	=	16'h	e613;
19264	:douta	=	16'h	cd91;
19265	:douta	=	16'h	cd72;
19266	:douta	=	16'h	bd12;
19267	:douta	=	16'h	bcf1;
19268	:douta	=	16'h	b4d1;
19269	:douta	=	16'h	b4d1;
19270	:douta	=	16'h	acb1;
19271	:douta	=	16'h	8c12;
19272	:douta	=	16'h	9452;
19273	:douta	=	16'h	8412;
19274	:douta	=	16'h	8c53;
19275	:douta	=	16'h	8c33;
19276	:douta	=	16'h	6b70;
19277	:douta	=	16'h	73f2;
19278	:douta	=	16'h	8c73;
19279	:douta	=	16'h	5b2f;
19280	:douta	=	16'h	2947;
19281	:douta	=	16'h	8b28;
19282	:douta	=	16'h	d590;
19283	:douta	=	16'h	9c2e;
19284	:douta	=	16'h	422b;
19285	:douta	=	16'h	5aac;
19286	:douta	=	16'h	422a;
19287	:douta	=	16'h	31ea;
19288	:douta	=	16'h	2147;
19289	:douta	=	16'h	10e5;
19290	:douta	=	16'h	1927;
19291	:douta	=	16'h	1906;
19292	:douta	=	16'h	4a8c;
19293	:douta	=	16'h	10a4;
19294	:douta	=	16'h	1084;
19295	:douta	=	16'h	10e4;
19296	:douta	=	16'h	10c4;
19297	:douta	=	16'h	10a4;
19298	:douta	=	16'h	10e4;
19299	:douta	=	16'h	10e4;
19300	:douta	=	16'h	10c5;
19301	:douta	=	16'h	1906;
19302	:douta	=	16'h	2187;
19303	:douta	=	16'h	0000;
19304	:douta	=	16'h	5371;
19305	:douta	=	16'h	6bb0;
19306	:douta	=	16'h	3a4c;
19307	:douta	=	16'h	940d;
19308	:douta	=	16'h	630c;
19309	:douta	=	16'h	accf;
19310	:douta	=	16'h	0883;
19311	:douta	=	16'h	0861;
19312	:douta	=	16'h	10c3;
19313	:douta	=	16'h	9cd1;
19314	:douta	=	16'h	1905;
19315	:douta	=	16'h	8c0d;
19316	:douta	=	16'h	8c4e;
19317	:douta	=	16'h	83ee;
19318	:douta	=	16'h	39e8;
19319	:douta	=	16'h	8bef;
19320	:douta	=	16'h	6c13;
19321	:douta	=	16'h	8cf8;
19322	:douta	=	16'h	8518;
19323	:douta	=	16'h	8d39;
19324	:douta	=	16'h	8d39;
19325	:douta	=	16'h	9d9a;
19326	:douta	=	16'h	8d38;
19327	:douta	=	16'h	8d38;
19328	:douta	=	16'h	9579;
19329	:douta	=	16'h	8517;
19330	:douta	=	16'h	8d18;
19331	:douta	=	16'h	7c96;
19332	:douta	=	16'h	7cb6;
19333	:douta	=	16'h	9579;
19334	:douta	=	16'h	9558;
19335	:douta	=	16'h	9538;
19336	:douta	=	16'h	84d7;
19337	:douta	=	16'h	8d38;
19338	:douta	=	16'h	8d39;
19339	:douta	=	16'h	8d58;
19340	:douta	=	16'h	7476;
19341	:douta	=	16'h	84f8;
19342	:douta	=	16'h	a5db;
19343	:douta	=	16'h	9579;
19344	:douta	=	16'h	8518;
19345	:douta	=	16'h	8d59;
19346	:douta	=	16'h	adda;
19347	:douta	=	16'h	a5ba;
19348	:douta	=	16'h	8d59;
19349	:douta	=	16'h	8d39;
19350	:douta	=	16'h	959a;
19351	:douta	=	16'h	7cb7;
19352	:douta	=	16'h	8d38;
19353	:douta	=	16'h	a5da;
19354	:douta	=	16'h	9d99;
19355	:douta	=	16'h	959a;
19356	:douta	=	16'h	9579;
19357	:douta	=	16'h	9d9a;
19358	:douta	=	16'h	9d9a;
19359	:douta	=	16'h	a5ba;
19360	:douta	=	16'h	9d99;
19361	:douta	=	16'h	9d7a;
19362	:douta	=	16'h	9db9;
19363	:douta	=	16'h	9579;
19364	:douta	=	16'h	957a;
19365	:douta	=	16'h	c4ee;
19366	:douta	=	16'h	c530;
19367	:douta	=	16'h	2926;
19368	:douta	=	16'h	1082;
19369	:douta	=	16'h	29ca;
19370	:douta	=	16'h	955a;
19371	:douta	=	16'h	9559;
19372	:douta	=	16'h	8d18;
19373	:douta	=	16'h	9dba;
19374	:douta	=	16'h	8d39;
19375	:douta	=	16'h	6c35;
19376	:douta	=	16'h	84b7;
19377	:douta	=	16'h	7c96;
19378	:douta	=	16'h	8cf7;
19379	:douta	=	16'h	84d7;
19380	:douta	=	16'h	7c75;
19381	:douta	=	16'h	84b6;
19382	:douta	=	16'h	9538;
19383	:douta	=	16'h	7c13;
19384	:douta	=	16'h	73f2;
19385	:douta	=	16'h	7c33;
19386	:douta	=	16'h	7c54;
19387	:douta	=	16'h	8cb6;
19388	:douta	=	16'h	84f8;
19389	:douta	=	16'h	7cb7;
19390	:douta	=	16'h	7477;
19391	:douta	=	16'h	7497;
19392	:douta	=	16'h	84f9;
19393	:douta	=	16'h	959a;
19394	:douta	=	16'h	851a;
19395	:douta	=	16'h	7476;
19396	:douta	=	16'h	2905;
19397	:douta	=	16'h	0884;
19398	:douta	=	16'h	2167;
19399	:douta	=	16'h	31c8;
19400	:douta	=	16'h	5bf4;
19401	:douta	=	16'h	74d9;
19402	:douta	=	16'h	74b8;
19403	:douta	=	16'h	7d3a;
19404	:douta	=	16'h	74f9;
19405	:douta	=	16'h	6436;
19406	:douta	=	16'h	6c78;
19407	:douta	=	16'h	6457;
19408	:douta	=	16'h	7d1a;
19409	:douta	=	16'h	74d9;
19410	:douta	=	16'h	8d7b;
19411	:douta	=	16'h	7cd9;
19412	:douta	=	16'h	9dfd;
19413	:douta	=	16'h	9e1d;
19414	:douta	=	16'h	9dfd;
19415	:douta	=	16'h	7cd9;
19416	:douta	=	16'h	6417;
19417	:douta	=	16'h	7498;
19418	:douta	=	16'h	6c98;
19419	:douta	=	16'h	74fa;
19420	:douta	=	16'h	5c37;
19421	:douta	=	16'h	53f6;
19422	:douta	=	16'h	7498;
19423	:douta	=	16'h	853a;
19424	:douta	=	16'h	7498;
19425	:douta	=	16'h	8d5a;
19426	:douta	=	16'h	7cd9;
19427	:douta	=	16'h	6c36;
19428	:douta	=	16'h	74b8;
19429	:douta	=	16'h	6c57;
19430	:douta	=	16'h	7cf9;
19431	:douta	=	16'h	8d7a;
19432	:douta	=	16'h	8539;
19433	:douta	=	16'h	851a;
19434	:douta	=	16'h	84d9;
19435	:douta	=	16'h	6c77;
19436	:douta	=	16'h	8d5b;
19437	:douta	=	16'h	959c;
19438	:douta	=	16'h	84f9;
19439	:douta	=	16'h	7cb8;
19440	:douta	=	16'h	855a;
19441	:douta	=	16'h	8d9b;
19442	:douta	=	16'h	6416;
19443	:douta	=	16'h	6391;
19444	:douta	=	16'h	8d3a;
19445	:douta	=	16'h	7454;
19446	:douta	=	16'h	7c95;
19447	:douta	=	16'h	9d58;
19448	:douta	=	16'h	7454;
19449	:douta	=	16'h	8475;
19450	:douta	=	16'h	7497;
19451	:douta	=	16'h	73f3;
19452	:douta	=	16'h	2167;
19453	:douta	=	16'h	adb8;
19454	:douta	=	16'h	9517;
19455	:douta	=	16'h	5351;
19456	:douta	=	16'h	1083;
19457	:douta	=	16'h	2127;
19458	:douta	=	16'h	3ad0;
19459	:douta	=	16'h	2a90;
19460	:douta	=	16'h	3af2;
19461	:douta	=	16'h	53b6;
19462	:douta	=	16'h	32d1;
19463	:douta	=	16'h	2a70;
19464	:douta	=	16'h	6478;
19465	:douta	=	16'h	3ad0;
19466	:douta	=	16'h	63d4;
19467	:douta	=	16'h	6416;
19468	:douta	=	16'h	7477;
19469	:douta	=	16'h	5330;
19470	:douta	=	16'h	63b3;
19471	:douta	=	16'h	63f3;
19472	:douta	=	16'h	6bd2;
19473	:douta	=	16'h	94b5;
19474	:douta	=	16'h	94d6;
19475	:douta	=	16'h	a536;
19476	:douta	=	16'h	ad35;
19477	:douta	=	16'h	a577;
19478	:douta	=	16'h	8c72;
19479	:douta	=	16'h	8b8a;
19480	:douta	=	16'h	8bab;
19481	:douta	=	16'h	93ac;
19482	:douta	=	16'h	ac6b;
19483	:douta	=	16'h	b4ab;
19484	:douta	=	16'h	c50e;
19485	:douta	=	16'h	d570;
19486	:douta	=	16'h	ddd1;
19487	:douta	=	16'h	d5b0;
19488	:douta	=	16'h	d5b1;
19489	:douta	=	16'h	e674;
19490	:douta	=	16'h	ee96;
19491	:douta	=	16'h	ee96;
19492	:douta	=	16'h	ee96;
19493	:douta	=	16'h	eeb6;
19494	:douta	=	16'h	cd4f;
19495	:douta	=	16'h	f6b6;
19496	:douta	=	16'h	ee96;
19497	:douta	=	16'h	cd70;
19498	:douta	=	16'h	cd6f;
19499	:douta	=	16'h	cd30;
19500	:douta	=	16'h	b4cd;
19501	:douta	=	16'h	a42c;
19502	:douta	=	16'h	834a;
19503	:douta	=	16'h	9c2d;
19504	:douta	=	16'h	a42c;
19505	:douta	=	16'h	a44d;
19506	:douta	=	16'h	b48d;
19507	:douta	=	16'h	c54f;
19508	:douta	=	16'h	cd90;
19509	:douta	=	16'h	d5d1;
19510	:douta	=	16'h	de13;
19511	:douta	=	16'h	de33;
19512	:douta	=	16'h	e674;
19513	:douta	=	16'h	ee75;
19514	:douta	=	16'h	e655;
19515	:douta	=	16'h	e654;
19516	:douta	=	16'h	e654;
19517	:douta	=	16'h	de14;
19518	:douta	=	16'h	ddf3;
19519	:douta	=	16'h	ddf3;
19520	:douta	=	16'h	cd91;
19521	:douta	=	16'h	cd71;
19522	:douta	=	16'h	bcf1;
19523	:douta	=	16'h	b4d1;
19524	:douta	=	16'h	b4b2;
19525	:douta	=	16'h	ac91;
19526	:douta	=	16'h	a4b1;
19527	:douta	=	16'h	7bf2;
19528	:douta	=	16'h	9432;
19529	:douta	=	16'h	8c32;
19530	:douta	=	16'h	7bf2;
19531	:douta	=	16'h	7c12;
19532	:douta	=	16'h	6b70;
19533	:douta	=	16'h	52cd;
19534	:douta	=	16'h	6b70;
19535	:douta	=	16'h	5249;
19536	:douta	=	16'h	59e5;
19537	:douta	=	16'h	b48c;
19538	:douta	=	16'h	ddd0;
19539	:douta	=	16'h	9c2e;
19540	:douta	=	16'h	524b;
19541	:douta	=	16'h	62cc;
19542	:douta	=	16'h	528b;
19543	:douta	=	16'h	3a2b;
19544	:douta	=	16'h	21a8;
19545	:douta	=	16'h	1926;
19546	:douta	=	16'h	1105;
19547	:douta	=	16'h	10a4;
19548	:douta	=	16'h	1904;
19549	:douta	=	16'h	524b;
19550	:douta	=	16'h	2987;
19551	:douta	=	16'h	10c4;
19552	:douta	=	16'h	10a4;
19553	:douta	=	16'h	10c4;
19554	:douta	=	16'h	10c4;
19555	:douta	=	16'h	10c4;
19556	:douta	=	16'h	10c5;
19557	:douta	=	16'h	1905;
19558	:douta	=	16'h	1905;
19559	:douta	=	16'h	18e4;
19560	:douta	=	16'h	0000;
19561	:douta	=	16'h	7412;
19562	:douta	=	16'h	5330;
19563	:douta	=	16'h	9cb4;
19564	:douta	=	16'h	528a;
19565	:douta	=	16'h	c593;
19566	:douta	=	16'h	630b;
19567	:douta	=	16'h	9470;
19568	:douta	=	16'h	8c2e;
19569	:douta	=	16'h	39e8;
19570	:douta	=	16'h	2145;
19571	:douta	=	16'h	62aa;
19572	:douta	=	16'h	2124;
19573	:douta	=	16'h	3166;
19574	:douta	=	16'h	7bad;
19575	:douta	=	16'h	738d;
19576	:douta	=	16'h	52ed;
19577	:douta	=	16'h	8d39;
19578	:douta	=	16'h	8d39;
19579	:douta	=	16'h	957a;
19580	:douta	=	16'h	8d39;
19581	:douta	=	16'h	8518;
19582	:douta	=	16'h	a5db;
19583	:douta	=	16'h	8d59;
19584	:douta	=	16'h	9559;
19585	:douta	=	16'h	8d38;
19586	:douta	=	16'h	8d38;
19587	:douta	=	16'h	9579;
19588	:douta	=	16'h	8d38;
19589	:douta	=	16'h	84d7;
19590	:douta	=	16'h	8d18;
19591	:douta	=	16'h	8cf7;
19592	:douta	=	16'h	84d7;
19593	:douta	=	16'h	84f7;
19594	:douta	=	16'h	9559;
19595	:douta	=	16'h	9579;
19596	:douta	=	16'h	9559;
19597	:douta	=	16'h	7c96;
19598	:douta	=	16'h	84f8;
19599	:douta	=	16'h	8d59;
19600	:douta	=	16'h	957a;
19601	:douta	=	16'h	8519;
19602	:douta	=	16'h	84f8;
19603	:douta	=	16'h	9d9a;
19604	:douta	=	16'h	9579;
19605	:douta	=	16'h	957a;
19606	:douta	=	16'h	9d9a;
19607	:douta	=	16'h	a5da;
19608	:douta	=	16'h	9d99;
19609	:douta	=	16'h	9579;
19610	:douta	=	16'h	9d99;
19611	:douta	=	16'h	a5da;
19612	:douta	=	16'h	9d79;
19613	:douta	=	16'h	a5da;
19614	:douta	=	16'h	9d9a;
19615	:douta	=	16'h	9d99;
19616	:douta	=	16'h	8d18;
19617	:douta	=	16'h	a5da;
19618	:douta	=	16'h	a5fa;
19619	:douta	=	16'h	a5da;
19620	:douta	=	16'h	9d9a;
19621	:douta	=	16'h	b511;
19622	:douta	=	16'h	ee73;
19623	:douta	=	16'h	9c0c;
19624	:douta	=	16'h	0882;
19625	:douta	=	16'h	0863;
19626	:douta	=	16'h	a5db;
19627	:douta	=	16'h	8d17;
19628	:douta	=	16'h	84d8;
19629	:douta	=	16'h	8d38;
19630	:douta	=	16'h	8d39;
19631	:douta	=	16'h	a5ba;
19632	:douta	=	16'h	9d79;
19633	:douta	=	16'h	9538;
19634	:douta	=	16'h	7c75;
19635	:douta	=	16'h	84d7;
19636	:douta	=	16'h	8495;
19637	:douta	=	16'h	7433;
19638	:douta	=	16'h	8495;
19639	:douta	=	16'h	9d57;
19640	:douta	=	16'h	8cb5;
19641	:douta	=	16'h	8cd6;
19642	:douta	=	16'h	94f6;
19643	:douta	=	16'h	7413;
19644	:douta	=	16'h	84f8;
19645	:douta	=	16'h	8539;
19646	:douta	=	16'h	8519;
19647	:douta	=	16'h	7cd8;
19648	:douta	=	16'h	7498;
19649	:douta	=	16'h	8d5a;
19650	:douta	=	16'h	8d7c;
19651	:douta	=	16'h	3a2b;
19652	:douta	=	16'h	2125;
19653	:douta	=	16'h	0884;
19654	:douta	=	16'h	2188;
19655	:douta	=	16'h	2125;
19656	:douta	=	16'h	63f5;
19657	:douta	=	16'h	5bf5;
19658	:douta	=	16'h	6c77;
19659	:douta	=	16'h	7cd8;
19660	:douta	=	16'h	853b;
19661	:douta	=	16'h	855a;
19662	:douta	=	16'h	7d19;
19663	:douta	=	16'h	7d1a;
19664	:douta	=	16'h	74d9;
19665	:douta	=	16'h	6c98;
19666	:douta	=	16'h	8d9c;
19667	:douta	=	16'h	95bc;
19668	:douta	=	16'h	74b8;
19669	:douta	=	16'h	9ddd;
19670	:douta	=	16'h	a63d;
19671	:douta	=	16'h	9dfd;
19672	:douta	=	16'h	95bc;
19673	:douta	=	16'h	6478;
19674	:douta	=	16'h	853a;
19675	:douta	=	16'h	7d3a;
19676	:douta	=	16'h	6cb8;
19677	:douta	=	16'h	5c37;
19678	:douta	=	16'h	6c77;
19679	:douta	=	16'h	6436;
19680	:douta	=	16'h	851a;
19681	:douta	=	16'h	7cb8;
19682	:douta	=	16'h	851a;
19683	:douta	=	16'h	7cb8;
19684	:douta	=	16'h	7498;
19685	:douta	=	16'h	7cd9;
19686	:douta	=	16'h	6437;
19687	:douta	=	16'h	6c57;
19688	:douta	=	16'h	853a;
19689	:douta	=	16'h	853a;
19690	:douta	=	16'h	8d5a;
19691	:douta	=	16'h	7cf9;
19692	:douta	=	16'h	7cd8;
19693	:douta	=	16'h	7cd8;
19694	:douta	=	16'h	95bc;
19695	:douta	=	16'h	8d5a;
19696	:douta	=	16'h	7477;
19697	:douta	=	16'h	6c56;
19698	:douta	=	16'h	6350;
19699	:douta	=	16'h	9d9a;
19700	:douta	=	16'h	8d3a;
19701	:douta	=	16'h	a59a;
19702	:douta	=	16'h	63b2;
19703	:douta	=	16'h	5b93;
19704	:douta	=	16'h	7c55;
19705	:douta	=	16'h	7c55;
19706	:douta	=	16'h	be5d;
19707	:douta	=	16'h	738f;
19708	:douta	=	16'h	5b50;
19709	:douta	=	16'h	7c53;
19710	:douta	=	16'h	8475;
19711	:douta	=	16'h	7413;
19712	:douta	=	16'h	18e4;
19713	:douta	=	16'h	2126;
19714	:douta	=	16'h	2a6f;
19715	:douta	=	16'h	2a4f;
19716	:douta	=	16'h	3af1;
19717	:douta	=	16'h	4bb6;
19718	:douta	=	16'h	3b33;
19719	:douta	=	16'h	2a6f;
19720	:douta	=	16'h	5bd5;
19721	:douta	=	16'h	5bb4;
19722	:douta	=	16'h	7478;
19723	:douta	=	16'h	7cd9;
19724	:douta	=	16'h	74b8;
19725	:douta	=	16'h	5b93;
19726	:douta	=	16'h	6bf4;
19727	:douta	=	16'h	5351;
19728	:douta	=	16'h	73f3;
19729	:douta	=	16'h	94f6;
19730	:douta	=	16'h	8c75;
19731	:douta	=	16'h	8454;
19732	:douta	=	16'h	9c94;
19733	:douta	=	16'h	6b70;
19734	:douta	=	16'h	8b29;
19735	:douta	=	16'h	8bab;
19736	:douta	=	16'h	93cc;
19737	:douta	=	16'h	a40b;
19738	:douta	=	16'h	c4ed;
19739	:douta	=	16'h	cd2e;
19740	:douta	=	16'h	d570;
19741	:douta	=	16'h	ddf1;
19742	:douta	=	16'h	de12;
19743	:douta	=	16'h	ddf2;
19744	:douta	=	16'h	d5b0;
19745	:douta	=	16'h	eeb6;
19746	:douta	=	16'h	e696;
19747	:douta	=	16'h	eeb6;
19748	:douta	=	16'h	e674;
19749	:douta	=	16'h	e654;
19750	:douta	=	16'h	ee95;
19751	:douta	=	16'h	c50e;
19752	:douta	=	16'h	d591;
19753	:douta	=	16'h	cd70;
19754	:douta	=	16'h	b4ad;
19755	:douta	=	16'h	c4ee;
19756	:douta	=	16'h	8b8a;
19757	:douta	=	16'h	8baa;
19758	:douta	=	16'h	9c2c;
19759	:douta	=	16'h	9c0c;
19760	:douta	=	16'h	ac8d;
19761	:douta	=	16'h	c52f;
19762	:douta	=	16'h	cd70;
19763	:douta	=	16'h	d5b1;
19764	:douta	=	16'h	d5f1;
19765	:douta	=	16'h	de13;
19766	:douta	=	16'h	e654;
19767	:douta	=	16'h	e654;
19768	:douta	=	16'h	e654;
19769	:douta	=	16'h	e675;
19770	:douta	=	16'h	ee95;
19771	:douta	=	16'h	de13;
19772	:douta	=	16'h	e634;
19773	:douta	=	16'h	ddf3;
19774	:douta	=	16'h	ddf2;
19775	:douta	=	16'h	d5b2;
19776	:douta	=	16'h	cd52;
19777	:douta	=	16'h	c552;
19778	:douta	=	16'h	acd1;
19779	:douta	=	16'h	a491;
19780	:douta	=	16'h	9c71;
19781	:douta	=	16'h	9c72;
19782	:douta	=	16'h	9c92;
19783	:douta	=	16'h	6371;
19784	:douta	=	16'h	5aef;
19785	:douta	=	16'h	9472;
19786	:douta	=	16'h	738f;
19787	:douta	=	16'h	6b2e;
19788	:douta	=	16'h	73b1;
19789	:douta	=	16'h	73d1;
19790	:douta	=	16'h	41a6;
19791	:douta	=	16'h	7309;
19792	:douta	=	16'h	7288;
19793	:douta	=	16'h	e613;
19794	:douta	=	16'h	d5b0;
19795	:douta	=	16'h	9c2e;
19796	:douta	=	16'h	734d;
19797	:douta	=	16'h	734d;
19798	:douta	=	16'h	62ec;
19799	:douta	=	16'h	5acd;
19800	:douta	=	16'h	4a8c;
19801	:douta	=	16'h	29c9;
19802	:douta	=	16'h	1926;
19803	:douta	=	16'h	2126;
19804	:douta	=	16'h	1906;
19805	:douta	=	16'h	0883;
19806	:douta	=	16'h	0863;
19807	:douta	=	16'h	4a6b;
19808	:douta	=	16'h	0863;
19809	:douta	=	16'h	10e4;
19810	:douta	=	16'h	10a4;
19811	:douta	=	16'h	10e4;
19812	:douta	=	16'h	10c3;
19813	:douta	=	16'h	18a4;
19814	:douta	=	16'h	10c5;
19815	:douta	=	16'h	10a4;
19816	:douta	=	16'h	1926;
19817	:douta	=	16'h	0863;
19818	:douta	=	16'h	52ad;
19819	:douta	=	16'h	6bd2;
19820	:douta	=	16'h	18e5;
19821	:douta	=	16'h	0884;
19822	:douta	=	16'h	4a08;
19823	:douta	=	16'h	7bad;
19824	:douta	=	16'h	9c4e;
19825	:douta	=	16'h	1125;
19826	:douta	=	16'h	1062;
19827	:douta	=	16'h	39e7;
19828	:douta	=	16'h	2966;
19829	:douta	=	16'h	5269;
19830	:douta	=	16'h	6b4d;
19831	:douta	=	16'h	732a;
19832	:douta	=	16'h	5248;
19833	:douta	=	16'h	a5fc;
19834	:douta	=	16'h	8d79;
19835	:douta	=	16'h	8d39;
19836	:douta	=	16'h	84f7;
19837	:douta	=	16'h	957a;
19838	:douta	=	16'h	8d39;
19839	:douta	=	16'h	8d39;
19840	:douta	=	16'h	84f8;
19841	:douta	=	16'h	8d18;
19842	:douta	=	16'h	8d39;
19843	:douta	=	16'h	9d79;
19844	:douta	=	16'h	9559;
19845	:douta	=	16'h	8d38;
19846	:douta	=	16'h	8d38;
19847	:douta	=	16'h	8d38;
19848	:douta	=	16'h	84f8;
19849	:douta	=	16'h	8d18;
19850	:douta	=	16'h	7c96;
19851	:douta	=	16'h	84b7;
19852	:douta	=	16'h	84d7;
19853	:douta	=	16'h	8d59;
19854	:douta	=	16'h	957a;
19855	:douta	=	16'h	8539;
19856	:douta	=	16'h	7cb8;
19857	:douta	=	16'h	6415;
19858	:douta	=	16'h	7cb7;
19859	:douta	=	16'h	84d8;
19860	:douta	=	16'h	8d39;
19861	:douta	=	16'h	84f9;
19862	:douta	=	16'h	8d59;
19863	:douta	=	16'h	959a;
19864	:douta	=	16'h	8d39;
19865	:douta	=	16'h	9d79;
19866	:douta	=	16'h	adda;
19867	:douta	=	16'h	adfa;
19868	:douta	=	16'h	a5ba;
19869	:douta	=	16'h	a5ba;
19870	:douta	=	16'h	a5da;
19871	:douta	=	16'h	b61b;
19872	:douta	=	16'h	adfa;
19873	:douta	=	16'h	9d59;
19874	:douta	=	16'h	9d99;
19875	:douta	=	16'h	9d9a;
19876	:douta	=	16'h	9d79;
19877	:douta	=	16'h	8d39;
19878	:douta	=	16'h	f693;
19879	:douta	=	16'h	ff37;
19880	:douta	=	16'h	3987;
19881	:douta	=	16'h	0043;
19882	:douta	=	16'h	2147;
19883	:douta	=	16'h	8d38;
19884	:douta	=	16'h	8d17;
19885	:douta	=	16'h	9d9a;
19886	:douta	=	16'h	9d99;
19887	:douta	=	16'h	84f8;
19888	:douta	=	16'h	8d39;
19889	:douta	=	16'h	84b6;
19890	:douta	=	16'h	b61b;
19891	:douta	=	16'h	b61a;
19892	:douta	=	16'h	7c33;
19893	:douta	=	16'h	7413;
19894	:douta	=	16'h	7413;
19895	:douta	=	16'h	73f2;
19896	:douta	=	16'h	7412;
19897	:douta	=	16'h	7c55;
19898	:douta	=	16'h	73f3;
19899	:douta	=	16'h	9559;
19900	:douta	=	16'h	957b;
19901	:douta	=	16'h	957b;
19902	:douta	=	16'h	74f9;
19903	:douta	=	16'h	7cd9;
19904	:douta	=	16'h	74b8;
19905	:douta	=	16'h	8d7c;
19906	:douta	=	16'h	5351;
19907	:douta	=	16'h	1905;
19908	:douta	=	16'h	0882;
19909	:douta	=	16'h	29c9;
19910	:douta	=	16'h	10c5;
19911	:douta	=	16'h	3a2b;
19912	:douta	=	16'h	5332;
19913	:douta	=	16'h	5351;
19914	:douta	=	16'h	6bf4;
19915	:douta	=	16'h	7cb8;
19916	:douta	=	16'h	6c77;
19917	:douta	=	16'h	7cf9;
19918	:douta	=	16'h	7cf9;
19919	:douta	=	16'h	84f9;
19920	:douta	=	16'h	7cd9;
19921	:douta	=	16'h	853a;
19922	:douta	=	16'h	853a;
19923	:douta	=	16'h	7cb9;
19924	:douta	=	16'h	8d7b;
19925	:douta	=	16'h	855a;
19926	:douta	=	16'h	7d19;
19927	:douta	=	16'h	857b;
19928	:douta	=	16'h	959b;
19929	:douta	=	16'h	9ddc;
19930	:douta	=	16'h	8d7b;
19931	:douta	=	16'h	8d7b;
19932	:douta	=	16'h	7cf9;
19933	:douta	=	16'h	8d5a;
19934	:douta	=	16'h	95bc;
19935	:douta	=	16'h	8d9c;
19936	:douta	=	16'h	6457;
19937	:douta	=	16'h	5bf6;
19938	:douta	=	16'h	5bd6;
19939	:douta	=	16'h	8d5b;
19940	:douta	=	16'h	6c98;
19941	:douta	=	16'h	7d5a;
19942	:douta	=	16'h	7cd9;
19943	:douta	=	16'h	8d5b;
19944	:douta	=	16'h	7cf9;
19945	:douta	=	16'h	6436;
19946	:douta	=	16'h	6c78;
19947	:douta	=	16'h	8d3a;
19948	:douta	=	16'h	7cd9;
19949	:douta	=	16'h	7cd9;
19950	:douta	=	16'h	853a;
19951	:douta	=	16'h	7cd9;
19952	:douta	=	16'h	7498;
19953	:douta	=	16'h	5bf5;
19954	:douta	=	16'h	632e;
19955	:douta	=	16'h	7c56;
19956	:douta	=	16'h	9538;
19957	:douta	=	16'h	2a2d;
19958	:douta	=	16'h	63d4;
19959	:douta	=	16'h	6c35;
19960	:douta	=	16'h	adda;
19961	:douta	=	16'h	b65c;
19962	:douta	=	16'h	6371;
19963	:douta	=	16'h	0800;
19964	:douta	=	16'h	7cb6;
19965	:douta	=	16'h	84b6;
19966	:douta	=	16'h	7413;
19967	:douta	=	16'h	9537;
19968	:douta	=	16'h	2105;
19969	:douta	=	16'h	1905;
19970	:douta	=	16'h	4334;
19971	:douta	=	16'h	32b1;
19972	:douta	=	16'h	3290;
19973	:douta	=	16'h	3b33;
19974	:douta	=	16'h	4354;
19975	:douta	=	16'h	2a90;
19976	:douta	=	16'h	4b53;
19977	:douta	=	16'h	5bb4;
19978	:douta	=	16'h	63d4;
19979	:douta	=	16'h	7497;
19980	:douta	=	16'h	6c56;
19981	:douta	=	16'h	4310;
19982	:douta	=	16'h	6372;
19983	:douta	=	16'h	7414;
19984	:douta	=	16'h	7414;
19985	:douta	=	16'h	7c54;
19986	:douta	=	16'h	7c33;
19987	:douta	=	16'h	73d2;
19988	:douta	=	16'h	ad77;
19989	:douta	=	16'h	730b;
19990	:douta	=	16'h	9c0b;
19991	:douta	=	16'h	93eb;
19992	:douta	=	16'h	93ab;
19993	:douta	=	16'h	bc8c;
19994	:douta	=	16'h	bcec;
19995	:douta	=	16'h	cd2e;
19996	:douta	=	16'h	d5b1;
19997	:douta	=	16'h	de12;
19998	:douta	=	16'h	de12;
19999	:douta	=	16'h	e654;
20000	:douta	=	16'h	ddf2;
20001	:douta	=	16'h	ee95;
20002	:douta	=	16'h	ee95;
20003	:douta	=	16'h	eed7;
20004	:douta	=	16'h	e675;
20005	:douta	=	16'h	e634;
20006	:douta	=	16'h	ddf3;
20007	:douta	=	16'h	ddf3;
20008	:douta	=	16'h	cd70;
20009	:douta	=	16'h	d5d1;
20010	:douta	=	16'h	c52f;
20011	:douta	=	16'h	ac6c;
20012	:douta	=	16'h	93ca;
20013	:douta	=	16'h	b4ae;
20014	:douta	=	16'h	a42c;
20015	:douta	=	16'h	a42c;
20016	:douta	=	16'h	b48d;
20017	:douta	=	16'h	cd91;
20018	:douta	=	16'h	d5d1;
20019	:douta	=	16'h	d5f2;
20020	:douta	=	16'h	ddf3;
20021	:douta	=	16'h	e654;
20022	:douta	=	16'h	e674;
20023	:douta	=	16'h	e634;
20024	:douta	=	16'h	e675;
20025	:douta	=	16'h	ee75;
20026	:douta	=	16'h	ee75;
20027	:douta	=	16'h	e654;
20028	:douta	=	16'h	e613;
20029	:douta	=	16'h	ddf3;
20030	:douta	=	16'h	ddd2;
20031	:douta	=	16'h	d591;
20032	:douta	=	16'h	c531;
20033	:douta	=	16'h	bd12;
20034	:douta	=	16'h	b4d1;
20035	:douta	=	16'h	a491;
20036	:douta	=	16'h	9452;
20037	:douta	=	16'h	9452;
20038	:douta	=	16'h	9c92;
20039	:douta	=	16'h	6b91;
20040	:douta	=	16'h	4aad;
20041	:douta	=	16'h	5aee;
20042	:douta	=	16'h	8c32;
20043	:douta	=	16'h	7b8f;
20044	:douta	=	16'h	630e;
20045	:douta	=	16'h	4a0a;
20046	:douta	=	16'h	8328;
20047	:douta	=	16'h	ac6c;
20048	:douta	=	16'h	a42a;
20049	:douta	=	16'h	ddd1;
20050	:douta	=	16'h	ddd2;
20051	:douta	=	16'h	a44d;
20052	:douta	=	16'h	8bae;
20053	:douta	=	16'h	7b6e;
20054	:douta	=	16'h	630d;
20055	:douta	=	16'h	630d;
20056	:douta	=	16'h	5aee;
20057	:douta	=	16'h	2a2b;
20058	:douta	=	16'h	2167;
20059	:douta	=	16'h	2126;
20060	:douta	=	16'h	2126;
20061	:douta	=	16'h	18e5;
20062	:douta	=	16'h	10a4;
20063	:douta	=	16'h	2947;
20064	:douta	=	16'h	29a8;
20065	:douta	=	16'h	0863;
20066	:douta	=	16'h	10a3;
20067	:douta	=	16'h	10c3;
20068	:douta	=	16'h	10a4;
20069	:douta	=	16'h	10a4;
20070	:douta	=	16'h	10c5;
20071	:douta	=	16'h	10c4;
20072	:douta	=	16'h	10a4;
20073	:douta	=	16'h	29c9;
20074	:douta	=	16'h	0042;
20075	:douta	=	16'h	1905;
20076	:douta	=	16'h	10e5;
20077	:douta	=	16'h	1926;
20078	:douta	=	16'h	2146;
20079	:douta	=	16'h	83cd;
20080	:douta	=	16'h	d655;
20081	:douta	=	16'h	6b0c;
20082	:douta	=	16'h	a490;
20083	:douta	=	16'h	6b0b;
20084	:douta	=	16'h	4a49;
20085	:douta	=	16'h	4a49;
20086	:douta	=	16'h	5acb;
20087	:douta	=	16'h	9c2e;
20088	:douta	=	16'h	62cb;
20089	:douta	=	16'h	7433;
20090	:douta	=	16'h	a5fc;
20091	:douta	=	16'h	9559;
20092	:douta	=	16'h	9559;
20093	:douta	=	16'h	9559;
20094	:douta	=	16'h	8518;
20095	:douta	=	16'h	957a;
20096	:douta	=	16'h	84f8;
20097	:douta	=	16'h	8d18;
20098	:douta	=	16'h	8d18;
20099	:douta	=	16'h	8d17;
20100	:douta	=	16'h	8d17;
20101	:douta	=	16'h	8d17;
20102	:douta	=	16'h	8d38;
20103	:douta	=	16'h	9538;
20104	:douta	=	16'h	84d7;
20105	:douta	=	16'h	84f7;
20106	:douta	=	16'h	8d18;
20107	:douta	=	16'h	84d7;
20108	:douta	=	16'h	8cf8;
20109	:douta	=	16'h	84d7;
20110	:douta	=	16'h	84d7;
20111	:douta	=	16'h	84d7;
20112	:douta	=	16'h	8d7a;
20113	:douta	=	16'h	8519;
20114	:douta	=	16'h	84d8;
20115	:douta	=	16'h	74b7;
20116	:douta	=	16'h	8d5a;
20117	:douta	=	16'h	8518;
20118	:douta	=	16'h	8d39;
20119	:douta	=	16'h	8d59;
20120	:douta	=	16'h	9dbb;
20121	:douta	=	16'h	9579;
20122	:douta	=	16'h	a5da;
20123	:douta	=	16'h	adfb;
20124	:douta	=	16'h	a5ba;
20125	:douta	=	16'h	a5fa;
20126	:douta	=	16'h	9d9a;
20127	:douta	=	16'h	959a;
20128	:douta	=	16'h	9d79;
20129	:douta	=	16'h	9d99;
20130	:douta	=	16'h	9579;
20131	:douta	=	16'h	a5da;
20132	:douta	=	16'h	a5ba;
20133	:douta	=	16'h	8d59;
20134	:douta	=	16'h	de13;
20135	:douta	=	16'h	ff37;
20136	:douta	=	16'h	ac0d;
20137	:douta	=	16'h	18e7;
20138	:douta	=	16'h	0001;
20139	:douta	=	16'h	2168;
20140	:douta	=	16'h	ae1b;
20141	:douta	=	16'h	8d58;
20142	:douta	=	16'h	9d9a;
20143	:douta	=	16'h	9d9a;
20144	:douta	=	16'h	9d79;
20145	:douta	=	16'h	9d78;
20146	:douta	=	16'h	8cf6;
20147	:douta	=	16'h	a598;
20148	:douta	=	16'h	9537;
20149	:douta	=	16'h	a558;
20150	:douta	=	16'h	8475;
20151	:douta	=	16'h	634f;
20152	:douta	=	16'h	73d2;
20153	:douta	=	16'h	94f7;
20154	:douta	=	16'h	7c95;
20155	:douta	=	16'h	7cb7;
20156	:douta	=	16'h	7cd8;
20157	:douta	=	16'h	7d19;
20158	:douta	=	16'h	7cf9;
20159	:douta	=	16'h	74d9;
20160	:douta	=	16'h	74b9;
20161	:douta	=	16'h	5bb3;
20162	:douta	=	16'h	2146;
20163	:douta	=	16'h	18c3;
20164	:douta	=	16'h	21a8;
20165	:douta	=	16'h	2187;
20166	:douta	=	16'h	0884;
20167	:douta	=	16'h	7cb8;
20168	:douta	=	16'h	6415;
20169	:douta	=	16'h	53b3;
20170	:douta	=	16'h	84b8;
20171	:douta	=	16'h	6c98;
20172	:douta	=	16'h	6c36;
20173	:douta	=	16'h	851a;
20174	:douta	=	16'h	8d3a;
20175	:douta	=	16'h	8539;
20176	:douta	=	16'h	8d5a;
20177	:douta	=	16'h	8d7b;
20178	:douta	=	16'h	8519;
20179	:douta	=	16'h	8519;
20180	:douta	=	16'h	7cd9;
20181	:douta	=	16'h	8d7b;
20182	:douta	=	16'h	851a;
20183	:douta	=	16'h	8d5b;
20184	:douta	=	16'h	8d5a;
20185	:douta	=	16'h	ae5d;
20186	:douta	=	16'h	8d5b;
20187	:douta	=	16'h	7d3a;
20188	:douta	=	16'h	7cf9;
20189	:douta	=	16'h	853a;
20190	:douta	=	16'h	8d7b;
20191	:douta	=	16'h	853a;
20192	:douta	=	16'h	95bd;
20193	:douta	=	16'h	74b9;
20194	:douta	=	16'h	5bf6;
20195	:douta	=	16'h	7d19;
20196	:douta	=	16'h	7498;
20197	:douta	=	16'h	74d9;
20198	:douta	=	16'h	851a;
20199	:douta	=	16'h	74d9;
20200	:douta	=	16'h	8d5a;
20201	:douta	=	16'h	853a;
20202	:douta	=	16'h	7cd9;
20203	:douta	=	16'h	6c57;
20204	:douta	=	16'h	7cd9;
20205	:douta	=	16'h	7cd8;
20206	:douta	=	16'h	7cd8;
20207	:douta	=	16'h	6c37;
20208	:douta	=	16'h	74d9;
20209	:douta	=	16'h	6371;
20210	:douta	=	16'h	5353;
20211	:douta	=	16'h	a5fc;
20212	:douta	=	16'h	9d79;
20213	:douta	=	16'h	84f8;
20214	:douta	=	16'h	4b31;
20215	:douta	=	16'h	63d2;
20216	:douta	=	16'h	84d7;
20217	:douta	=	16'h	6457;
20218	:douta	=	16'h	49e9;
20219	:douta	=	16'h	1881;
20220	:douta	=	16'h	9517;
20221	:douta	=	16'h	6bd1;
20222	:douta	=	16'h	6391;
20223	:douta	=	16'h	7c75;
20224	:douta	=	16'h	2905;
20225	:douta	=	16'h	18a4;
20226	:douta	=	16'h	29ea;
20227	:douta	=	16'h	2250;
20228	:douta	=	16'h	3ad1;
20229	:douta	=	16'h	4374;
20230	:douta	=	16'h	32d2;
20231	:douta	=	16'h	32d1;
20232	:douta	=	16'h	53b5;
20233	:douta	=	16'h	5394;
20234	:douta	=	16'h	5b93;
20235	:douta	=	16'h	5bb4;
20236	:douta	=	16'h	6c56;
20237	:douta	=	16'h	6c36;
20238	:douta	=	16'h	7c14;
20239	:douta	=	16'h	7435;
20240	:douta	=	16'h	7c76;
20241	:douta	=	16'h	8454;
20242	:douta	=	16'h	9d17;
20243	:douta	=	16'h	94b5;
20244	:douta	=	16'h	734e;
20245	:douta	=	16'h	93ca;
20246	:douta	=	16'h	93aa;
20247	:douta	=	16'h	a42c;
20248	:douta	=	16'h	ac4b;
20249	:douta	=	16'h	c4cd;
20250	:douta	=	16'h	cd2e;
20251	:douta	=	16'h	d570;
20252	:douta	=	16'h	ddd2;
20253	:douta	=	16'h	e654;
20254	:douta	=	16'h	e674;
20255	:douta	=	16'h	eed7;
20256	:douta	=	16'h	f6f7;
20257	:douta	=	16'h	e654;
20258	:douta	=	16'h	e613;
20259	:douta	=	16'h	ddd2;
20260	:douta	=	16'h	e695;
20261	:douta	=	16'h	de13;
20262	:douta	=	16'h	d5b1;
20263	:douta	=	16'h	c52f;
20264	:douta	=	16'h	cd90;
20265	:douta	=	16'h	c52f;
20266	:douta	=	16'h	bcce;
20267	:douta	=	16'h	8b69;
20268	:douta	=	16'h	ac6d;
20269	:douta	=	16'h	ac6d;
20270	:douta	=	16'h	ac8d;
20271	:douta	=	16'h	b4ed;
20272	:douta	=	16'h	c50e;
20273	:douta	=	16'h	d5f2;
20274	:douta	=	16'h	de13;
20275	:douta	=	16'h	e655;
20276	:douta	=	16'h	e654;
20277	:douta	=	16'h	e654;
20278	:douta	=	16'h	ee96;
20279	:douta	=	16'h	eeb6;
20280	:douta	=	16'h	ee75;
20281	:douta	=	16'h	e675;
20282	:douta	=	16'h	e634;
20283	:douta	=	16'h	e654;
20284	:douta	=	16'h	e654;
20285	:douta	=	16'h	ddd2;
20286	:douta	=	16'h	d591;
20287	:douta	=	16'h	bd10;
20288	:douta	=	16'h	ac91;
20289	:douta	=	16'h	9c51;
20290	:douta	=	16'h	9c52;
20291	:douta	=	16'h	9c72;
20292	:douta	=	16'h	9c92;
20293	:douta	=	16'h	8412;
20294	:douta	=	16'h	8431;
20295	:douta	=	16'h	73d1;
20296	:douta	=	16'h	5aee;
20297	:douta	=	16'h	31ea;
20298	:douta	=	16'h	39ea;
20299	:douta	=	16'h	4a6b;
20300	:douta	=	16'h	5a26;
20301	:douta	=	16'h	ac2c;
20302	:douta	=	16'h	93cb;
20303	:douta	=	16'h	cd2e;
20304	:douta	=	16'h	e5f2;
20305	:douta	=	16'h	e634;
20306	:douta	=	16'h	d58f;
20307	:douta	=	16'h	b48d;
20308	:douta	=	16'h	93ac;
20309	:douta	=	16'h	7b6e;
20310	:douta	=	16'h	630d;
20311	:douta	=	16'h	630e;
20312	:douta	=	16'h	630e;
20313	:douta	=	16'h	52ee;
20314	:douta	=	16'h	3a4c;
20315	:douta	=	16'h	322c;
20316	:douta	=	16'h	322b;
20317	:douta	=	16'h	29a9;
20318	:douta	=	16'h	2988;
20319	:douta	=	16'h	1906;
20320	:douta	=	16'h	1084;
20321	:douta	=	16'h	42ad;
20322	:douta	=	16'h	0883;
20323	:douta	=	16'h	10a3;
20324	:douta	=	16'h	10c4;
20325	:douta	=	16'h	18e5;
20326	:douta	=	16'h	1905;
20327	:douta	=	16'h	10a4;
20328	:douta	=	16'h	10c5;
20329	:douta	=	16'h	1083;
20330	:douta	=	16'h	2146;
20331	:douta	=	16'h	29a8;
20332	:douta	=	16'h	10c5;
20333	:douta	=	16'h	1926;
20334	:douta	=	16'h	2126;
20335	:douta	=	16'h	1926;
20336	:douta	=	16'h	2167;
20337	:douta	=	16'h	d633;
20338	:douta	=	16'h	8c6f;
20339	:douta	=	16'h	8c2e;
20340	:douta	=	16'h	1063;
20341	:douta	=	16'h	10a4;
20342	:douta	=	16'h	3986;
20343	:douta	=	16'h	31a6;
20344	:douta	=	16'h	6b0b;
20345	:douta	=	16'h	5aaa;
20346	:douta	=	16'h	6391;
20347	:douta	=	16'h	7cb7;
20348	:douta	=	16'h	7496;
20349	:douta	=	16'h	9579;
20350	:douta	=	16'h	9d7a;
20351	:douta	=	16'h	9559;
20352	:douta	=	16'h	9579;
20353	:douta	=	16'h	9579;
20354	:douta	=	16'h	8d38;
20355	:douta	=	16'h	8d38;
20356	:douta	=	16'h	9579;
20357	:douta	=	16'h	8d38;
20358	:douta	=	16'h	8d38;
20359	:douta	=	16'h	8d18;
20360	:douta	=	16'h	84f8;
20361	:douta	=	16'h	8d39;
20362	:douta	=	16'h	9d99;
20363	:douta	=	16'h	8d58;
20364	:douta	=	16'h	8d18;
20365	:douta	=	16'h	9559;
20366	:douta	=	16'h	8d18;
20367	:douta	=	16'h	9559;
20368	:douta	=	16'h	84d8;
20369	:douta	=	16'h	8518;
20370	:douta	=	16'h	8d18;
20371	:douta	=	16'h	9559;
20372	:douta	=	16'h	9d9a;
20373	:douta	=	16'h	957a;
20374	:douta	=	16'h	8d39;
20375	:douta	=	16'h	8518;
20376	:douta	=	16'h	8d18;
20377	:douta	=	16'h	8d39;
20378	:douta	=	16'h	957a;
20379	:douta	=	16'h	9d9a;
20380	:douta	=	16'h	9559;
20381	:douta	=	16'h	8d18;
20382	:douta	=	16'h	8d39;
20383	:douta	=	16'h	8d39;
20384	:douta	=	16'h	9d9a;
20385	:douta	=	16'h	9d9a;
20386	:douta	=	16'h	9d9a;
20387	:douta	=	16'h	9d9a;
20388	:douta	=	16'h	9d79;
20389	:douta	=	16'h	9d99;
20390	:douta	=	16'h	8d5a;
20391	:douta	=	16'h	ad34;
20392	:douta	=	16'h	ff98;
20393	:douta	=	16'h	e590;
20394	:douta	=	16'h	29eb;
20395	:douta	=	16'h	1106;
20396	:douta	=	16'h	0043;
20397	:douta	=	16'h	7cb7;
20398	:douta	=	16'h	a5fb;
20399	:douta	=	16'h	9d79;
20400	:douta	=	16'h	9538;
20401	:douta	=	16'h	9558;
20402	:douta	=	16'h	9d58;
20403	:douta	=	16'h	9d58;
20404	:douta	=	16'h	8c94;
20405	:douta	=	16'h	94f6;
20406	:douta	=	16'h	8473;
20407	:douta	=	16'h	9d16;
20408	:douta	=	16'h	9537;
20409	:douta	=	16'h	7c35;
20410	:douta	=	16'h	73f4;
20411	:douta	=	16'h	6cb8;
20412	:douta	=	16'h	53f5;
20413	:douta	=	16'h	6457;
20414	:douta	=	16'h	753c;
20415	:douta	=	16'h	7d5c;
20416	:douta	=	16'h	39ea;
20417	:douta	=	16'h	2125;
20418	:douta	=	16'h	20e5;
20419	:douta	=	16'h	322c;
20420	:douta	=	16'h	1927;
20421	:douta	=	16'h	1107;
20422	:douta	=	16'h	7d1a;
20423	:douta	=	16'h	7d3a;
20424	:douta	=	16'h	853a;
20425	:douta	=	16'h	8d7b;
20426	:douta	=	16'h	853a;
20427	:douta	=	16'h	8d5a;
20428	:douta	=	16'h	84f9;
20429	:douta	=	16'h	6415;
20430	:douta	=	16'h	6c36;
20431	:douta	=	16'h	7498;
20432	:douta	=	16'h	853a;
20433	:douta	=	16'h	855a;
20434	:douta	=	16'h	853a;
20435	:douta	=	16'h	853a;
20436	:douta	=	16'h	8519;
20437	:douta	=	16'h	7498;
20438	:douta	=	16'h	8519;
20439	:douta	=	16'h	8d5a;
20440	:douta	=	16'h	8d7b;
20441	:douta	=	16'h	8519;
20442	:douta	=	16'h	851a;
20443	:douta	=	16'h	855a;
20444	:douta	=	16'h	8d7b;
20445	:douta	=	16'h	853a;
20446	:douta	=	16'h	853a;
20447	:douta	=	16'h	853b;
20448	:douta	=	16'h	853a;
20449	:douta	=	16'h	74d9;
20450	:douta	=	16'h	7cfa;
20451	:douta	=	16'h	855a;
20452	:douta	=	16'h	5394;
20453	:douta	=	16'h	5c16;
20454	:douta	=	16'h	8d7b;
20455	:douta	=	16'h	7cd9;
20456	:douta	=	16'h	959b;
20457	:douta	=	16'h	7cf9;
20458	:douta	=	16'h	8d5a;
20459	:douta	=	16'h	7498;
20460	:douta	=	16'h	74d8;
20461	:douta	=	16'h	6457;
20462	:douta	=	16'h	74d8;
20463	:douta	=	16'h	6cda;
20464	:douta	=	16'h	72cb;
20465	:douta	=	16'h	630e;
20466	:douta	=	16'h	a5fb;
20467	:douta	=	16'h	7414;
20468	:douta	=	16'h	5351;
20469	:douta	=	16'h	5310;
20470	:douta	=	16'h	7c76;
20471	:douta	=	16'h	7cb7;
20472	:douta	=	16'h	84f8;
20473	:douta	=	16'h	b69f;
20474	:douta	=	16'h	0800;
20475	:douta	=	16'h	5330;
20476	:douta	=	16'h	6c14;
20477	:douta	=	16'h	7434;
20478	:douta	=	16'h	7454;
20479	:douta	=	16'h	7c95;
20480	:douta	=	16'h	2925;
20481	:douta	=	16'h	18a3;
20482	:douta	=	16'h	29a9;
20483	:douta	=	16'h	4bd6;
20484	:douta	=	16'h	222e;
20485	:douta	=	16'h	32b1;
20486	:douta	=	16'h	3312;
20487	:douta	=	16'h	220d;
20488	:douta	=	16'h	3ad1;
20489	:douta	=	16'h	6416;
20490	:douta	=	16'h	5b94;
20491	:douta	=	16'h	7cb8;
20492	:douta	=	16'h	7498;
20493	:douta	=	16'h	53b4;
20494	:douta	=	16'h	324c;
20495	:douta	=	16'h	5b92;
20496	:douta	=	16'h	6c14;
20497	:douta	=	16'h	8c96;
20498	:douta	=	16'h	8c94;
20499	:douta	=	16'h	94d4;
20500	:douta	=	16'h	62a9;
20501	:douta	=	16'h	9bea;
20502	:douta	=	16'h	93cb;
20503	:douta	=	16'h	ac4b;
20504	:douta	=	16'h	b48b;
20505	:douta	=	16'h	c50d;
20506	:douta	=	16'h	cd4f;
20507	:douta	=	16'h	d590;
20508	:douta	=	16'h	ddf2;
20509	:douta	=	16'h	e654;
20510	:douta	=	16'h	ee96;
20511	:douta	=	16'h	eeb6;
20512	:douta	=	16'h	eeb6;
20513	:douta	=	16'h	eeb6;
20514	:douta	=	16'h	e695;
20515	:douta	=	16'h	de13;
20516	:douta	=	16'h	e634;
20517	:douta	=	16'h	e613;
20518	:douta	=	16'h	d570;
20519	:douta	=	16'h	cd4f;
20520	:douta	=	16'h	c52e;
20521	:douta	=	16'h	c50e;
20522	:douta	=	16'h	938a;
20523	:douta	=	16'h	b48d;
20524	:douta	=	16'h	a44c;
20525	:douta	=	16'h	ac8d;
20526	:douta	=	16'h	bcee;
20527	:douta	=	16'h	bced;
20528	:douta	=	16'h	d591;
20529	:douta	=	16'h	de33;
20530	:douta	=	16'h	e634;
20531	:douta	=	16'h	e675;
20532	:douta	=	16'h	e675;
20533	:douta	=	16'h	e654;
20534	:douta	=	16'h	ee96;
20535	:douta	=	16'h	ee96;
20536	:douta	=	16'h	e654;
20537	:douta	=	16'h	e654;
20538	:douta	=	16'h	e613;
20539	:douta	=	16'h	de13;
20540	:douta	=	16'h	e613;
20541	:douta	=	16'h	d5b2;
20542	:douta	=	16'h	d592;
20543	:douta	=	16'h	bcef;
20544	:douta	=	16'h	9c51;
20545	:douta	=	16'h	9c51;
20546	:douta	=	16'h	9c71;
20547	:douta	=	16'h	9c72;
20548	:douta	=	16'h	9452;
20549	:douta	=	16'h	8c32;
20550	:douta	=	16'h	8432;
20551	:douta	=	16'h	7bf2;
20552	:douta	=	16'h	6b6f;
20553	:douta	=	16'h	5aee;
20554	:douta	=	16'h	2988;
20555	:douta	=	16'h	20e6;
20556	:douta	=	16'h	82e7;
20557	:douta	=	16'h	c50e;
20558	:douta	=	16'h	ac6c;
20559	:douta	=	16'h	ddb1;
20560	:douta	=	16'h	e654;
20561	:douta	=	16'h	e612;
20562	:douta	=	16'h	ddd1;
20563	:douta	=	16'h	bcac;
20564	:douta	=	16'h	9bed;
20565	:douta	=	16'h	838e;
20566	:douta	=	16'h	632d;
20567	:douta	=	16'h	5b0d;
20568	:douta	=	16'h	6b6f;
20569	:douta	=	16'h	632f;
20570	:douta	=	16'h	5310;
20571	:douta	=	16'h	42af;
20572	:douta	=	16'h	42ae;
20573	:douta	=	16'h	3a2c;
20574	:douta	=	16'h	29cb;
20575	:douta	=	16'h	2168;
20576	:douta	=	16'h	10c4;
20577	:douta	=	16'h	0884;
20578	:douta	=	16'h	428d;
20579	:douta	=	16'h	10a4;
20580	:douta	=	16'h	18e5;
20581	:douta	=	16'h	10c5;
20582	:douta	=	16'h	10e5;
20583	:douta	=	16'h	10a4;
20584	:douta	=	16'h	10a4;
20585	:douta	=	16'h	18c5;
20586	:douta	=	16'h	10a3;
20587	:douta	=	16'h	1905;
20588	:douta	=	16'h	10e5;
20589	:douta	=	16'h	0863;
20590	:douta	=	16'h	1926;
20591	:douta	=	16'h	1926;
20592	:douta	=	16'h	08c5;
20593	:douta	=	16'h	738d;
20594	:douta	=	16'h	52aa;
20595	:douta	=	16'h	c5d4;
20596	:douta	=	16'h	a4d2;
20597	:douta	=	16'h	6b4d;
20598	:douta	=	16'h	9c2f;
20599	:douta	=	16'h	630b;
20600	:douta	=	16'h	20c3;
20601	:douta	=	16'h	39a8;
20602	:douta	=	16'h	3988;
20603	:douta	=	16'h	9dbb;
20604	:douta	=	16'h	84d7;
20605	:douta	=	16'h	7cd7;
20606	:douta	=	16'h	9559;
20607	:douta	=	16'h	9d9a;
20608	:douta	=	16'h	9dba;
20609	:douta	=	16'h	a5db;
20610	:douta	=	16'h	9dba;
20611	:douta	=	16'h	84f7;
20612	:douta	=	16'h	8d39;
20613	:douta	=	16'h	8d18;
20614	:douta	=	16'h	84f8;
20615	:douta	=	16'h	84f8;
20616	:douta	=	16'h	84f8;
20617	:douta	=	16'h	84f8;
20618	:douta	=	16'h	8d38;
20619	:douta	=	16'h	8d39;
20620	:douta	=	16'h	9d7a;
20621	:douta	=	16'h	8d59;
20622	:douta	=	16'h	8d39;
20623	:douta	=	16'h	84f8;
20624	:douta	=	16'h	8539;
20625	:douta	=	16'h	84f8;
20626	:douta	=	16'h	8d18;
20627	:douta	=	16'h	7cb7;
20628	:douta	=	16'h	8d39;
20629	:douta	=	16'h	957a;
20630	:douta	=	16'h	8d39;
20631	:douta	=	16'h	957a;
20632	:douta	=	16'h	9559;
20633	:douta	=	16'h	84f8;
20634	:douta	=	16'h	84d7;
20635	:douta	=	16'h	8d38;
20636	:douta	=	16'h	9dba;
20637	:douta	=	16'h	9dba;
20638	:douta	=	16'h	84f8;
20639	:douta	=	16'h	8517;
20640	:douta	=	16'h	8d39;
20641	:douta	=	16'h	9559;
20642	:douta	=	16'h	a5da;
20643	:douta	=	16'h	957a;
20644	:douta	=	16'h	8d39;
20645	:douta	=	16'h	9d99;
20646	:douta	=	16'h	9dbb;
20647	:douta	=	16'h	8519;
20648	:douta	=	16'h	f6b4;
20649	:douta	=	16'h	ff14;
20650	:douta	=	16'h	426d;
20651	:douta	=	16'h	4b0f;
20652	:douta	=	16'h	0001;
20653	:douta	=	16'h	08c5;
20654	:douta	=	16'h	3aae;
20655	:douta	=	16'h	9dbb;
20656	:douta	=	16'h	a5fb;
20657	:douta	=	16'h	8d18;
20658	:douta	=	16'h	9d79;
20659	:douta	=	16'h	9517;
20660	:douta	=	16'h	a557;
20661	:douta	=	16'h	9d16;
20662	:douta	=	16'h	8c93;
20663	:douta	=	16'h	8493;
20664	:douta	=	16'h	7c74;
20665	:douta	=	16'h	7cb8;
20666	:douta	=	16'h	7d3a;
20667	:douta	=	16'h	5c37;
20668	:douta	=	16'h	5c58;
20669	:douta	=	16'h	6cda;
20670	:douta	=	16'h	4b94;
20671	:douta	=	16'h	322c;
20672	:douta	=	16'h	2904;
20673	:douta	=	16'h	2125;
20674	:douta	=	16'h	3a8d;
20675	:douta	=	16'h	2189;
20676	:douta	=	16'h	4311;
20677	:douta	=	16'h	1126;
20678	:douta	=	16'h	7cfa;
20679	:douta	=	16'h	5c15;
20680	:douta	=	16'h	7d19;
20681	:douta	=	16'h	95bc;
20682	:douta	=	16'h	95bb;
20683	:douta	=	16'h	8d7a;
20684	:douta	=	16'h	959b;
20685	:douta	=	16'h	8d5a;
20686	:douta	=	16'h	8d1a;
20687	:douta	=	16'h	53b4;
20688	:douta	=	16'h	7497;
20689	:douta	=	16'h	6c16;
20690	:douta	=	16'h	8d5a;
20691	:douta	=	16'h	959c;
20692	:douta	=	16'h	853a;
20693	:douta	=	16'h	7cd9;
20694	:douta	=	16'h	7498;
20695	:douta	=	16'h	7498;
20696	:douta	=	16'h	84f9;
20697	:douta	=	16'h	8d5a;
20698	:douta	=	16'h	8d7b;
20699	:douta	=	16'h	959c;
20700	:douta	=	16'h	8d7c;
20701	:douta	=	16'h	7d1a;
20702	:douta	=	16'h	8d7b;
20703	:douta	=	16'h	7cf9;
20704	:douta	=	16'h	853a;
20705	:douta	=	16'h	959c;
20706	:douta	=	16'h	853a;
20707	:douta	=	16'h	95bc;
20708	:douta	=	16'h	6457;
20709	:douta	=	16'h	4332;
20710	:douta	=	16'h	7498;
20711	:douta	=	16'h	8d5b;
20712	:douta	=	16'h	74b8;
20713	:douta	=	16'h	6c57;
20714	:douta	=	16'h	6c78;
20715	:douta	=	16'h	7d3a;
20716	:douta	=	16'h	7cf9;
20717	:douta	=	16'h	74b9;
20718	:douta	=	16'h	53d6;
20719	:douta	=	16'h	3af1;
20720	:douta	=	16'h	736f;
20721	:douta	=	16'h	7cd9;
20722	:douta	=	16'h	5330;
20723	:douta	=	16'h	9d9a;
20724	:douta	=	16'h	8cf8;
20725	:douta	=	16'h	8496;
20726	:douta	=	16'h	8d18;
20727	:douta	=	16'h	63f4;
20728	:douta	=	16'h	63d4;
20729	:douta	=	16'h	63f3;
20730	:douta	=	16'h	2946;
20731	:douta	=	16'h	7cd8;
20732	:douta	=	16'h	adfa;
20733	:douta	=	16'h	a599;
20734	:douta	=	16'h	5b72;
20735	:douta	=	16'h	6c13;
20736	:douta	=	16'h	2945;
20737	:douta	=	16'h	1062;
20738	:douta	=	16'h	2146;
20739	:douta	=	16'h	4394;
20740	:douta	=	16'h	21cc;
20741	:douta	=	16'h	32b0;
20742	:douta	=	16'h	2ab1;
20743	:douta	=	16'h	2a4f;
20744	:douta	=	16'h	4333;
20745	:douta	=	16'h	6436;
20746	:douta	=	16'h	5393;
20747	:douta	=	16'h	5393;
20748	:douta	=	16'h	6415;
20749	:douta	=	16'h	63d4;
20750	:douta	=	16'h	6bd3;
20751	:douta	=	16'h	6bd3;
20752	:douta	=	16'h	9d58;
20753	:douta	=	16'h	7c55;
20754	:douta	=	16'h	a577;
20755	:douta	=	16'h	732c;
20756	:douta	=	16'h	8b8a;
20757	:douta	=	16'h	ac4c;
20758	:douta	=	16'h	b48b;
20759	:douta	=	16'h	ac6c;
20760	:douta	=	16'h	d54f;
20761	:douta	=	16'h	cd4f;
20762	:douta	=	16'h	d58f;
20763	:douta	=	16'h	d5d0;
20764	:douta	=	16'h	ee75;
20765	:douta	=	16'h	eeb6;
20766	:douta	=	16'h	ee95;
20767	:douta	=	16'h	eeb6;
20768	:douta	=	16'h	eeb7;
20769	:douta	=	16'h	ee75;
20770	:douta	=	16'h	ee75;
20771	:douta	=	16'h	e654;
20772	:douta	=	16'h	ddd2;
20773	:douta	=	16'h	d591;
20774	:douta	=	16'h	c4ef;
20775	:douta	=	16'h	b46c;
20776	:douta	=	16'h	b48e;
20777	:douta	=	16'h	8b69;
20778	:douta	=	16'h	a44c;
20779	:douta	=	16'h	9c2b;
20780	:douta	=	16'h	b4ad;
20781	:douta	=	16'h	bcee;
20782	:douta	=	16'h	c52e;
20783	:douta	=	16'h	cd6f;
20784	:douta	=	16'h	d5b2;
20785	:douta	=	16'h	e655;
20786	:douta	=	16'h	e655;
20787	:douta	=	16'h	e675;
20788	:douta	=	16'h	eeb6;
20789	:douta	=	16'h	ee96;
20790	:douta	=	16'h	e675;
20791	:douta	=	16'h	e675;
20792	:douta	=	16'h	e675;
20793	:douta	=	16'h	e654;
20794	:douta	=	16'h	e613;
20795	:douta	=	16'h	ddd2;
20796	:douta	=	16'h	d5b1;
20797	:douta	=	16'h	cd90;
20798	:douta	=	16'h	cd50;
20799	:douta	=	16'h	a450;
20800	:douta	=	16'h	9431;
20801	:douta	=	16'h	8c11;
20802	:douta	=	16'h	8412;
20803	:douta	=	16'h	7bd1;
20804	:douta	=	16'h	7bb0;
20805	:douta	=	16'h	7b6f;
20806	:douta	=	16'h	7b6f;
20807	:douta	=	16'h	630e;
20808	:douta	=	16'h	630e;
20809	:douta	=	16'h	524a;
20810	:douta	=	16'h	5a27;
20811	:douta	=	16'h	9389;
20812	:douta	=	16'h	93cc;
20813	:douta	=	16'h	938b;
20814	:douta	=	16'h	cd70;
20815	:douta	=	16'h	ddf2;
20816	:douta	=	16'h	e613;
20817	:douta	=	16'h	e613;
20818	:douta	=	16'h	d58f;
20819	:douta	=	16'h	d52f;
20820	:douta	=	16'h	a42d;
20821	:douta	=	16'h	a40e;
20822	:douta	=	16'h	7b6e;
20823	:douta	=	16'h	6b2e;
20824	:douta	=	16'h	632e;
20825	:douta	=	16'h	632f;
20826	:douta	=	16'h	5b50;
20827	:douta	=	16'h	5330;
20828	:douta	=	16'h	5310;
20829	:douta	=	16'h	42cf;
20830	:douta	=	16'h	42ae;
20831	:douta	=	16'h	322c;
20832	:douta	=	16'h	29ca;
20833	:douta	=	16'h	2168;
20834	:douta	=	16'h	0884;
20835	:douta	=	16'h	424c;
20836	:douta	=	16'h	1906;
20837	:douta	=	16'h	10a4;
20838	:douta	=	16'h	10a4;
20839	:douta	=	16'h	18e5;
20840	:douta	=	16'h	18e5;
20841	:douta	=	16'h	10e4;
20842	:douta	=	16'h	10c5;
20843	:douta	=	16'h	1905;
20844	:douta	=	16'h	10a3;
20845	:douta	=	16'h	1925;
20846	:douta	=	16'h	10e4;
20847	:douta	=	16'h	2126;
20848	:douta	=	16'h	1927;
20849	:douta	=	16'h	0043;
20850	:douta	=	16'h	a491;
20851	:douta	=	16'h	2167;
20852	:douta	=	16'h	a513;
20853	:douta	=	16'h	2967;
20854	:douta	=	16'h	6b6d;
20855	:douta	=	16'h	2166;
20856	:douta	=	16'h	6b2b;
20857	:douta	=	16'h	62cb;
20858	:douta	=	16'h	7bce;
20859	:douta	=	16'h	4aae;
20860	:douta	=	16'h	95bb;
20861	:douta	=	16'h	8d18;
20862	:douta	=	16'h	8518;
20863	:douta	=	16'h	84d7;
20864	:douta	=	16'h	84d7;
20865	:douta	=	16'h	7cb6;
20866	:douta	=	16'h	9559;
20867	:douta	=	16'h	a5fb;
20868	:douta	=	16'h	ae1b;
20869	:douta	=	16'h	9599;
20870	:douta	=	16'h	9dba;
20871	:douta	=	16'h	8d18;
20872	:douta	=	16'h	8d18;
20873	:douta	=	16'h	84f7;
20874	:douta	=	16'h	84d7;
20875	:douta	=	16'h	84f8;
20876	:douta	=	16'h	8d18;
20877	:douta	=	16'h	84d7;
20878	:douta	=	16'h	9559;
20879	:douta	=	16'h	8d39;
20880	:douta	=	16'h	84d7;
20881	:douta	=	16'h	8d18;
20882	:douta	=	16'h	84d7;
20883	:douta	=	16'h	8d38;
20884	:douta	=	16'h	84f7;
20885	:douta	=	16'h	84b7;
20886	:douta	=	16'h	84d7;
20887	:douta	=	16'h	84d7;
20888	:douta	=	16'h	8d39;
20889	:douta	=	16'h	9559;
20890	:douta	=	16'h	9d9a;
20891	:douta	=	16'h	9d9a;
20892	:douta	=	16'h	9579;
20893	:douta	=	16'h	9559;
20894	:douta	=	16'h	8d18;
20895	:douta	=	16'h	8d19;
20896	:douta	=	16'h	9559;
20897	:douta	=	16'h	8d39;
20898	:douta	=	16'h	8d39;
20899	:douta	=	16'h	8d59;
20900	:douta	=	16'h	9559;
20901	:douta	=	16'h	8d59;
20902	:douta	=	16'h	a5ba;
20903	:douta	=	16'h	9d99;
20904	:douta	=	16'h	8d19;
20905	:douta	=	16'h	838e;
20906	:douta	=	16'h	940e;
20907	:douta	=	16'h	6b0f;
20908	:douta	=	16'h	6cb8;
20909	:douta	=	16'h	1948;
20910	:douta	=	16'h	1906;
20911	:douta	=	16'h	0001;
20912	:douta	=	16'h	0043;
20913	:douta	=	16'h	42cf;
20914	:douta	=	16'h	9579;
20915	:douta	=	16'h	adfb;
20916	:douta	=	16'h	8c52;
20917	:douta	=	16'h	5aea;
20918	:douta	=	16'h	10c5;
20919	:douta	=	16'h	19ab;
20920	:douta	=	16'h	2ad2;
20921	:douta	=	16'h	54fb;
20922	:douta	=	16'h	54bb;
20923	:douta	=	16'h	4311;
20924	:douta	=	16'h	18e5;
20925	:douta	=	16'h	2082;
20926	:douta	=	16'h	49e8;
20927	:douta	=	16'h	4a09;
20928	:douta	=	16'h	4a8c;
20929	:douta	=	16'h	42d0;
20930	:douta	=	16'h	3189;
20931	:douta	=	16'h	1105;
20932	:douta	=	16'h	2148;
20933	:douta	=	16'h	857b;
20934	:douta	=	16'h	851a;
20935	:douta	=	16'h	7cd9;
20936	:douta	=	16'h	7cd9;
20937	:douta	=	16'h	7cf9;
20938	:douta	=	16'h	7cb9;
20939	:douta	=	16'h	8519;
20940	:douta	=	16'h	8d3a;
20941	:douta	=	16'h	957a;
20942	:douta	=	16'h	8d7a;
20943	:douta	=	16'h	9dbc;
20944	:douta	=	16'h	959c;
20945	:douta	=	16'h	8d5b;
20946	:douta	=	16'h	851a;
20947	:douta	=	16'h	84d9;
20948	:douta	=	16'h	6c77;
20949	:douta	=	16'h	853a;
20950	:douta	=	16'h	853a;
20951	:douta	=	16'h	8d7b;
20952	:douta	=	16'h	8d7b;
20953	:douta	=	16'h	8d5a;
20954	:douta	=	16'h	8d7b;
20955	:douta	=	16'h	8d19;
20956	:douta	=	16'h	7cd8;
20957	:douta	=	16'h	8d5a;
20958	:douta	=	16'h	7cf9;
20959	:douta	=	16'h	8d5a;
20960	:douta	=	16'h	95bb;
20961	:douta	=	16'h	7cf9;
20962	:douta	=	16'h	853a;
20963	:douta	=	16'h	853a;
20964	:douta	=	16'h	7cd9;
20965	:douta	=	16'h	851a;
20966	:douta	=	16'h	853a;
20967	:douta	=	16'h	7d1a;
20968	:douta	=	16'h	6457;
20969	:douta	=	16'h	6478;
20970	:douta	=	16'h	6457;
20971	:douta	=	16'h	6c57;
20972	:douta	=	16'h	6457;
20973	:douta	=	16'h	6cb9;
20974	:douta	=	16'h	7c13;
20975	:douta	=	16'h	6a46;
20976	:douta	=	16'h	324e;
20977	:douta	=	16'h	4372;
20978	:douta	=	16'h	9dbb;
20979	:douta	=	16'h	84b6;
20980	:douta	=	16'h	84f8;
20981	:douta	=	16'h	84b8;
20982	:douta	=	16'h	5bd4;
20983	:douta	=	16'h	5bf3;
20984	:douta	=	16'h	957a;
20985	:douta	=	16'h	4a28;
20986	:douta	=	16'h	7c55;
20987	:douta	=	16'h	9539;
20988	:douta	=	16'h	6c14;
20989	:douta	=	16'h	7c54;
20990	:douta	=	16'h	6bd2;
20991	:douta	=	16'h	638f;
20992	:douta	=	16'h	3146;
20993	:douta	=	16'h	0862;
20994	:douta	=	16'h	2126;
20995	:douta	=	16'h	3ad1;
20996	:douta	=	16'h	2a90;
20997	:douta	=	16'h	3b33;
20998	:douta	=	16'h	53f7;
20999	:douta	=	16'h	4374;
21000	:douta	=	16'h	32f1;
21001	:douta	=	16'h	4312;
21002	:douta	=	16'h	326f;
21003	:douta	=	16'h	7c98;
21004	:douta	=	16'h	6c57;
21005	:douta	=	16'h	957c;
21006	:douta	=	16'h	4acf;
21007	:douta	=	16'h	5b72;
21008	:douta	=	16'h	6bd3;
21009	:douta	=	16'h	73f3;
21010	:douta	=	16'h	9d37;
21011	:douta	=	16'h	8b8b;
21012	:douta	=	16'h	93aa;
21013	:douta	=	16'h	ac4c;
21014	:douta	=	16'h	ac6b;
21015	:douta	=	16'h	bc8b;
21016	:douta	=	16'h	d56f;
21017	:douta	=	16'h	cd6f;
21018	:douta	=	16'h	d5b0;
21019	:douta	=	16'h	ddd1;
21020	:douta	=	16'h	ee95;
21021	:douta	=	16'h	ee95;
21022	:douta	=	16'h	ee95;
21023	:douta	=	16'h	ee96;
21024	:douta	=	16'h	eeb6;
21025	:douta	=	16'h	ee74;
21026	:douta	=	16'h	e674;
21027	:douta	=	16'h	e654;
21028	:douta	=	16'h	cd70;
21029	:douta	=	16'h	c50f;
21030	:douta	=	16'h	c4cf;
21031	:douta	=	16'h	b48d;
21032	:douta	=	16'h	8b69;
21033	:douta	=	16'h	a42c;
21034	:douta	=	16'h	9bea;
21035	:douta	=	16'h	ac6c;
21036	:douta	=	16'h	b4ad;
21037	:douta	=	16'h	c52e;
21038	:douta	=	16'h	cd6f;
21039	:douta	=	16'h	d5b0;
21040	:douta	=	16'h	ddf3;
21041	:douta	=	16'h	e675;
21042	:douta	=	16'h	e655;
21043	:douta	=	16'h	e675;
21044	:douta	=	16'h	e675;
21045	:douta	=	16'h	eeb6;
21046	:douta	=	16'h	e674;
21047	:douta	=	16'h	e654;
21048	:douta	=	16'h	e654;
21049	:douta	=	16'h	e654;
21050	:douta	=	16'h	ddf2;
21051	:douta	=	16'h	dd92;
21052	:douta	=	16'h	cd70;
21053	:douta	=	16'h	bd0e;
21054	:douta	=	16'h	bcef;
21055	:douta	=	16'h	9c30;
21056	:douta	=	16'h	9451;
21057	:douta	=	16'h	8c11;
21058	:douta	=	16'h	7bd1;
21059	:douta	=	16'h	7bf2;
21060	:douta	=	16'h	734e;
21061	:douta	=	16'h	734e;
21062	:douta	=	16'h	7b8f;
21063	:douta	=	16'h	6b4f;
21064	:douta	=	16'h	630e;
21065	:douta	=	16'h	49a5;
21066	:douta	=	16'h	7b08;
21067	:douta	=	16'h	938a;
21068	:douta	=	16'h	a42c;
21069	:douta	=	16'h	93cc;
21070	:douta	=	16'h	d590;
21071	:douta	=	16'h	e634;
21072	:douta	=	16'h	e613;
21073	:douta	=	16'h	de12;
21074	:douta	=	16'h	dd8f;
21075	:douta	=	16'h	cd0e;
21076	:douta	=	16'h	a42d;
21077	:douta	=	16'h	ac2e;
21078	:douta	=	16'h	838e;
21079	:douta	=	16'h	732e;
21080	:douta	=	16'h	634e;
21081	:douta	=	16'h	632f;
21082	:douta	=	16'h	6350;
21083	:douta	=	16'h	4aef;
21084	:douta	=	16'h	5b51;
21085	:douta	=	16'h	4b10;
21086	:douta	=	16'h	42cf;
21087	:douta	=	16'h	324d;
21088	:douta	=	16'h	29ec;
21089	:douta	=	16'h	21a9;
21090	:douta	=	16'h	2168;
21091	:douta	=	16'h	0884;
21092	:douta	=	16'h	5b0e;
21093	:douta	=	16'h	0883;
21094	:douta	=	16'h	10c4;
21095	:douta	=	16'h	18e4;
21096	:douta	=	16'h	10e5;
21097	:douta	=	16'h	18c4;
21098	:douta	=	16'h	10c4;
21099	:douta	=	16'h	10c5;
21100	:douta	=	16'h	10a3;
21101	:douta	=	16'h	10a3;
21102	:douta	=	16'h	2146;
21103	:douta	=	16'h	10e4;
21104	:douta	=	16'h	18e5;
21105	:douta	=	16'h	3a0a;
21106	:douta	=	16'h	6bb1;
21107	:douta	=	16'h	2966;
21108	:douta	=	16'h	d678;
21109	:douta	=	16'h	9cb1;
21110	:douta	=	16'h	840e;
21111	:douta	=	16'h	2946;
21112	:douta	=	16'h	528a;
21113	:douta	=	16'h	5acb;
21114	:douta	=	16'h	0002;
21115	:douta	=	16'h	41c7;
21116	:douta	=	16'h	5b70;
21117	:douta	=	16'h	7c96;
21118	:douta	=	16'h	84f8;
21119	:douta	=	16'h	84f7;
21120	:douta	=	16'h	8d39;
21121	:douta	=	16'h	84f8;
21122	:douta	=	16'h	7c96;
21123	:douta	=	16'h	8d39;
21124	:douta	=	16'h	957a;
21125	:douta	=	16'h	a5fb;
21126	:douta	=	16'h	a5fb;
21127	:douta	=	16'h	9d7a;
21128	:douta	=	16'h	84d7;
21129	:douta	=	16'h	8d18;
21130	:douta	=	16'h	84f8;
21131	:douta	=	16'h	84f8;
21132	:douta	=	16'h	9559;
21133	:douta	=	16'h	84d7;
21134	:douta	=	16'h	84d7;
21135	:douta	=	16'h	84d7;
21136	:douta	=	16'h	7496;
21137	:douta	=	16'h	8d39;
21138	:douta	=	16'h	84f8;
21139	:douta	=	16'h	7c96;
21140	:douta	=	16'h	7cb6;
21141	:douta	=	16'h	84b6;
21142	:douta	=	16'h	84f8;
21143	:douta	=	16'h	7c96;
21144	:douta	=	16'h	84d7;
21145	:douta	=	16'h	84f7;
21146	:douta	=	16'h	84d7;
21147	:douta	=	16'h	9d9a;
21148	:douta	=	16'h	8d38;
21149	:douta	=	16'h	9579;
21150	:douta	=	16'h	9559;
21151	:douta	=	16'h	9559;
21152	:douta	=	16'h	8d39;
21153	:douta	=	16'h	9559;
21154	:douta	=	16'h	9579;
21155	:douta	=	16'h	9d9a;
21156	:douta	=	16'h	9d9a;
21157	:douta	=	16'h	84f8;
21158	:douta	=	16'h	84f8;
21159	:douta	=	16'h	9559;
21160	:douta	=	16'h	a5db;
21161	:douta	=	16'h	957a;
21162	:douta	=	16'h	7b4c;
21163	:douta	=	16'h	7b6e;
21164	:douta	=	16'h	7476;
21165	:douta	=	16'h	326f;
21166	:douta	=	16'h	322d;
21167	:douta	=	16'h	1906;
21168	:douta	=	16'h	18c4;
21169	:douta	=	16'h	0022;
21170	:douta	=	16'h	21eb;
21171	:douta	=	16'h	63d3;
21172	:douta	=	16'h	7bce;
21173	:douta	=	16'h	39a5;
21174	:douta	=	16'h	0882;
21175	:douta	=	16'h	1968;
21176	:douta	=	16'h	4c39;
21177	:douta	=	16'h	3312;
21178	:douta	=	16'h	2a2c;
21179	:douta	=	16'h	1082;
21180	:douta	=	16'h	3145;
21181	:douta	=	16'h	41e7;
21182	:douta	=	16'h	5a6a;
21183	:douta	=	16'h	49a7;
21184	:douta	=	16'h	6c98;
21185	:douta	=	16'h	31eb;
21186	:douta	=	16'h	29a9;
21187	:douta	=	16'h	324c;
21188	:douta	=	16'h	7cf9;
21189	:douta	=	16'h	7498;
21190	:douta	=	16'h	7cd8;
21191	:douta	=	16'h	84f9;
21192	:douta	=	16'h	7c98;
21193	:douta	=	16'h	84f9;
21194	:douta	=	16'h	7cd9;
21195	:douta	=	16'h	8d5a;
21196	:douta	=	16'h	957b;
21197	:douta	=	16'h	95bb;
21198	:douta	=	16'h	959b;
21199	:douta	=	16'h	9dbc;
21200	:douta	=	16'h	9dbc;
21201	:douta	=	16'h	9dbb;
21202	:douta	=	16'h	8d7a;
21203	:douta	=	16'h	9ddc;
21204	:douta	=	16'h	8d3a;
21205	:douta	=	16'h	7cd8;
21206	:douta	=	16'h	6436;
21207	:douta	=	16'h	7497;
21208	:douta	=	16'h	7cd8;
21209	:douta	=	16'h	851a;
21210	:douta	=	16'h	8d3a;
21211	:douta	=	16'h	957b;
21212	:douta	=	16'h	8d7b;
21213	:douta	=	16'h	853a;
21214	:douta	=	16'h	74b8;
21215	:douta	=	16'h	6415;
21216	:douta	=	16'h	6c56;
21217	:douta	=	16'h	959b;
21218	:douta	=	16'h	9ddc;
21219	:douta	=	16'h	8d5a;
21220	:douta	=	16'h	8d5b;
21221	:douta	=	16'h	7cf9;
21222	:douta	=	16'h	851a;
21223	:douta	=	16'h	74d9;
21224	:douta	=	16'h	853a;
21225	:douta	=	16'h	53d5;
21226	:douta	=	16'h	6437;
21227	:douta	=	16'h	5bd5;
21228	:douta	=	16'h	4b53;
21229	:douta	=	16'h	4bd6;
21230	:douta	=	16'h	7b8e;
21231	:douta	=	16'h	6b90;
21232	:douta	=	16'h	3880;
21233	:douta	=	16'h	1862;
21234	:douta	=	16'h	4b72;
21235	:douta	=	16'h	9559;
21236	:douta	=	16'h	adb9;
21237	:douta	=	16'h	8d39;
21238	:douta	=	16'h	53b4;
21239	:douta	=	16'h	7456;
21240	:douta	=	16'h	5350;
21241	:douta	=	16'h	28a1;
21242	:douta	=	16'h	9559;
21243	:douta	=	16'h	a599;
21244	:douta	=	16'h	9d98;
21245	:douta	=	16'h	9d78;
21246	:douta	=	16'h	1084;
21247	:douta	=	16'h	0000;
21248	:douta	=	16'h	2945;
21249	:douta	=	16'h	18e4;
21250	:douta	=	16'h	18e4;
21251	:douta	=	16'h	328f;
21252	:douta	=	16'h	3290;
21253	:douta	=	16'h	2a6f;
21254	:douta	=	16'h	4bb5;
21255	:douta	=	16'h	4374;
21256	:douta	=	16'h	2a2e;
21257	:douta	=	16'h	6415;
21258	:douta	=	16'h	5bf5;
21259	:douta	=	16'h	84d8;
21260	:douta	=	16'h	7456;
21261	:douta	=	16'h	7c77;
21262	:douta	=	16'h	5b72;
21263	:douta	=	16'h	5b51;
21264	:douta	=	16'h	7434;
21265	:douta	=	16'h	5b71;
21266	:douta	=	16'h	a599;
21267	:douta	=	16'h	9bca;
21268	:douta	=	16'h	ac4c;
21269	:douta	=	16'h	bccd;
21270	:douta	=	16'h	b4ad;
21271	:douta	=	16'h	c4ed;
21272	:douta	=	16'h	d5af;
21273	:douta	=	16'h	ddd1;
21274	:douta	=	16'h	e613;
21275	:douta	=	16'h	e633;
21276	:douta	=	16'h	eeb6;
21277	:douta	=	16'h	ee96;
21278	:douta	=	16'h	ee75;
21279	:douta	=	16'h	eeb6;
21280	:douta	=	16'h	e674;
21281	:douta	=	16'h	e654;
21282	:douta	=	16'h	d5b2;
21283	:douta	=	16'h	d5b1;
21284	:douta	=	16'h	cd70;
21285	:douta	=	16'h	bd0f;
21286	:douta	=	16'h	ac6c;
21287	:douta	=	16'h	8308;
21288	:douta	=	16'h	a40b;
21289	:douta	=	16'h	93ca;
21290	:douta	=	16'h	9beb;
21291	:douta	=	16'h	bccd;
21292	:douta	=	16'h	c50e;
21293	:douta	=	16'h	c52e;
21294	:douta	=	16'h	cd90;
21295	:douta	=	16'h	de12;
21296	:douta	=	16'h	e675;
21297	:douta	=	16'h	ee96;
21298	:douta	=	16'h	ee96;
21299	:douta	=	16'h	ee95;
21300	:douta	=	16'h	e675;
21301	:douta	=	16'h	eeb6;
21302	:douta	=	16'h	e674;
21303	:douta	=	16'h	e613;
21304	:douta	=	16'h	ddd2;
21305	:douta	=	16'h	ddd2;
21306	:douta	=	16'h	d591;
21307	:douta	=	16'h	c530;
21308	:douta	=	16'h	c510;
21309	:douta	=	16'h	b4af;
21310	:douta	=	16'h	9c50;
21311	:douta	=	16'h	9431;
21312	:douta	=	16'h	9431;
21313	:douta	=	16'h	8412;
21314	:douta	=	16'h	6aed;
21315	:douta	=	16'h	630e;
21316	:douta	=	16'h	736f;
21317	:douta	=	16'h	734e;
21318	:douta	=	16'h	6b0e;
21319	:douta	=	16'h	49e8;
21320	:douta	=	16'h	4185;
21321	:douta	=	16'h	a40b;
21322	:douta	=	16'h	9c0c;
21323	:douta	=	16'h	9bcb;
21324	:douta	=	16'h	c52f;
21325	:douta	=	16'h	cd6f;
21326	:douta	=	16'h	e5f2;
21327	:douta	=	16'h	e654;
21328	:douta	=	16'h	e654;
21329	:douta	=	16'h	e5f2;
21330	:douta	=	16'h	d58f;
21331	:douta	=	16'h	c4ee;
21332	:douta	=	16'h	a42d;
21333	:douta	=	16'h	a40d;
21334	:douta	=	16'h	838d;
21335	:douta	=	16'h	7b4d;
21336	:douta	=	16'h	632e;
21337	:douta	=	16'h	6b4f;
21338	:douta	=	16'h	634f;
21339	:douta	=	16'h	6b71;
21340	:douta	=	16'h	5b50;
21341	:douta	=	16'h	5331;
21342	:douta	=	16'h	52f0;
21343	:douta	=	16'h	3a8e;
21344	:douta	=	16'h	320c;
21345	:douta	=	16'h	29eb;
21346	:douta	=	16'h	2189;
21347	:douta	=	16'h	2168;
21348	:douta	=	16'h	0884;
21349	:douta	=	16'h	4ace;
21350	:douta	=	16'h	10a4;
21351	:douta	=	16'h	10e4;
21352	:douta	=	16'h	18c4;
21353	:douta	=	16'h	10c4;
21354	:douta	=	16'h	10c4;
21355	:douta	=	16'h	10a4;
21356	:douta	=	16'h	10c4;
21357	:douta	=	16'h	10c4;
21358	:douta	=	16'h	18e4;
21359	:douta	=	16'h	1905;
21360	:douta	=	16'h	1906;
21361	:douta	=	16'h	29a8;
21362	:douta	=	16'h	6b90;
21363	:douta	=	16'h	6b90;
21364	:douta	=	16'h	52ed;
21365	:douta	=	16'h	83ee;
21366	:douta	=	16'h	4228;
21367	:douta	=	16'h	5269;
21368	:douta	=	16'h	62cb;
21369	:douta	=	16'h	18e5;
21370	:douta	=	16'h	8c0f;
21371	:douta	=	16'h	6b2b;
21372	:douta	=	16'h	5269;
21373	:douta	=	16'h	6c13;
21374	:douta	=	16'h	84f8;
21375	:douta	=	16'h	8d38;
21376	:douta	=	16'h	7cb6;
21377	:douta	=	16'h	84d7;
21378	:douta	=	16'h	8d18;
21379	:douta	=	16'h	84b7;
21380	:douta	=	16'h	8d59;
21381	:douta	=	16'h	9579;
21382	:douta	=	16'h	84f8;
21383	:douta	=	16'h	8d39;
21384	:douta	=	16'h	9579;
21385	:douta	=	16'h	a5da;
21386	:douta	=	16'h	a5ba;
21387	:douta	=	16'h	9558;
21388	:douta	=	16'h	7476;
21389	:douta	=	16'h	7cb7;
21390	:douta	=	16'h	8d18;
21391	:douta	=	16'h	7496;
21392	:douta	=	16'h	7cb7;
21393	:douta	=	16'h	84f7;
21394	:douta	=	16'h	7c96;
21395	:douta	=	16'h	84d7;
21396	:douta	=	16'h	8d38;
21397	:douta	=	16'h	8d18;
21398	:douta	=	16'h	9579;
21399	:douta	=	16'h	8d39;
21400	:douta	=	16'h	84f8;
21401	:douta	=	16'h	84d7;
21402	:douta	=	16'h	84f7;
21403	:douta	=	16'h	8d18;
21404	:douta	=	16'h	9559;
21405	:douta	=	16'h	8d39;
21406	:douta	=	16'h	84f8;
21407	:douta	=	16'h	8d18;
21408	:douta	=	16'h	9559;
21409	:douta	=	16'h	957a;
21410	:douta	=	16'h	9559;
21411	:douta	=	16'h	84f8;
21412	:douta	=	16'h	8d18;
21413	:douta	=	16'h	7cd7;
21414	:douta	=	16'h	a5db;
21415	:douta	=	16'h	9559;
21416	:douta	=	16'h	7496;
21417	:douta	=	16'h	7cd7;
21418	:douta	=	16'h	a5fc;
21419	:douta	=	16'h	9db9;
21420	:douta	=	16'h	6330;
21421	:douta	=	16'h	6bd3;
21422	:douta	=	16'h	4a8d;
21423	:douta	=	16'h	1989;
21424	:douta	=	16'h	1968;
21425	:douta	=	16'h	21aa;
21426	:douta	=	16'h	1948;
21427	:douta	=	16'h	10e5;
21428	:douta	=	16'h	0064;
21429	:douta	=	16'h	10c5;
21430	:douta	=	16'h	2146;
21431	:douta	=	16'h	1905;
21432	:douta	=	16'h	1061;
21433	:douta	=	16'h	3186;
21434	:douta	=	16'h	4a08;
21435	:douta	=	16'h	834c;
21436	:douta	=	16'h	8b4b;
21437	:douta	=	16'h	832b;
21438	:douta	=	16'h	6c14;
21439	:douta	=	16'h	63f4;
21440	:douta	=	16'h	5350;
21441	:douta	=	16'h	4a8d;
21442	:douta	=	16'h	7c97;
21443	:douta	=	16'h	853b;
21444	:douta	=	16'h	8519;
21445	:douta	=	16'h	7cb8;
21446	:douta	=	16'h	6c78;
21447	:douta	=	16'h	6c37;
21448	:douta	=	16'h	959c;
21449	:douta	=	16'h	959b;
21450	:douta	=	16'h	74b8;
21451	:douta	=	16'h	7cb8;
21452	:douta	=	16'h	7c98;
21453	:douta	=	16'h	7cb8;
21454	:douta	=	16'h	8d3a;
21455	:douta	=	16'h	8d5a;
21456	:douta	=	16'h	a61c;
21457	:douta	=	16'h	a5fc;
21458	:douta	=	16'h	851a;
21459	:douta	=	16'h	8d5b;
21460	:douta	=	16'h	95bb;
21461	:douta	=	16'h	8d5b;
21462	:douta	=	16'h	95dc;
21463	:douta	=	16'h	95bc;
21464	:douta	=	16'h	95bc;
21465	:douta	=	16'h	84d9;
21466	:douta	=	16'h	7d19;
21467	:douta	=	16'h	74b8;
21468	:douta	=	16'h	7477;
21469	:douta	=	16'h	74b8;
21470	:douta	=	16'h	959c;
21471	:douta	=	16'h	8d7b;
21472	:douta	=	16'h	95bb;
21473	:douta	=	16'h	851a;
21474	:douta	=	16'h	6c16;
21475	:douta	=	16'h	5bf5;
21476	:douta	=	16'h	74b8;
21477	:douta	=	16'h	853a;
21478	:douta	=	16'h	7cf9;
21479	:douta	=	16'h	851a;
21480	:douta	=	16'h	7cd9;
21481	:douta	=	16'h	74d9;
21482	:douta	=	16'h	7d1a;
21483	:douta	=	16'h	857b;
21484	:douta	=	16'h	857c;
21485	:douta	=	16'h	73b1;
21486	:douta	=	16'h	7c98;
21487	:douta	=	16'h	63d4;
21488	:douta	=	16'h	4374;
21489	:douta	=	16'h	63d3;
21490	:douta	=	16'h	72a6;
21491	:douta	=	16'h	3965;
21492	:douta	=	16'h	2a4d;
21493	:douta	=	16'h	7d3b;
21494	:douta	=	16'h	7499;
21495	:douta	=	16'h	6c56;
21496	:douta	=	16'h	4165;
21497	:douta	=	16'h	2924;
21498	:douta	=	16'h	a5db;
21499	:douta	=	16'h	84b6;
21500	:douta	=	16'h	63d5;
21501	:douta	=	16'h	3a4c;
21502	:douta	=	16'h	2125;
21503	:douta	=	16'h	1083;
21504	:douta	=	16'h	3166;
21505	:douta	=	16'h	18e4;
21506	:douta	=	16'h	1083;
21507	:douta	=	16'h	328e;
21508	:douta	=	16'h	4b94;
21509	:douta	=	16'h	32b0;
21510	:douta	=	16'h	4353;
21511	:douta	=	16'h	3af2;
21512	:douta	=	16'h	4353;
21513	:douta	=	16'h	6c36;
21514	:douta	=	16'h	5bf5;
21515	:douta	=	16'h	84d8;
21516	:douta	=	16'h	7457;
21517	:douta	=	16'h	7cb8;
21518	:douta	=	16'h	5b52;
21519	:douta	=	16'h	6bb3;
21520	:douta	=	16'h	84b6;
21521	:douta	=	16'h	8cb6;
21522	:douta	=	16'h	73f3;
21523	:douta	=	16'h	ac4b;
21524	:douta	=	16'h	b4ac;
21525	:douta	=	16'h	bccd;
21526	:douta	=	16'h	bcad;
21527	:douta	=	16'h	c50e;
21528	:douta	=	16'h	d5d0;
21529	:douta	=	16'h	ddf2;
21530	:douta	=	16'h	e634;
21531	:douta	=	16'h	e654;
21532	:douta	=	16'h	ee96;
21533	:douta	=	16'h	eeb6;
21534	:douta	=	16'h	e675;
21535	:douta	=	16'h	e633;
21536	:douta	=	16'h	ee95;
21537	:douta	=	16'h	ddf2;
21538	:douta	=	16'h	d591;
21539	:douta	=	16'h	d590;
21540	:douta	=	16'h	cd4f;
21541	:douta	=	16'h	bcee;
21542	:douta	=	16'h	93aa;
21543	:douta	=	16'h	9bcb;
21544	:douta	=	16'h	ac6c;
21545	:douta	=	16'h	9c0b;
21546	:douta	=	16'h	a44c;
21547	:douta	=	16'h	bcee;
21548	:douta	=	16'h	c50e;
21549	:douta	=	16'h	cd6f;
21550	:douta	=	16'h	d5b1;
21551	:douta	=	16'h	de13;
21552	:douta	=	16'h	e675;
21553	:douta	=	16'h	ee96;
21554	:douta	=	16'h	ee96;
21555	:douta	=	16'h	ee75;
21556	:douta	=	16'h	ee75;
21557	:douta	=	16'h	ee75;
21558	:douta	=	16'h	ee75;
21559	:douta	=	16'h	e632;
21560	:douta	=	16'h	ddb2;
21561	:douta	=	16'h	d590;
21562	:douta	=	16'h	cd71;
21563	:douta	=	16'h	c4f0;
21564	:douta	=	16'h	bcd0;
21565	:douta	=	16'h	ac8f;
21566	:douta	=	16'h	9c50;
21567	:douta	=	16'h	8c11;
21568	:douta	=	16'h	83f1;
21569	:douta	=	16'h	7b90;
21570	:douta	=	16'h	62cd;
21571	:douta	=	16'h	62cd;
21572	:douta	=	16'h	5acc;
21573	:douta	=	16'h	5aee;
21574	:douta	=	16'h	5aab;
21575	:douta	=	16'h	4164;
21576	:douta	=	16'h	7ac7;
21577	:douta	=	16'h	ac2c;
21578	:douta	=	16'h	b48e;
21579	:douta	=	16'h	bcae;
21580	:douta	=	16'h	d5b1;
21581	:douta	=	16'h	ddf2;
21582	:douta	=	16'h	e634;
21583	:douta	=	16'h	ee55;
21584	:douta	=	16'h	e633;
21585	:douta	=	16'h	ddd1;
21586	:douta	=	16'h	d58f;
21587	:douta	=	16'h	bcad;
21588	:douta	=	16'h	a42d;
21589	:douta	=	16'h	9bed;
21590	:douta	=	16'h	a42e;
21591	:douta	=	16'h	838d;
21592	:douta	=	16'h	734f;
21593	:douta	=	16'h	6b4f;
21594	:douta	=	16'h	634f;
21595	:douta	=	16'h	6b71;
21596	:douta	=	16'h	6371;
21597	:douta	=	16'h	5b72;
21598	:douta	=	16'h	4af0;
21599	:douta	=	16'h	42ae;
21600	:douta	=	16'h	322c;
21601	:douta	=	16'h	2a0c;
21602	:douta	=	16'h	29ea;
21603	:douta	=	16'h	21a9;
21604	:douta	=	16'h	2128;
21605	:douta	=	16'h	428d;
21606	:douta	=	16'h	4a8d;
21607	:douta	=	16'h	10a3;
21608	:douta	=	16'h	10e5;
21609	:douta	=	16'h	10c4;
21610	:douta	=	16'h	10a3;
21611	:douta	=	16'h	18e4;
21612	:douta	=	16'h	10a4;
21613	:douta	=	16'h	10e4;
21614	:douta	=	16'h	10a3;
21615	:douta	=	16'h	10c5;
21616	:douta	=	16'h	18e5;
21617	:douta	=	16'h	0042;
21618	:douta	=	16'h	18e5;
21619	:douta	=	16'h	7433;
21620	:douta	=	16'h	5b50;
21621	:douta	=	16'h	9cd2;
21622	:douta	=	16'h	6b2c;
21623	:douta	=	16'h	8bce;
21624	:douta	=	16'h	8bcd;
21625	:douta	=	16'h	41e8;
21626	:douta	=	16'h	8c30;
21627	:douta	=	16'h	734d;
21628	:douta	=	16'h	a4f1;
21629	:douta	=	16'h	2968;
21630	:douta	=	16'h	8d7a;
21631	:douta	=	16'h	7cb6;
21632	:douta	=	16'h	7c96;
21633	:douta	=	16'h	7c96;
21634	:douta	=	16'h	7475;
21635	:douta	=	16'h	84d7;
21636	:douta	=	16'h	6c14;
21637	:douta	=	16'h	84d7;
21638	:douta	=	16'h	8d38;
21639	:douta	=	16'h	8cf8;
21640	:douta	=	16'h	7c96;
21641	:douta	=	16'h	8d38;
21642	:douta	=	16'h	9d9a;
21643	:douta	=	16'h	a5db;
21644	:douta	=	16'h	a599;
21645	:douta	=	16'h	8d39;
21646	:douta	=	16'h	84f8;
21647	:douta	=	16'h	84f8;
21648	:douta	=	16'h	7c97;
21649	:douta	=	16'h	84b6;
21650	:douta	=	16'h	8d38;
21651	:douta	=	16'h	84f8;
21652	:douta	=	16'h	84b7;
21653	:douta	=	16'h	84b7;
21654	:douta	=	16'h	8d17;
21655	:douta	=	16'h	8d18;
21656	:douta	=	16'h	8d18;
21657	:douta	=	16'h	9539;
21658	:douta	=	16'h	8cd8;
21659	:douta	=	16'h	84d7;
21660	:douta	=	16'h	8d39;
21661	:douta	=	16'h	a5ba;
21662	:douta	=	16'h	9559;
21663	:douta	=	16'h	8d18;
21664	:douta	=	16'h	8d18;
21665	:douta	=	16'h	957a;
21666	:douta	=	16'h	9dba;
21667	:douta	=	16'h	9559;
21668	:douta	=	16'h	8d59;
21669	:douta	=	16'h	7cb7;
21670	:douta	=	16'h	8d18;
21671	:douta	=	16'h	959a;
21672	:douta	=	16'h	957a;
21673	:douta	=	16'h	9559;
21674	:douta	=	16'h	7c97;
21675	:douta	=	16'h	957b;
21676	:douta	=	16'h	8495;
21677	:douta	=	16'h	630e;
21678	:douta	=	16'h	424b;
21679	:douta	=	16'h	4aae;
21680	:douta	=	16'h	3a6d;
21681	:douta	=	16'h	1127;
21682	:douta	=	16'h	21a9;
21683	:douta	=	16'h	21a9;
21684	:douta	=	16'h	1947;
21685	:douta	=	16'h	10c5;
21686	:douta	=	16'h	0882;
21687	:douta	=	16'h	2125;
21688	:douta	=	16'h	49e8;
21689	:douta	=	16'h	8b6b;
21690	:douta	=	16'h	a40e;
21691	:douta	=	16'h	936c;
21692	:douta	=	16'h	7bf2;
21693	:douta	=	16'h	7476;
21694	:douta	=	16'h	5350;
21695	:douta	=	16'h	3a0a;
21696	:douta	=	16'h	4a8d;
21697	:douta	=	16'h	95bc;
21698	:douta	=	16'h	a61d;
21699	:douta	=	16'h	8d19;
21700	:douta	=	16'h	8d3a;
21701	:douta	=	16'h	9dbb;
21702	:douta	=	16'h	9539;
21703	:douta	=	16'h	7c77;
21704	:douta	=	16'h	5394;
21705	:douta	=	16'h	7498;
21706	:douta	=	16'h	957b;
21707	:douta	=	16'h	7cb8;
21708	:douta	=	16'h	74b8;
21709	:douta	=	16'h	7c97;
21710	:douta	=	16'h	7c98;
21711	:douta	=	16'h	851a;
21712	:douta	=	16'h	8d5b;
21713	:douta	=	16'h	9dbb;
21714	:douta	=	16'h	a63d;
21715	:douta	=	16'h	8d7a;
21716	:douta	=	16'h	8d5a;
21717	:douta	=	16'h	84f9;
21718	:douta	=	16'h	8d5b;
21719	:douta	=	16'h	851a;
21720	:douta	=	16'h	8d9b;
21721	:douta	=	16'h	9ddc;
21722	:douta	=	16'h	853a;
21723	:douta	=	16'h	7c98;
21724	:douta	=	16'h	7cd8;
21725	:douta	=	16'h	74b7;
21726	:douta	=	16'h	6415;
21727	:douta	=	16'h	95bc;
21728	:douta	=	16'h	853a;
21729	:douta	=	16'h	95dc;
21730	:douta	=	16'h	95bc;
21731	:douta	=	16'h	6c57;
21732	:douta	=	16'h	6c77;
21733	:douta	=	16'h	6416;
21734	:douta	=	16'h	7cd9;
21735	:douta	=	16'h	74b8;
21736	:douta	=	16'h	6c77;
21737	:douta	=	16'h	7cf9;
21738	:douta	=	16'h	74b8;
21739	:douta	=	16'h	751b;
21740	:douta	=	16'h	7d3a;
21741	:douta	=	16'h	52ce;
21742	:douta	=	16'h	63f5;
21743	:douta	=	16'h	9d9a;
21744	:douta	=	16'h	63f4;
21745	:douta	=	16'h	7cb8;
21746	:douta	=	16'h	959a;
21747	:douta	=	16'h	6249;
21748	:douta	=	16'h	40e1;
21749	:douta	=	16'h	29aa;
21750	:douta	=	16'h	53b5;
21751	:douta	=	16'h	7d5c;
21752	:douta	=	16'h	1000;
21753	:douta	=	16'h	42ce;
21754	:douta	=	16'h	9559;
21755	:douta	=	16'h	be7b;
21756	:douta	=	16'h	7455;
21757	:douta	=	16'h	6414;
21758	:douta	=	16'h	2967;
21759	:douta	=	16'h	1083;
21760	:douta	=	16'h	39a7;
21761	:douta	=	16'h	2104;
21762	:douta	=	16'h	1083;
21763	:douta	=	16'h	29ca;
21764	:douta	=	16'h	3b33;
21765	:douta	=	16'h	32b0;
21766	:douta	=	16'h	4b95;
21767	:douta	=	16'h	4374;
21768	:douta	=	16'h	222e;
21769	:douta	=	16'h	53b4;
21770	:douta	=	16'h	4b73;
21771	:douta	=	16'h	5351;
21772	:douta	=	16'h	5bb3;
21773	:douta	=	16'h	5bb4;
21774	:douta	=	16'h	5351;
21775	:douta	=	16'h	6bb2;
21776	:douta	=	16'h	8cd7;
21777	:douta	=	16'h	7c55;
21778	:douta	=	16'h	94d5;
21779	:douta	=	16'h	bcad;
21780	:douta	=	16'h	b4cd;
21781	:douta	=	16'h	c50e;
21782	:douta	=	16'h	c52e;
21783	:douta	=	16'h	cd4f;
21784	:douta	=	16'h	ddf2;
21785	:douta	=	16'h	e634;
21786	:douta	=	16'h	e675;
21787	:douta	=	16'h	ee95;
21788	:douta	=	16'h	ee95;
21789	:douta	=	16'h	ee75;
21790	:douta	=	16'h	e654;
21791	:douta	=	16'h	ddf1;
21792	:douta	=	16'h	cd2f;
21793	:douta	=	16'h	e633;
21794	:douta	=	16'h	c50e;
21795	:douta	=	16'h	c4ee;
21796	:douta	=	16'h	b4cd;
21797	:douta	=	16'h	a40b;
21798	:douta	=	16'h	8b69;
21799	:douta	=	16'h	ac6d;
21800	:douta	=	16'h	b4ad;
21801	:douta	=	16'h	ac4c;
21802	:douta	=	16'h	a42b;
21803	:douta	=	16'h	bcee;
21804	:douta	=	16'h	d590;
21805	:douta	=	16'h	ddd1;
21806	:douta	=	16'h	de13;
21807	:douta	=	16'h	e654;
21808	:douta	=	16'h	ee96;
21809	:douta	=	16'h	ee96;
21810	:douta	=	16'h	ee96;
21811	:douta	=	16'h	ee95;
21812	:douta	=	16'h	ee95;
21813	:douta	=	16'h	e654;
21814	:douta	=	16'h	e654;
21815	:douta	=	16'h	e654;
21816	:douta	=	16'h	d591;
21817	:douta	=	16'h	cd50;
21818	:douta	=	16'h	bcce;
21819	:douta	=	16'h	ac8f;
21820	:douta	=	16'h	9430;
21821	:douta	=	16'h	8c10;
21822	:douta	=	16'h	9430;
21823	:douta	=	16'h	8bf1;
21824	:douta	=	16'h	734f;
21825	:douta	=	16'h	6b2e;
21826	:douta	=	16'h	6b0d;
21827	:douta	=	16'h	6b0d;
21828	:douta	=	16'h	5a6b;
21829	:douta	=	16'h	2904;
21830	:douta	=	16'h	4963;
21831	:douta	=	16'h	93ca;
21832	:douta	=	16'h	9bcb;
21833	:douta	=	16'h	a46c;
21834	:douta	=	16'h	cd2f;
21835	:douta	=	16'h	d5b1;
21836	:douta	=	16'h	e654;
21837	:douta	=	16'h	ee75;
21838	:douta	=	16'h	ee75;
21839	:douta	=	16'h	e655;
21840	:douta	=	16'h	de12;
21841	:douta	=	16'h	dd90;
21842	:douta	=	16'h	d56f;
21843	:douta	=	16'h	c4cd;
21844	:douta	=	16'h	a40d;
21845	:douta	=	16'h	a40d;
21846	:douta	=	16'h	9bed;
21847	:douta	=	16'h	9bef;
21848	:douta	=	16'h	83af;
21849	:douta	=	16'h	8bd0;
21850	:douta	=	16'h	7390;
21851	:douta	=	16'h	6370;
21852	:douta	=	16'h	6bb1;
21853	:douta	=	16'h	6371;
21854	:douta	=	16'h	5b51;
21855	:douta	=	16'h	42cf;
21856	:douta	=	16'h	42ae;
21857	:douta	=	16'h	428e;
21858	:douta	=	16'h	2a2c;
21859	:douta	=	16'h	322c;
21860	:douta	=	16'h	2a0b;
21861	:douta	=	16'h	29ea;
21862	:douta	=	16'h	1927;
21863	:douta	=	16'h	530e;
21864	:douta	=	16'h	2127;
21865	:douta	=	16'h	18c4;
21866	:douta	=	16'h	10c4;
21867	:douta	=	16'h	10a4;
21868	:douta	=	16'h	10a3;
21869	:douta	=	16'h	08a3;
21870	:douta	=	16'h	10e4;
21871	:douta	=	16'h	10c4;
21872	:douta	=	16'h	10a3;
21873	:douta	=	16'h	10e4;
21874	:douta	=	16'h	18e4;
21875	:douta	=	16'h	0021;
21876	:douta	=	16'h	7411;
21877	:douta	=	16'h	6bf1;
21878	:douta	=	16'h	7bd0;
21879	:douta	=	16'h	ad33;
21880	:douta	=	16'h	94b1;
21881	:douta	=	16'h	a4b0;
21882	:douta	=	16'h	ad12;
21883	:douta	=	16'h	ad31;
21884	:douta	=	16'h	632b;
21885	:douta	=	16'h	62aa;
21886	:douta	=	16'h	20e6;
21887	:douta	=	16'h	7cb7;
21888	:douta	=	16'h	7455;
21889	:douta	=	16'h	7455;
21890	:douta	=	16'h	8cf8;
21891	:douta	=	16'h	84d7;
21892	:douta	=	16'h	8d39;
21893	:douta	=	16'h	8d18;
21894	:douta	=	16'h	84f8;
21895	:douta	=	16'h	84b7;
21896	:douta	=	16'h	8518;
21897	:douta	=	16'h	84f7;
21898	:douta	=	16'h	7476;
21899	:douta	=	16'h	7cb7;
21900	:douta	=	16'h	7cd7;
21901	:douta	=	16'h	84f7;
21902	:douta	=	16'h	84f7;
21903	:douta	=	16'h	84b6;
21904	:douta	=	16'h	9517;
21905	:douta	=	16'h	9dba;
21906	:douta	=	16'h	9559;
21907	:douta	=	16'h	84b6;
21908	:douta	=	16'h	8d18;
21909	:douta	=	16'h	957a;
21910	:douta	=	16'h	8d18;
21911	:douta	=	16'h	9d79;
21912	:douta	=	16'h	9579;
21913	:douta	=	16'h	959a;
21914	:douta	=	16'h	9dba;
21915	:douta	=	16'h	9d79;
21916	:douta	=	16'h	8518;
21917	:douta	=	16'h	84b6;
21918	:douta	=	16'h	84f8;
21919	:douta	=	16'h	84d7;
21920	:douta	=	16'h	9559;
21921	:douta	=	16'h	a5bb;
21922	:douta	=	16'h	9d9a;
21923	:douta	=	16'h	8d18;
21924	:douta	=	16'h	84d8;
21925	:douta	=	16'h	8518;
21926	:douta	=	16'h	9d9a;
21927	:douta	=	16'h	8d19;
21928	:douta	=	16'h	8d39;
21929	:douta	=	16'h	8518;
21930	:douta	=	16'h	9559;
21931	:douta	=	16'h	955a;
21932	:douta	=	16'h	957a;
21933	:douta	=	16'h	8519;
21934	:douta	=	16'h	8d18;
21935	:douta	=	16'h	634f;
21936	:douta	=	16'h	5a8c;
21937	:douta	=	16'h	52ee;
21938	:douta	=	16'h	5bb3;
21939	:douta	=	16'h	4b51;
21940	:douta	=	16'h	324d;
21941	:douta	=	16'h	1927;
21942	:douta	=	16'h	1968;
21943	:douta	=	16'h	5acd;
21944	:douta	=	16'h	ac8f;
21945	:douta	=	16'h	6b71;
21946	:douta	=	16'h	63b2;
21947	:douta	=	16'h	4a6e;
21948	:douta	=	16'h	4a4b;
21949	:douta	=	16'h	5ace;
21950	:douta	=	16'h	957b;
21951	:douta	=	16'h	a63d;
21952	:douta	=	16'h	9d9b;
21953	:douta	=	16'h	9559;
21954	:douta	=	16'h	8d3a;
21955	:douta	=	16'h	9ddb;
21956	:douta	=	16'h	9dba;
21957	:douta	=	16'h	9ddb;
21958	:douta	=	16'h	8d7a;
21959	:douta	=	16'h	8d5a;
21960	:douta	=	16'h	ae3d;
21961	:douta	=	16'h	ae1c;
21962	:douta	=	16'h	74b7;
21963	:douta	=	16'h	7cb8;
21964	:douta	=	16'h	6c36;
21965	:douta	=	16'h	7cd8;
21966	:douta	=	16'h	853a;
21967	:douta	=	16'h	8519;
21968	:douta	=	16'h	8d5a;
21969	:douta	=	16'h	8d7a;
21970	:douta	=	16'h	6c56;
21971	:douta	=	16'h	7cd8;
21972	:douta	=	16'h	8d5a;
21973	:douta	=	16'h	7cb9;
21974	:douta	=	16'h	853a;
21975	:douta	=	16'h	8d9b;
21976	:douta	=	16'h	a61d;
21977	:douta	=	16'h	9d9b;
21978	:douta	=	16'h	95bb;
21979	:douta	=	16'h	959a;
21980	:douta	=	16'h	a5fc;
21981	:douta	=	16'h	959b;
21982	:douta	=	16'h	95bc;
21983	:douta	=	16'h	7498;
21984	:douta	=	16'h	74b8;
21985	:douta	=	16'h	7498;
21986	:douta	=	16'h	7457;
21987	:douta	=	16'h	853a;
21988	:douta	=	16'h	7d3a;
21989	:douta	=	16'h	7cf9;
21990	:douta	=	16'h	7cd9;
21991	:douta	=	16'h	7d19;
21992	:douta	=	16'h	8d9c;
21993	:douta	=	16'h	6477;
21994	:douta	=	16'h	5c18;
21995	:douta	=	16'h	6aec;
21996	:douta	=	16'h	530f;
21997	:douta	=	16'h	5bb3;
21998	:douta	=	16'h	8d39;
21999	:douta	=	16'h	63f5;
22000	:douta	=	16'h	7cb7;
22001	:douta	=	16'h	84f9;
22002	:douta	=	16'h	4b73;
22003	:douta	=	16'h	9559;
22004	:douta	=	16'h	8d7a;
22005	:douta	=	16'h	9517;
22006	:douta	=	16'h	840e;
22007	:douta	=	16'h	5164;
22008	:douta	=	16'h	0883;
22009	:douta	=	16'h	3b30;
22010	:douta	=	16'h	adfc;
22011	:douta	=	16'h	84d7;
22012	:douta	=	16'h	6c35;
22013	:douta	=	16'h	7cb7;
22014	:douta	=	16'h	632e;
22015	:douta	=	16'h	10a3;
22016	:douta	=	16'h	39a7;
22017	:douta	=	16'h	2925;
22018	:douta	=	16'h	18a4;
22019	:douta	=	16'h	322b;
22020	:douta	=	16'h	3b12;
22021	:douta	=	16'h	3290;
22022	:douta	=	16'h	3b13;
22023	:douta	=	16'h	53f6;
22024	:douta	=	16'h	2a4f;
22025	:douta	=	16'h	5bd5;
22026	:douta	=	16'h	6c36;
22027	:douta	=	16'h	7cb7;
22028	:douta	=	16'h	7476;
22029	:douta	=	16'h	6c15;
22030	:douta	=	16'h	5b52;
22031	:douta	=	16'h	6b92;
22032	:douta	=	16'h	84b6;
22033	:douta	=	16'h	63d2;
22034	:douta	=	16'h	7bf2;
22035	:douta	=	16'h	bcad;
22036	:douta	=	16'h	bced;
22037	:douta	=	16'h	c50e;
22038	:douta	=	16'h	cd4f;
22039	:douta	=	16'h	d590;
22040	:douta	=	16'h	de13;
22041	:douta	=	16'h	e654;
22042	:douta	=	16'h	ee75;
22043	:douta	=	16'h	e654;
22044	:douta	=	16'h	ee95;
22045	:douta	=	16'h	e674;
22046	:douta	=	16'h	e653;
22047	:douta	=	16'h	ddf2;
22048	:douta	=	16'h	c50d;
22049	:douta	=	16'h	c50f;
22050	:douta	=	16'h	d590;
22051	:douta	=	16'h	c4ee;
22052	:douta	=	16'h	9bea;
22053	:douta	=	16'h	72c6;
22054	:douta	=	16'h	ac4c;
22055	:douta	=	16'h	ac6d;
22056	:douta	=	16'h	b4ad;
22057	:douta	=	16'h	ac6d;
22058	:douta	=	16'h	ac6c;
22059	:douta	=	16'h	cd8f;
22060	:douta	=	16'h	cd90;
22061	:douta	=	16'h	ddf2;
22062	:douta	=	16'h	de33;
22063	:douta	=	16'h	ee75;
22064	:douta	=	16'h	e695;
22065	:douta	=	16'h	eeb7;
22066	:douta	=	16'h	ee96;
22067	:douta	=	16'h	ee95;
22068	:douta	=	16'h	e675;
22069	:douta	=	16'h	e654;
22070	:douta	=	16'h	e613;
22071	:douta	=	16'h	de33;
22072	:douta	=	16'h	d5d2;
22073	:douta	=	16'h	cd4f;
22074	:douta	=	16'h	a46f;
22075	:douta	=	16'h	a450;
22076	:douta	=	16'h	9c50;
22077	:douta	=	16'h	7bb0;
22078	:douta	=	16'h	83d0;
22079	:douta	=	16'h	83f0;
22080	:douta	=	16'h	6b0d;
22081	:douta	=	16'h	62ec;
22082	:douta	=	16'h	630c;
22083	:douta	=	16'h	630c;
22084	:douta	=	16'h	41e8;
22085	:douta	=	16'h	51a4;
22086	:douta	=	16'h	8b48;
22087	:douta	=	16'h	9c0b;
22088	:douta	=	16'h	9c0c;
22089	:douta	=	16'h	bccd;
22090	:douta	=	16'h	d5b1;
22091	:douta	=	16'h	de13;
22092	:douta	=	16'h	ee95;
22093	:douta	=	16'h	ee95;
22094	:douta	=	16'h	ee75;
22095	:douta	=	16'h	de13;
22096	:douta	=	16'h	ddd1;
22097	:douta	=	16'h	d54f;
22098	:douta	=	16'h	cd0e;
22099	:douta	=	16'h	c4cd;
22100	:douta	=	16'h	a42d;
22101	:douta	=	16'h	ac2d;
22102	:douta	=	16'h	9c0e;
22103	:douta	=	16'h	93ce;
22104	:douta	=	16'h	8bcf;
22105	:douta	=	16'h	8bd0;
22106	:douta	=	16'h	7bb0;
22107	:douta	=	16'h	6b91;
22108	:douta	=	16'h	6bb1;
22109	:douta	=	16'h	6bb2;
22110	:douta	=	16'h	6392;
22111	:douta	=	16'h	4b10;
22112	:douta	=	16'h	42ae;
22113	:douta	=	16'h	428e;
22114	:douta	=	16'h	322c;
22115	:douta	=	16'h	324d;
22116	:douta	=	16'h	2a0b;
22117	:douta	=	16'h	322b;
22118	:douta	=	16'h	2189;
22119	:douta	=	16'h	3a4b;
22120	:douta	=	16'h	5b0f;
22121	:douta	=	16'h	0862;
22122	:douta	=	16'h	18e4;
22123	:douta	=	16'h	10c4;
22124	:douta	=	16'h	10a3;
22125	:douta	=	16'h	10a3;
22126	:douta	=	16'h	10c4;
22127	:douta	=	16'h	10c5;
22128	:douta	=	16'h	18e5;
22129	:douta	=	16'h	1905;
22130	:douta	=	16'h	1926;
22131	:douta	=	16'h	18e5;
22132	:douta	=	16'h	2988;
22133	:douta	=	16'h	6b90;
22134	:douta	=	16'h	5b50;
22135	:douta	=	16'h	4b2f;
22136	:douta	=	16'h	0842;
22137	:douta	=	16'h	a4b1;
22138	:douta	=	16'h	9cb0;
22139	:douta	=	16'h	83ee;
22140	:douta	=	16'h	5aaa;
22141	:douta	=	16'h	c5f4;
22142	:douta	=	16'h	7b8c;
22143	:douta	=	16'h	31ea;
22144	:douta	=	16'h	9559;
22145	:douta	=	16'h	84d6;
22146	:douta	=	16'h	6c34;
22147	:douta	=	16'h	7c96;
22148	:douta	=	16'h	7cb7;
22149	:douta	=	16'h	84d7;
22150	:douta	=	16'h	9559;
22151	:douta	=	16'h	84f8;
22152	:douta	=	16'h	84f8;
22153	:douta	=	16'h	8d18;
22154	:douta	=	16'h	84f8;
22155	:douta	=	16'h	84d7;
22156	:douta	=	16'h	84d7;
22157	:douta	=	16'h	8518;
22158	:douta	=	16'h	9559;
22159	:douta	=	16'h	6c14;
22160	:douta	=	16'h	6c14;
22161	:douta	=	16'h	84d6;
22162	:douta	=	16'h	a5db;
22163	:douta	=	16'h	9dba;
22164	:douta	=	16'h	9559;
22165	:douta	=	16'h	8d59;
22166	:douta	=	16'h	9579;
22167	:douta	=	16'h	9559;
22168	:douta	=	16'h	9d9a;
22169	:douta	=	16'h	8d38;
22170	:douta	=	16'h	9558;
22171	:douta	=	16'h	9d7a;
22172	:douta	=	16'h	84f7;
22173	:douta	=	16'h	8d38;
22174	:douta	=	16'h	9559;
22175	:douta	=	16'h	8518;
22176	:douta	=	16'h	8d18;
22177	:douta	=	16'h	84f8;
22178	:douta	=	16'h	9559;
22179	:douta	=	16'h	9dbb;
22180	:douta	=	16'h	9559;
22181	:douta	=	16'h	7c97;
22182	:douta	=	16'h	84f8;
22183	:douta	=	16'h	957a;
22184	:douta	=	16'h	9559;
22185	:douta	=	16'h	9559;
22186	:douta	=	16'h	957a;
22187	:douta	=	16'h	8d59;
22188	:douta	=	16'h	9559;
22189	:douta	=	16'h	9d9a;
22190	:douta	=	16'h	9579;
22191	:douta	=	16'h	8d18;
22192	:douta	=	16'h	7cb6;
22193	:douta	=	16'h	73b1;
22194	:douta	=	16'h	528c;
22195	:douta	=	16'h	4aad;
22196	:douta	=	16'h	5c56;
22197	:douta	=	16'h	5c57;
22198	:douta	=	16'h	32ae;
22199	:douta	=	16'h	6414;
22200	:douta	=	16'h	6c76;
22201	:douta	=	16'h	422b;
22202	:douta	=	16'h	3a09;
22203	:douta	=	16'h	5aef;
22204	:douta	=	16'h	9d9a;
22205	:douta	=	16'h	ae3d;
22206	:douta	=	16'h	8d7a;
22207	:douta	=	16'h	8539;
22208	:douta	=	16'h	8d59;
22209	:douta	=	16'h	8d7a;
22210	:douta	=	16'h	957a;
22211	:douta	=	16'h	957a;
22212	:douta	=	16'h	8d39;
22213	:douta	=	16'h	957a;
22214	:douta	=	16'h	9dbb;
22215	:douta	=	16'h	8d7a;
22216	:douta	=	16'h	8d5a;
22217	:douta	=	16'h	8d5a;
22218	:douta	=	16'h	a61c;
22219	:douta	=	16'h	8539;
22220	:douta	=	16'h	8518;
22221	:douta	=	16'h	7477;
22222	:douta	=	16'h	7cb8;
22223	:douta	=	16'h	7cd9;
22224	:douta	=	16'h	8519;
22225	:douta	=	16'h	959b;
22226	:douta	=	16'h	8d7b;
22227	:douta	=	16'h	84d9;
22228	:douta	=	16'h	853a;
22229	:douta	=	16'h	7498;
22230	:douta	=	16'h	74b8;
22231	:douta	=	16'h	7cf9;
22232	:douta	=	16'h	959b;
22233	:douta	=	16'h	9dfc;
22234	:douta	=	16'h	95bb;
22235	:douta	=	16'h	957b;
22236	:douta	=	16'h	851a;
22237	:douta	=	16'h	8d7b;
22238	:douta	=	16'h	8d5a;
22239	:douta	=	16'h	95bb;
22240	:douta	=	16'h	959c;
22241	:douta	=	16'h	7cf9;
22242	:douta	=	16'h	7cb8;
22243	:douta	=	16'h	7498;
22244	:douta	=	16'h	7cd9;
22245	:douta	=	16'h	851a;
22246	:douta	=	16'h	7d1a;
22247	:douta	=	16'h	7cd9;
22248	:douta	=	16'h	7cd9;
22249	:douta	=	16'h	85be;
22250	:douta	=	16'h	7414;
22251	:douta	=	16'h	6c55;
22252	:douta	=	16'h	7d3b;
22253	:douta	=	16'h	63f3;
22254	:douta	=	16'h	4b11;
22255	:douta	=	16'h	63f5;
22256	:douta	=	16'h	95bc;
22257	:douta	=	16'h	c6de;
22258	:douta	=	16'h	63f5;
22259	:douta	=	16'h	5bf5;
22260	:douta	=	16'h	7477;
22261	:douta	=	16'h	6c57;
22262	:douta	=	16'h	851a;
22263	:douta	=	16'h	838d;
22264	:douta	=	16'h	0000;
22265	:douta	=	16'h	28e2;
22266	:douta	=	16'h	2290;
22267	:douta	=	16'h	43b5;
22268	:douta	=	16'h	74b7;
22269	:douta	=	16'h	a5fb;
22270	:douta	=	16'h	8433;
22271	:douta	=	16'h	10a3;
22272	:douta	=	16'h	3986;
22273	:douta	=	16'h	2926;
22274	:douta	=	16'h	18e3;
22275	:douta	=	16'h	31ca;
22276	:douta	=	16'h	4bb5;
22277	:douta	=	16'h	3312;
22278	:douta	=	16'h	4374;
22279	:douta	=	16'h	4bb5;
22280	:douta	=	16'h	3ad1;
22281	:douta	=	16'h	4b53;
22282	:douta	=	16'h	6415;
22283	:douta	=	16'h	63d4;
22284	:douta	=	16'h	7477;
22285	:douta	=	16'h	6c36;
22286	:douta	=	16'h	5b72;
22287	:douta	=	16'h	6392;
22288	:douta	=	16'h	84b6;
22289	:douta	=	16'h	8d18;
22290	:douta	=	16'h	7bf2;
22291	:douta	=	16'h	c4ed;
22292	:douta	=	16'h	bced;
22293	:douta	=	16'h	d56f;
22294	:douta	=	16'h	cd8f;
22295	:douta	=	16'h	de13;
22296	:douta	=	16'h	ee75;
22297	:douta	=	16'h	ee95;
22298	:douta	=	16'h	eeb6;
22299	:douta	=	16'h	ee95;
22300	:douta	=	16'h	e654;
22301	:douta	=	16'h	e654;
22302	:douta	=	16'h	e633;
22303	:douta	=	16'h	d5b0;
22304	:douta	=	16'h	d570;
22305	:douta	=	16'h	ac4d;
22306	:douta	=	16'h	ac4c;
22307	:douta	=	16'h	bcee;
22308	:douta	=	16'h	8348;
22309	:douta	=	16'h	b4ae;
22310	:douta	=	16'h	b48d;
22311	:douta	=	16'h	b4cd;
22312	:douta	=	16'h	bccd;
22313	:douta	=	16'h	bcee;
22314	:douta	=	16'h	c4ee;
22315	:douta	=	16'h	de33;
22316	:douta	=	16'h	d5b0;
22317	:douta	=	16'h	e634;
22318	:douta	=	16'h	e654;
22319	:douta	=	16'h	e675;
22320	:douta	=	16'h	ee95;
22321	:douta	=	16'h	eeb6;
22322	:douta	=	16'h	eeb6;
22323	:douta	=	16'h	ee75;
22324	:douta	=	16'h	e654;
22325	:douta	=	16'h	e654;
22326	:douta	=	16'h	ddd1;
22327	:douta	=	16'h	d590;
22328	:douta	=	16'h	d570;
22329	:douta	=	16'h	bcb0;
22330	:douta	=	16'h	9c30;
22331	:douta	=	16'h	83d0;
22332	:douta	=	16'h	8c10;
22333	:douta	=	16'h	7370;
22334	:douta	=	16'h	6b2e;
22335	:douta	=	16'h	734f;
22336	:douta	=	16'h	732e;
22337	:douta	=	16'h	5aaa;
22338	:douta	=	16'h	4a29;
22339	:douta	=	16'h	2925;
22340	:douta	=	16'h	9308;
22341	:douta	=	16'h	a3eb;
22342	:douta	=	16'h	ac2b;
22343	:douta	=	16'h	cd2f;
22344	:douta	=	16'h	d56f;
22345	:douta	=	16'h	e613;
22346	:douta	=	16'h	ee75;
22347	:douta	=	16'h	ee95;
22348	:douta	=	16'h	eeb6;
22349	:douta	=	16'h	ee75;
22350	:douta	=	16'h	ee75;
22351	:douta	=	16'h	ee54;
22352	:douta	=	16'h	ddf2;
22353	:douta	=	16'h	cd0f;
22354	:douta	=	16'h	cd0f;
22355	:douta	=	16'h	c4cf;
22356	:douta	=	16'h	b46e;
22357	:douta	=	16'h	ac4e;
22358	:douta	=	16'h	9bee;
22359	:douta	=	16'h	93ce;
22360	:douta	=	16'h	93ef;
22361	:douta	=	16'h	8c10;
22362	:douta	=	16'h	8410;
22363	:douta	=	16'h	7bf2;
22364	:douta	=	16'h	7bf2;
22365	:douta	=	16'h	6bb2;
22366	:douta	=	16'h	63b2;
22367	:douta	=	16'h	5b91;
22368	:douta	=	16'h	4b10;
22369	:douta	=	16'h	42ce;
22370	:douta	=	16'h	320c;
22371	:douta	=	16'h	29cb;
22372	:douta	=	16'h	29aa;
22373	:douta	=	16'h	322c;
22374	:douta	=	16'h	2a0c;
22375	:douta	=	16'h	31eb;
22376	:douta	=	16'h	2146;
22377	:douta	=	16'h	3a4c;
22378	:douta	=	16'h	3a0b;
22379	:douta	=	16'h	1905;
22380	:douta	=	16'h	1926;
22381	:douta	=	16'h	1927;
22382	:douta	=	16'h	18e5;
22383	:douta	=	16'h	2147;
22384	:douta	=	16'h	1926;
22385	:douta	=	16'h	1906;
22386	:douta	=	16'h	18e5;
22387	:douta	=	16'h	18e5;
22388	:douta	=	16'h	18e5;
22389	:douta	=	16'h	18e5;
22390	:douta	=	16'h	31ea;
22391	:douta	=	16'h	10e4;
22392	:douta	=	16'h	18e5;
22393	:douta	=	16'h	0022;
22394	:douta	=	16'h	630c;
22395	:douta	=	16'h	6b6d;
22396	:douta	=	16'h	526a;
22397	:douta	=	16'h	83ee;
22398	:douta	=	16'h	8c2f;
22399	:douta	=	16'h	8bed;
22400	:douta	=	16'h	29a9;
22401	:douta	=	16'h	8518;
22402	:douta	=	16'h	84f7;
22403	:douta	=	16'h	7cb7;
22404	:douta	=	16'h	84b7;
22405	:douta	=	16'h	8d38;
22406	:douta	=	16'h	8d38;
22407	:douta	=	16'h	84f8;
22408	:douta	=	16'h	84d7;
22409	:douta	=	16'h	7476;
22410	:douta	=	16'h	7c96;
22411	:douta	=	16'h	63f4;
22412	:douta	=	16'h	8d18;
22413	:douta	=	16'h	8d18;
22414	:douta	=	16'h	84f8;
22415	:douta	=	16'h	8d38;
22416	:douta	=	16'h	84d7;
22417	:douta	=	16'h	7c96;
22418	:douta	=	16'h	84f7;
22419	:douta	=	16'h	8d18;
22420	:douta	=	16'h	9559;
22421	:douta	=	16'h	9599;
22422	:douta	=	16'h	a5fb;
22423	:douta	=	16'h	be7c;
22424	:douta	=	16'h	ae1b;
22425	:douta	=	16'h	84d8;
22426	:douta	=	16'h	a5ba;
22427	:douta	=	16'h	8d39;
22428	:douta	=	16'h	8d59;
22429	:douta	=	16'h	8d39;
22430	:douta	=	16'h	9559;
22431	:douta	=	16'h	9559;
22432	:douta	=	16'h	a5fb;
22433	:douta	=	16'h	9559;
22434	:douta	=	16'h	8d18;
22435	:douta	=	16'h	8d39;
22436	:douta	=	16'h	84f8;
22437	:douta	=	16'h	8d18;
22438	:douta	=	16'h	957a;
22439	:douta	=	16'h	8d18;
22440	:douta	=	16'h	7456;
22441	:douta	=	16'h	7476;
22442	:douta	=	16'h	8d18;
22443	:douta	=	16'h	957a;
22444	:douta	=	16'h	957a;
22445	:douta	=	16'h	8518;
22446	:douta	=	16'h	8d18;
22447	:douta	=	16'h	9d9a;
22448	:douta	=	16'h	9ddb;
22449	:douta	=	16'h	8d39;
22450	:douta	=	16'h	8539;
22451	:douta	=	16'h	853a;
22452	:douta	=	16'h	734f;
22453	:douta	=	16'h	49e6;
22454	:douta	=	16'h	4a4b;
22455	:douta	=	16'h	2188;
22456	:douta	=	16'h	2906;
22457	:douta	=	16'h	ae3e;
22458	:douta	=	16'h	9ddc;
22459	:douta	=	16'h	8d59;
22460	:douta	=	16'h	8518;
22461	:douta	=	16'h	7cf8;
22462	:douta	=	16'h	959a;
22463	:douta	=	16'h	959a;
22464	:douta	=	16'h	a5db;
22465	:douta	=	16'h	8d79;
22466	:douta	=	16'h	9d9a;
22467	:douta	=	16'h	8539;
22468	:douta	=	16'h	74b8;
22469	:douta	=	16'h	9dbb;
22470	:douta	=	16'h	8519;
22471	:douta	=	16'h	7cf8;
22472	:douta	=	16'h	8d59;
22473	:douta	=	16'h	a5db;
22474	:douta	=	16'h	8519;
22475	:douta	=	16'h	9dbb;
22476	:douta	=	16'h	959a;
22477	:douta	=	16'h	959b;
22478	:douta	=	16'h	9ddb;
22479	:douta	=	16'h	959a;
22480	:douta	=	16'h	8519;
22481	:douta	=	16'h	7498;
22482	:douta	=	16'h	853a;
22483	:douta	=	16'h	8d3a;
22484	:douta	=	16'h	7d19;
22485	:douta	=	16'h	959b;
22486	:douta	=	16'h	8d5b;
22487	:douta	=	16'h	855a;
22488	:douta	=	16'h	8d3a;
22489	:douta	=	16'h	7478;
22490	:douta	=	16'h	8d1a;
22491	:douta	=	16'h	7498;
22492	:douta	=	16'h	95bb;
22493	:douta	=	16'h	8d3a;
22494	:douta	=	16'h	957b;
22495	:douta	=	16'h	853a;
22496	:douta	=	16'h	8d9b;
22497	:douta	=	16'h	853a;
22498	:douta	=	16'h	853a;
22499	:douta	=	16'h	95bc;
22500	:douta	=	16'h	8d7b;
22501	:douta	=	16'h	7d19;
22502	:douta	=	16'h	6c56;
22503	:douta	=	16'h	74b8;
22504	:douta	=	16'h	6c98;
22505	:douta	=	16'h	52ac;
22506	:douta	=	16'h	84d8;
22507	:douta	=	16'h	32ae;
22508	:douta	=	16'h	5372;
22509	:douta	=	16'h	6415;
22510	:douta	=	16'h	8d18;
22511	:douta	=	16'h	ae1c;
22512	:douta	=	16'h	6416;
22513	:douta	=	16'h	6c76;
22514	:douta	=	16'h	5bd4;
22515	:douta	=	16'h	4b33;
22516	:douta	=	16'h	5372;
22517	:douta	=	16'h	8d18;
22518	:douta	=	16'h	9ddc;
22519	:douta	=	16'h	0000;
22520	:douta	=	16'h	b71f;
22521	:douta	=	16'h	7c96;
22522	:douta	=	16'h	6b0a;
22523	:douta	=	16'h	61e4;
22524	:douta	=	16'h	2947;
22525	:douta	=	16'h	64d9;
22526	:douta	=	16'h	7c96;
22527	:douta	=	16'h	0882;
22528	:douta	=	16'h	3166;
22529	:douta	=	16'h	3146;
22530	:douta	=	16'h	18e4;
22531	:douta	=	16'h	31c9;
22532	:douta	=	16'h	4374;
22533	:douta	=	16'h	4bb5;
22534	:douta	=	16'h	3290;
22535	:douta	=	16'h	5c16;
22536	:douta	=	16'h	2a50;
22537	:douta	=	16'h	4b53;
22538	:douta	=	16'h	5bf5;
22539	:douta	=	16'h	6c36;
22540	:douta	=	16'h	6c36;
22541	:douta	=	16'h	6c16;
22542	:douta	=	16'h	5b92;
22543	:douta	=	16'h	6392;
22544	:douta	=	16'h	7414;
22545	:douta	=	16'h	7c55;
22546	:douta	=	16'h	73d1;
22547	:douta	=	16'h	c4ed;
22548	:douta	=	16'h	c50e;
22549	:douta	=	16'h	d56f;
22550	:douta	=	16'h	cd8f;
22551	:douta	=	16'h	e613;
22552	:douta	=	16'h	ee95;
22553	:douta	=	16'h	ee95;
22554	:douta	=	16'h	f6b6;
22555	:douta	=	16'h	f6d7;
22556	:douta	=	16'h	e654;
22557	:douta	=	16'h	e633;
22558	:douta	=	16'h	ddf2;
22559	:douta	=	16'h	d56f;
22560	:douta	=	16'h	cd2f;
22561	:douta	=	16'h	ac4b;
22562	:douta	=	16'h	9baa;
22563	:douta	=	16'h	7ae7;
22564	:douta	=	16'h	b48d;
22565	:douta	=	16'h	ac6d;
22566	:douta	=	16'h	bd2e;
22567	:douta	=	16'h	bd0d;
22568	:douta	=	16'h	bcee;
22569	:douta	=	16'h	cd4f;
22570	:douta	=	16'h	cd6f;
22571	:douta	=	16'h	e655;
22572	:douta	=	16'h	d5b0;
22573	:douta	=	16'h	e654;
22574	:douta	=	16'h	eeb6;
22575	:douta	=	16'h	ee75;
22576	:douta	=	16'h	eeb6;
22577	:douta	=	16'h	e675;
22578	:douta	=	16'h	ee96;
22579	:douta	=	16'h	ee95;
22580	:douta	=	16'h	e654;
22581	:douta	=	16'h	e613;
22582	:douta	=	16'h	ddb2;
22583	:douta	=	16'h	cd50;
22584	:douta	=	16'h	cd30;
22585	:douta	=	16'h	c4f0;
22586	:douta	=	16'h	8bd0;
22587	:douta	=	16'h	7bb0;
22588	:douta	=	16'h	7bd0;
22589	:douta	=	16'h	736f;
22590	:douta	=	16'h	6b2f;
22591	:douta	=	16'h	6b2d;
22592	:douta	=	16'h	7b8f;
22593	:douta	=	16'h	62cc;
22594	:douta	=	16'h	28e3;
22595	:douta	=	16'h	51a5;
22596	:douta	=	16'h	9be9;
22597	:douta	=	16'h	b46b;
22598	:douta	=	16'h	c4ee;
22599	:douta	=	16'h	d5b1;
22600	:douta	=	16'h	ddf2;
22601	:douta	=	16'h	ee95;
22602	:douta	=	16'h	ee96;
22603	:douta	=	16'h	eeb6;
22604	:douta	=	16'h	ee95;
22605	:douta	=	16'h	ee75;
22606	:douta	=	16'h	e634;
22607	:douta	=	16'h	e634;
22608	:douta	=	16'h	ddf2;
22609	:douta	=	16'h	cd2f;
22610	:douta	=	16'h	cd0f;
22611	:douta	=	16'h	bcae;
22612	:douta	=	16'h	ac4e;
22613	:douta	=	16'h	ac2e;
22614	:douta	=	16'h	a42e;
22615	:douta	=	16'h	a42f;
22616	:douta	=	16'h	8c10;
22617	:douta	=	16'h	8c10;
22618	:douta	=	16'h	8c11;
22619	:douta	=	16'h	8412;
22620	:douta	=	16'h	8433;
22621	:douta	=	16'h	7c13;
22622	:douta	=	16'h	7414;
22623	:douta	=	16'h	63b2;
22624	:douta	=	16'h	5b51;
22625	:douta	=	16'h	5330;
22626	:douta	=	16'h	428e;
22627	:douta	=	16'h	3a8d;
22628	:douta	=	16'h	3a6d;
22629	:douta	=	16'h	42ef;
22630	:douta	=	16'h	3af0;
22631	:douta	=	16'h	31c9;
22632	:douta	=	16'h	31c9;
22633	:douta	=	16'h	2168;
22634	:douta	=	16'h	42ae;
22635	:douta	=	16'h	5310;
22636	:douta	=	16'h	1927;
22637	:douta	=	16'h	2147;
22638	:douta	=	16'h	18e5;
22639	:douta	=	16'h	1906;
22640	:douta	=	16'h	1926;
22641	:douta	=	16'h	1926;
22642	:douta	=	16'h	1925;
22643	:douta	=	16'h	18e5;
22644	:douta	=	16'h	1905;
22645	:douta	=	16'h	18e5;
22646	:douta	=	16'h	10c5;
22647	:douta	=	16'h	18e5;
22648	:douta	=	16'h	10e5;
22649	:douta	=	16'h	18c5;
22650	:douta	=	16'h	0001;
22651	:douta	=	16'h	2987;
22652	:douta	=	16'h	7b6e;
22653	:douta	=	16'h	2126;
22654	:douta	=	16'h	5acb;
22655	:douta	=	16'h	9c70;
22656	:douta	=	16'h	4a28;
22657	:douta	=	16'h	31c9;
22658	:douta	=	16'h	ae3d;
22659	:douta	=	16'h	7c96;
22660	:douta	=	16'h	7455;
22661	:douta	=	16'h	9559;
22662	:douta	=	16'h	9579;
22663	:douta	=	16'h	9d9a;
22664	:douta	=	16'h	84f8;
22665	:douta	=	16'h	84d7;
22666	:douta	=	16'h	7c96;
22667	:douta	=	16'h	7455;
22668	:douta	=	16'h	7c76;
22669	:douta	=	16'h	84b7;
22670	:douta	=	16'h	8d18;
22671	:douta	=	16'h	9559;
22672	:douta	=	16'h	9579;
22673	:douta	=	16'h	84b7;
22674	:douta	=	16'h	84d7;
22675	:douta	=	16'h	84d7;
22676	:douta	=	16'h	84b6;
22677	:douta	=	16'h	84d7;
22678	:douta	=	16'h	9539;
22679	:douta	=	16'h	adda;
22680	:douta	=	16'h	b63b;
22681	:douta	=	16'h	9579;
22682	:douta	=	16'h	8d18;
22683	:douta	=	16'h	8d39;
22684	:douta	=	16'h	9559;
22685	:douta	=	16'h	8d39;
22686	:douta	=	16'h	957a;
22687	:douta	=	16'h	8d39;
22688	:douta	=	16'h	7cb7;
22689	:douta	=	16'h	84f8;
22690	:douta	=	16'h	8d59;
22691	:douta	=	16'h	9559;
22692	:douta	=	16'h	955a;
22693	:douta	=	16'h	84f8;
22694	:douta	=	16'h	8518;
22695	:douta	=	16'h	8d59;
22696	:douta	=	16'h	84f8;
22697	:douta	=	16'h	84f8;
22698	:douta	=	16'h	6c55;
22699	:douta	=	16'h	6c15;
22700	:douta	=	16'h	84f9;
22701	:douta	=	16'h	959a;
22702	:douta	=	16'h	8d39;
22703	:douta	=	16'h	8d59;
22704	:douta	=	16'h	84f8;
22705	:douta	=	16'h	9ddb;
22706	:douta	=	16'h	957a;
22707	:douta	=	16'h	8d5a;
22708	:douta	=	16'h	8432;
22709	:douta	=	16'h	7b09;
22710	:douta	=	16'h	4a6b;
22711	:douta	=	16'h	1041;
22712	:douta	=	16'h	39e9;
22713	:douta	=	16'h	9dbb;
22714	:douta	=	16'h	8519;
22715	:douta	=	16'h	959a;
22716	:douta	=	16'h	9d9a;
22717	:douta	=	16'h	8539;
22718	:douta	=	16'h	957a;
22719	:douta	=	16'h	957a;
22720	:douta	=	16'h	957a;
22721	:douta	=	16'h	a61b;
22722	:douta	=	16'h	959a;
22723	:douta	=	16'h	9dbb;
22724	:douta	=	16'h	8d59;
22725	:douta	=	16'h	9ddb;
22726	:douta	=	16'h	9dbb;
22727	:douta	=	16'h	957a;
22728	:douta	=	16'h	957a;
22729	:douta	=	16'h	a5db;
22730	:douta	=	16'h	9ddb;
22731	:douta	=	16'h	8d7a;
22732	:douta	=	16'h	9dbb;
22733	:douta	=	16'h	957a;
22734	:douta	=	16'h	959b;
22735	:douta	=	16'h	959a;
22736	:douta	=	16'h	a61c;
22737	:douta	=	16'h	8d59;
22738	:douta	=	16'h	7cf9;
22739	:douta	=	16'h	8519;
22740	:douta	=	16'h	7cf9;
22741	:douta	=	16'h	8d7b;
22742	:douta	=	16'h	957a;
22743	:douta	=	16'h	853a;
22744	:douta	=	16'h	7cd9;
22745	:douta	=	16'h	8d3a;
22746	:douta	=	16'h	8d5a;
22747	:douta	=	16'h	7cd8;
22748	:douta	=	16'h	7cd9;
22749	:douta	=	16'h	7498;
22750	:douta	=	16'h	8d3a;
22751	:douta	=	16'h	9e1d;
22752	:douta	=	16'h	9e1e;
22753	:douta	=	16'h	959c;
22754	:douta	=	16'h	853a;
22755	:douta	=	16'h	8d5b;
22756	:douta	=	16'h	8d7b;
22757	:douta	=	16'h	8d5a;
22758	:douta	=	16'h	8d7b;
22759	:douta	=	16'h	7d7c;
22760	:douta	=	16'h	6b2c;
22761	:douta	=	16'h	53d4;
22762	:douta	=	16'h	9dfd;
22763	:douta	=	16'h	74b9;
22764	:douta	=	16'h	74b9;
22765	:douta	=	16'h	7c56;
22766	:douta	=	16'h	7cb7;
22767	:douta	=	16'h	6c57;
22768	:douta	=	16'h	5bd4;
22769	:douta	=	16'h	8519;
22770	:douta	=	16'h	9dbb;
22771	:douta	=	16'h	6c35;
22772	:douta	=	16'h	9d7a;
22773	:douta	=	16'h	5bf5;
22774	:douta	=	16'h	5394;
22775	:douta	=	16'h	1860;
22776	:douta	=	16'h	8d5a;
22777	:douta	=	16'h	8d7b;
22778	:douta	=	16'h	95bb;
22779	:douta	=	16'h	84b6;
22780	:douta	=	16'h	7225;
22781	:douta	=	16'h	3145;
22782	:douta	=	16'h	3a4c;
22783	:douta	=	16'h	1883;
22784	:douta	=	16'h	3166;
22785	:douta	=	16'h	3146;
22786	:douta	=	16'h	2945;
22787	:douta	=	16'h	2126;
22788	:douta	=	16'h	326f;
22789	:douta	=	16'h	3b33;
22790	:douta	=	16'h	2a2e;
22791	:douta	=	16'h	4333;
22792	:douta	=	16'h	32b0;
22793	:douta	=	16'h	4b53;
22794	:douta	=	16'h	6c36;
22795	:douta	=	16'h	4b11;
22796	:douta	=	16'h	63f4;
22797	:douta	=	16'h	5bb4;
22798	:douta	=	16'h	6392;
22799	:douta	=	16'h	63b3;
22800	:douta	=	16'h	9518;
22801	:douta	=	16'h	63f4;
22802	:douta	=	16'h	7c54;
22803	:douta	=	16'h	c50d;
22804	:douta	=	16'h	c54e;
22805	:douta	=	16'h	cd70;
22806	:douta	=	16'h	ddd3;
22807	:douta	=	16'h	e654;
22808	:douta	=	16'h	ee95;
22809	:douta	=	16'h	eeb6;
22810	:douta	=	16'h	eeb6;
22811	:douta	=	16'h	e675;
22812	:douta	=	16'h	ee75;
22813	:douta	=	16'h	d5b1;
22814	:douta	=	16'h	ddd0;
22815	:douta	=	16'h	c4cf;
22816	:douta	=	16'h	ac6d;
22817	:douta	=	16'h	938a;
22818	:douta	=	16'h	72c6;
22819	:douta	=	16'h	a42c;
22820	:douta	=	16'h	b4ed;
22821	:douta	=	16'h	b4ad;
22822	:douta	=	16'h	c54f;
22823	:douta	=	16'h	d591;
22824	:douta	=	16'h	bd0e;
22825	:douta	=	16'h	ddf2;
22826	:douta	=	16'h	e675;
22827	:douta	=	16'h	ee95;
22828	:douta	=	16'h	ddf2;
22829	:douta	=	16'h	ddf2;
22830	:douta	=	16'h	ee96;
22831	:douta	=	16'h	eeb6;
22832	:douta	=	16'h	e654;
22833	:douta	=	16'h	ee95;
22834	:douta	=	16'h	e654;
22835	:douta	=	16'h	ee54;
22836	:douta	=	16'h	e654;
22837	:douta	=	16'h	ddd1;
22838	:douta	=	16'h	c52f;
22839	:douta	=	16'h	d550;
22840	:douta	=	16'h	ac6f;
22841	:douta	=	16'h	9c10;
22842	:douta	=	16'h	8bf0;
22843	:douta	=	16'h	7bb0;
22844	:douta	=	16'h	736f;
22845	:douta	=	16'h	62ed;
22846	:douta	=	16'h	62ed;
22847	:douta	=	16'h	5a6a;
22848	:douta	=	16'h	4a2a;
22849	:douta	=	16'h	2904;
22850	:douta	=	16'h	abca;
22851	:douta	=	16'h	b46c;
22852	:douta	=	16'h	b46c;
22853	:douta	=	16'h	cd2d;
22854	:douta	=	16'h	d5b0;
22855	:douta	=	16'h	e613;
22856	:douta	=	16'h	e675;
22857	:douta	=	16'h	ee96;
22858	:douta	=	16'h	ee95;
22859	:douta	=	16'h	ee75;
22860	:douta	=	16'h	ee75;
22861	:douta	=	16'h	ee75;
22862	:douta	=	16'h	e613;
22863	:douta	=	16'h	ddd2;
22864	:douta	=	16'h	d591;
22865	:douta	=	16'h	cd0f;
22866	:douta	=	16'h	bccf;
22867	:douta	=	16'h	bccf;
22868	:douta	=	16'h	b46f;
22869	:douta	=	16'h	b46e;
22870	:douta	=	16'h	a450;
22871	:douta	=	16'h	9410;
22872	:douta	=	16'h	9431;
22873	:douta	=	16'h	8c31;
22874	:douta	=	16'h	9432;
22875	:douta	=	16'h	8c73;
22876	:douta	=	16'h	8433;
22877	:douta	=	16'h	7c13;
22878	:douta	=	16'h	7c13;
22879	:douta	=	16'h	7434;
22880	:douta	=	16'h	73f2;
22881	:douta	=	16'h	6bd2;
22882	:douta	=	16'h	6bb2;
22883	:douta	=	16'h	6392;
22884	:douta	=	16'h	5bb3;
22885	:douta	=	16'h	0909;
22886	:douta	=	16'h	3925;
22887	:douta	=	16'h	4b0e;
22888	:douta	=	16'h	320c;
22889	:douta	=	16'h	4a8e;
22890	:douta	=	16'h	1947;
22891	:douta	=	16'h	0042;
22892	:douta	=	16'h	42af;
22893	:douta	=	16'h	1905;
22894	:douta	=	16'h	0883;
22895	:douta	=	16'h	10a4;
22896	:douta	=	16'h	1083;
22897	:douta	=	16'h	10a4;
22898	:douta	=	16'h	10c5;
22899	:douta	=	16'h	1905;
22900	:douta	=	16'h	18e5;
22901	:douta	=	16'h	18e5;
22902	:douta	=	16'h	1905;
22903	:douta	=	16'h	1084;
22904	:douta	=	16'h	1906;
22905	:douta	=	16'h	18c4;
22906	:douta	=	16'h	2106;
22907	:douta	=	16'h	10e4;
22908	:douta	=	16'h	0001;
22909	:douta	=	16'h	736d;
22910	:douta	=	16'h	ce14;
22911	:douta	=	16'h	de97;
22912	:douta	=	16'h	9491;
22913	:douta	=	16'h	4a8c;
22914	:douta	=	16'h	3147;
22915	:douta	=	16'h	9d7a;
22916	:douta	=	16'h	adfc;
22917	:douta	=	16'h	7cb7;
22918	:douta	=	16'h	84b7;
22919	:douta	=	16'h	7cb7;
22920	:douta	=	16'h	9d9a;
22921	:douta	=	16'h	959a;
22922	:douta	=	16'h	9d7a;
22923	:douta	=	16'h	9599;
22924	:douta	=	16'h	9599;
22925	:douta	=	16'h	84f8;
22926	:douta	=	16'h	84f8;
22927	:douta	=	16'h	84d6;
22928	:douta	=	16'h	7c95;
22929	:douta	=	16'h	6c14;
22930	:douta	=	16'h	8cf8;
22931	:douta	=	16'h	8d18;
22932	:douta	=	16'h	84d7;
22933	:douta	=	16'h	8d18;
22934	:douta	=	16'h	7455;
22935	:douta	=	16'h	84d7;
22936	:douta	=	16'h	7476;
22937	:douta	=	16'h	7455;
22938	:douta	=	16'h	7476;
22939	:douta	=	16'h	a5db;
22940	:douta	=	16'h	9d9a;
22941	:douta	=	16'h	9dba;
22942	:douta	=	16'h	8d18;
22943	:douta	=	16'h	8d19;
22944	:douta	=	16'h	8d59;
22945	:douta	=	16'h	9559;
22946	:douta	=	16'h	8d39;
22947	:douta	=	16'h	84d7;
22948	:douta	=	16'h	7cd7;
22949	:douta	=	16'h	84b7;
22950	:douta	=	16'h	8d59;
22951	:douta	=	16'h	8518;
22952	:douta	=	16'h	957a;
22953	:douta	=	16'h	84f8;
22954	:douta	=	16'h	8d39;
22955	:douta	=	16'h	957a;
22956	:douta	=	16'h	8d5a;
22957	:douta	=	16'h	7497;
22958	:douta	=	16'h	7476;
22959	:douta	=	16'h	84f8;
22960	:douta	=	16'h	8d59;
22961	:douta	=	16'h	8d7a;
22962	:douta	=	16'h	8d59;
22963	:douta	=	16'h	8d19;
22964	:douta	=	16'h	8c52;
22965	:douta	=	16'h	8b6b;
22966	:douta	=	16'h	4a8c;
22967	:douta	=	16'h	1882;
22968	:douta	=	16'h	39e9;
22969	:douta	=	16'h	7cb8;
22970	:douta	=	16'h	84f8;
22971	:douta	=	16'h	9dbb;
22972	:douta	=	16'h	9559;
22973	:douta	=	16'h	95bb;
22974	:douta	=	16'h	9d9a;
22975	:douta	=	16'h	959a;
22976	:douta	=	16'h	9dda;
22977	:douta	=	16'h	8d18;
22978	:douta	=	16'h	7c97;
22979	:douta	=	16'h	8d59;
22980	:douta	=	16'h	959a;
22981	:douta	=	16'h	74b8;
22982	:douta	=	16'h	a5fb;
22983	:douta	=	16'h	9dbb;
22984	:douta	=	16'h	7d19;
22985	:douta	=	16'h	8d7a;
22986	:douta	=	16'h	95ba;
22987	:douta	=	16'h	95bb;
22988	:douta	=	16'h	957b;
22989	:douta	=	16'h	957a;
22990	:douta	=	16'h	8d5a;
22991	:douta	=	16'h	959b;
22992	:douta	=	16'h	9dbb;
22993	:douta	=	16'h	959a;
22994	:douta	=	16'h	9ddb;
22995	:douta	=	16'h	957a;
22996	:douta	=	16'h	a5fc;
22997	:douta	=	16'h	7477;
22998	:douta	=	16'h	7457;
22999	:douta	=	16'h	7cd8;
23000	:douta	=	16'h	8d7a;
23001	:douta	=	16'h	959b;
23002	:douta	=	16'h	84f9;
23003	:douta	=	16'h	8d3a;
23004	:douta	=	16'h	8d5a;
23005	:douta	=	16'h	9d9a;
23006	:douta	=	16'h	7d19;
23007	:douta	=	16'h	7477;
23008	:douta	=	16'h	7cb8;
23009	:douta	=	16'h	7cf9;
23010	:douta	=	16'h	8519;
23011	:douta	=	16'h	8d7b;
23012	:douta	=	16'h	851a;
23013	:douta	=	16'h	8d5b;
23014	:douta	=	16'h	851a;
23015	:douta	=	16'h	632e;
23016	:douta	=	16'h	328d;
23017	:douta	=	16'h	5921;
23018	:douta	=	16'h	2168;
23019	:douta	=	16'h	3af1;
23020	:douta	=	16'h	5372;
23021	:douta	=	16'h	6c56;
23022	:douta	=	16'h	9539;
23023	:douta	=	16'h	6c57;
23024	:douta	=	16'h	74b7;
23025	:douta	=	16'h	8d39;
23026	:douta	=	16'h	4311;
23027	:douta	=	16'h	4311;
23028	:douta	=	16'h	5bd4;
23029	:douta	=	16'h	84fa;
23030	:douta	=	16'h	6b4e;
23031	:douta	=	16'h	63f4;
23032	:douta	=	16'h	5b94;
23033	:douta	=	16'h	5bf4;
23034	:douta	=	16'h	7455;
23035	:douta	=	16'h	7456;
23036	:douta	=	16'h	6415;
23037	:douta	=	16'h	7477;
23038	:douta	=	16'h	8c52;
23039	:douta	=	16'h	5a25;
23040	:douta	=	16'h	3986;
23041	:douta	=	16'h	3165;
23042	:douta	=	16'h	2925;
23043	:douta	=	16'h	31a8;
23044	:douta	=	16'h	2a6f;
23045	:douta	=	16'h	4c18;
23046	:douta	=	16'h	2a4e;
23047	:douta	=	16'h	3b12;
23048	:douta	=	16'h	32b0;
23049	:douta	=	16'h	4353;
23050	:douta	=	16'h	6436;
23051	:douta	=	16'h	5352;
23052	:douta	=	16'h	7455;
23053	:douta	=	16'h	7476;
23054	:douta	=	16'h	6393;
23055	:douta	=	16'h	5b72;
23056	:douta	=	16'h	7434;
23057	:douta	=	16'h	7455;
23058	:douta	=	16'h	7c13;
23059	:douta	=	16'h	cd2e;
23060	:douta	=	16'h	cd6f;
23061	:douta	=	16'h	d590;
23062	:douta	=	16'h	ddf2;
23063	:douta	=	16'h	ee75;
23064	:douta	=	16'h	eeb6;
23065	:douta	=	16'h	eeb6;
23066	:douta	=	16'h	ee75;
23067	:douta	=	16'h	e654;
23068	:douta	=	16'h	ee95;
23069	:douta	=	16'h	b4cd;
23070	:douta	=	16'h	ac6d;
23071	:douta	=	16'h	b46e;
23072	:douta	=	16'h	b48d;
23073	:douta	=	16'h	7ae7;
23074	:douta	=	16'h	a42c;
23075	:douta	=	16'h	b4ad;
23076	:douta	=	16'h	accd;
23077	:douta	=	16'h	c56f;
23078	:douta	=	16'h	c52e;
23079	:douta	=	16'h	de13;
23080	:douta	=	16'h	c54f;
23081	:douta	=	16'h	e654;
23082	:douta	=	16'h	e676;
23083	:douta	=	16'h	ee96;
23084	:douta	=	16'h	e654;
23085	:douta	=	16'h	de12;
23086	:douta	=	16'h	ee96;
23087	:douta	=	16'h	ee96;
23088	:douta	=	16'h	e633;
23089	:douta	=	16'h	ee75;
23090	:douta	=	16'h	e675;
23091	:douta	=	16'h	e613;
23092	:douta	=	16'h	e633;
23093	:douta	=	16'h	ddf1;
23094	:douta	=	16'h	b4af;
23095	:douta	=	16'h	b48f;
23096	:douta	=	16'h	ac8f;
23097	:douta	=	16'h	9430;
23098	:douta	=	16'h	83cf;
23099	:douta	=	16'h	734f;
23100	:douta	=	16'h	732e;
23101	:douta	=	16'h	6b0c;
23102	:douta	=	16'h	62ec;
23103	:douta	=	16'h	5aab;
23104	:douta	=	16'h	20c4;
23105	:douta	=	16'h	59c4;
23106	:douta	=	16'h	b46c;
23107	:douta	=	16'h	ac4c;
23108	:douta	=	16'h	bccc;
23109	:douta	=	16'h	d58f;
23110	:douta	=	16'h	e612;
23111	:douta	=	16'h	e654;
23112	:douta	=	16'h	ee75;
23113	:douta	=	16'h	eeb6;
23114	:douta	=	16'h	eeb6;
23115	:douta	=	16'h	eeb6;
23116	:douta	=	16'h	e655;
23117	:douta	=	16'h	e655;
23118	:douta	=	16'h	e613;
23119	:douta	=	16'h	ddd2;
23120	:douta	=	16'h	ddb2;
23121	:douta	=	16'h	c4ef;
23122	:douta	=	16'h	bccf;
23123	:douta	=	16'h	bcaf;
23124	:douta	=	16'h	ac6e;
23125	:douta	=	16'h	ac4f;
23126	:douta	=	16'h	8bef;
23127	:douta	=	16'h	9410;
23128	:douta	=	16'h	9451;
23129	:douta	=	16'h	9c72;
23130	:douta	=	16'h	9452;
23131	:douta	=	16'h	9473;
23132	:douta	=	16'h	8c53;
23133	:douta	=	16'h	8474;
23134	:douta	=	16'h	8454;
23135	:douta	=	16'h	7c54;
23136	:douta	=	16'h	7414;
23137	:douta	=	16'h	73d3;
23138	:douta	=	16'h	6bd2;
23139	:douta	=	16'h	6bf2;
23140	:douta	=	16'h	4b32;
23141	:douta	=	16'h	8b09;
23142	:douta	=	16'h	b46f;
23143	:douta	=	16'h	42ae;
23144	:douta	=	16'h	322b;
23145	:douta	=	16'h	4aae;
23146	:douta	=	16'h	31ea;
23147	:douta	=	16'h	1906;
23148	:douta	=	16'h	2988;
23149	:douta	=	16'h	29c9;
23150	:douta	=	16'h	0863;
23151	:douta	=	16'h	0883;
23152	:douta	=	16'h	10a3;
23153	:douta	=	16'h	10a3;
23154	:douta	=	16'h	10c3;
23155	:douta	=	16'h	10a4;
23156	:douta	=	16'h	10c4;
23157	:douta	=	16'h	18e5;
23158	:douta	=	16'h	18e5;
23159	:douta	=	16'h	1905;
23160	:douta	=	16'h	10c4;
23161	:douta	=	16'h	10a4;
23162	:douta	=	16'h	10a3;
23163	:douta	=	16'h	18e5;
23164	:douta	=	16'h	1905;
23165	:douta	=	16'h	0022;
23166	:douta	=	16'h	bd72;
23167	:douta	=	16'h	8430;
23168	:douta	=	16'h	9491;
23169	:douta	=	16'h	5b0c;
23170	:douta	=	16'h	d635;
23171	:douta	=	16'h	31eb;
23172	:douta	=	16'h	7cb7;
23173	:douta	=	16'h	9579;
23174	:douta	=	16'h	8d38;
23175	:douta	=	16'h	8d18;
23176	:douta	=	16'h	9d9a;
23177	:douta	=	16'h	9559;
23178	:douta	=	16'h	84f8;
23179	:douta	=	16'h	7cb7;
23180	:douta	=	16'h	9d7a;
23181	:douta	=	16'h	9559;
23182	:douta	=	16'h	8d38;
23183	:douta	=	16'h	9579;
23184	:douta	=	16'h	9559;
23185	:douta	=	16'h	8cf8;
23186	:douta	=	16'h	7434;
23187	:douta	=	16'h	63d3;
23188	:douta	=	16'h	84d7;
23189	:douta	=	16'h	9539;
23190	:douta	=	16'h	8d18;
23191	:douta	=	16'h	7c96;
23192	:douta	=	16'h	7c97;
23193	:douta	=	16'h	7c97;
23194	:douta	=	16'h	6c15;
23195	:douta	=	16'h	6c35;
23196	:douta	=	16'h	8518;
23197	:douta	=	16'h	957a;
23198	:douta	=	16'h	9559;
23199	:douta	=	16'h	959a;
23200	:douta	=	16'h	959a;
23201	:douta	=	16'h	84f8;
23202	:douta	=	16'h	7cb7;
23203	:douta	=	16'h	8518;
23204	:douta	=	16'h	8518;
23205	:douta	=	16'h	8d19;
23206	:douta	=	16'h	7cb7;
23207	:douta	=	16'h	7cd8;
23208	:douta	=	16'h	8518;
23209	:douta	=	16'h	8d39;
23210	:douta	=	16'h	955a;
23211	:douta	=	16'h	8d39;
23212	:douta	=	16'h	8539;
23213	:douta	=	16'h	8d7a;
23214	:douta	=	16'h	957a;
23215	:douta	=	16'h	7cd7;
23216	:douta	=	16'h	7cd8;
23217	:douta	=	16'h	84f8;
23218	:douta	=	16'h	959a;
23219	:douta	=	16'h	8d59;
23220	:douta	=	16'h	9473;
23221	:douta	=	16'h	834b;
23222	:douta	=	16'h	4a6c;
23223	:douta	=	16'h	1062;
23224	:douta	=	16'h	39e9;
23225	:douta	=	16'h	95bb;
23226	:douta	=	16'h	8519;
23227	:douta	=	16'h	8d59;
23228	:douta	=	16'h	7cf8;
23229	:douta	=	16'h	8d5a;
23230	:douta	=	16'h	9ddb;
23231	:douta	=	16'h	959a;
23232	:douta	=	16'h	9dbb;
23233	:douta	=	16'h	b65d;
23234	:douta	=	16'h	ae3c;
23235	:douta	=	16'h	8539;
23236	:douta	=	16'h	8539;
23237	:douta	=	16'h	9dbb;
23238	:douta	=	16'h	8539;
23239	:douta	=	16'h	959a;
23240	:douta	=	16'h	8d39;
23241	:douta	=	16'h	8d39;
23242	:douta	=	16'h	959b;
23243	:douta	=	16'h	9ddb;
23244	:douta	=	16'h	7cf9;
23245	:douta	=	16'h	a5fc;
23246	:douta	=	16'h	a5fb;
23247	:douta	=	16'h	959b;
23248	:douta	=	16'h	8d5a;
23249	:douta	=	16'h	959a;
23250	:douta	=	16'h	a61c;
23251	:douta	=	16'h	a5fb;
23252	:douta	=	16'h	8539;
23253	:douta	=	16'h	a61d;
23254	:douta	=	16'h	a5fc;
23255	:douta	=	16'h	7497;
23256	:douta	=	16'h	7497;
23257	:douta	=	16'h	8519;
23258	:douta	=	16'h	9dbb;
23259	:douta	=	16'h	957b;
23260	:douta	=	16'h	95bb;
23261	:douta	=	16'h	95bb;
23262	:douta	=	16'h	8d3a;
23263	:douta	=	16'h	8519;
23264	:douta	=	16'h	7cd9;
23265	:douta	=	16'h	7cd9;
23266	:douta	=	16'h	7cd8;
23267	:douta	=	16'h	853a;
23268	:douta	=	16'h	7d3a;
23269	:douta	=	16'h	8dbc;
23270	:douta	=	16'h	524a;
23271	:douta	=	16'h	0000;
23272	:douta	=	16'h	2127;
23273	:douta	=	16'h	7bef;
23274	:douta	=	16'h	4921;
23275	:douta	=	16'h	74fa;
23276	:douta	=	16'h	95dc;
23277	:douta	=	16'h	8d5a;
23278	:douta	=	16'h	53b4;
23279	:douta	=	16'h	53b4;
23280	:douta	=	16'h	9dbc;
23281	:douta	=	16'h	8d19;
23282	:douta	=	16'h	9dbb;
23283	:douta	=	16'h	8d39;
23284	:douta	=	16'h	8518;
23285	:douta	=	16'h	84d7;
23286	:douta	=	16'h	5184;
23287	:douta	=	16'h	53f5;
23288	:douta	=	16'h	7477;
23289	:douta	=	16'h	8539;
23290	:douta	=	16'h	cefe;
23291	:douta	=	16'h	8d19;
23292	:douta	=	16'h	8d39;
23293	:douta	=	16'h	5bf5;
23294	:douta	=	16'h	6cba;
23295	:douta	=	16'h	3964;
23296	:douta	=	16'h	3966;
23297	:douta	=	16'h	3145;
23298	:douta	=	16'h	3145;
23299	:douta	=	16'h	1083;
23300	:douta	=	16'h	32d1;
23301	:douta	=	16'h	32d1;
23302	:douta	=	16'h	32b1;
23303	:douta	=	16'h	32b1;
23304	:douta	=	16'h	4353;
23305	:douta	=	16'h	53b5;
23306	:douta	=	16'h	5394;
23307	:douta	=	16'h	7456;
23308	:douta	=	16'h	7cb7;
23309	:douta	=	16'h	7cb8;
23310	:douta	=	16'h	63f5;
23311	:douta	=	16'h	6372;
23312	:douta	=	16'h	7c55;
23313	:douta	=	16'h	8496;
23314	:douta	=	16'h	6bd2;
23315	:douta	=	16'h	bcef;
23316	:douta	=	16'h	d58e;
23317	:douta	=	16'h	ddf3;
23318	:douta	=	16'h	e654;
23319	:douta	=	16'h	ee76;
23320	:douta	=	16'h	eeb6;
23321	:douta	=	16'h	ee95;
23322	:douta	=	16'h	e634;
23323	:douta	=	16'h	e613;
23324	:douta	=	16'h	d570;
23325	:douta	=	16'h	cd70;
23326	:douta	=	16'h	cd70;
23327	:douta	=	16'h	7b07;
23328	:douta	=	16'h	51c4;
23329	:douta	=	16'h	b48d;
23330	:douta	=	16'h	b4ad;
23331	:douta	=	16'h	bcee;
23332	:douta	=	16'h	d5b1;
23333	:douta	=	16'h	d613;
23334	:douta	=	16'h	d5b1;
23335	:douta	=	16'h	d5d3;
23336	:douta	=	16'h	c570;
23337	:douta	=	16'h	e675;
23338	:douta	=	16'h	eeb6;
23339	:douta	=	16'h	ddf3;
23340	:douta	=	16'h	f6f8;
23341	:douta	=	16'h	eeb7;
23342	:douta	=	16'h	e675;
23343	:douta	=	16'h	ee95;
23344	:douta	=	16'h	e654;
23345	:douta	=	16'h	e613;
23346	:douta	=	16'h	e613;
23347	:douta	=	16'h	de12;
23348	:douta	=	16'h	d5b1;
23349	:douta	=	16'h	cd2f;
23350	:douta	=	16'h	b4ae;
23351	:douta	=	16'h	a46f;
23352	:douta	=	16'h	83af;
23353	:douta	=	16'h	838f;
23354	:douta	=	16'h	7b8f;
23355	:douta	=	16'h	6b2c;
23356	:douta	=	16'h	62ec;
23357	:douta	=	16'h	5a6b;
23358	:douta	=	16'h	5a6a;
23359	:douta	=	16'h	3145;
23360	:douta	=	16'h	a388;
23361	:douta	=	16'h	ac4a;
23362	:douta	=	16'h	b46b;
23363	:douta	=	16'h	c4cc;
23364	:douta	=	16'h	ddd1;
23365	:douta	=	16'h	e654;
23366	:douta	=	16'h	e634;
23367	:douta	=	16'h	de33;
23368	:douta	=	16'h	e654;
23369	:douta	=	16'h	e654;
23370	:douta	=	16'h	eeb6;
23371	:douta	=	16'h	eeb6;
23372	:douta	=	16'h	e654;
23373	:douta	=	16'h	e654;
23374	:douta	=	16'h	e613;
23375	:douta	=	16'h	d572;
23376	:douta	=	16'h	cd71;
23377	:douta	=	16'h	c510;
23378	:douta	=	16'h	bcb0;
23379	:douta	=	16'h	ac50;
23380	:douta	=	16'h	9c30;
23381	:douta	=	16'h	9430;
23382	:douta	=	16'h	9451;
23383	:douta	=	16'h	8c31;
23384	:douta	=	16'h	8c11;
23385	:douta	=	16'h	8432;
23386	:douta	=	16'h	8c32;
23387	:douta	=	16'h	8412;
23388	:douta	=	16'h	8412;
23389	:douta	=	16'h	7bf2;
23390	:douta	=	16'h	73b1;
23391	:douta	=	16'h	736f;
23392	:douta	=	16'h	632e;
23393	:douta	=	16'h	52ac;
23394	:douta	=	16'h	62ac;
23395	:douta	=	16'h	6a8a;
23396	:douta	=	16'h	d52b;
23397	:douta	=	16'h	de13;
23398	:douta	=	16'h	a48f;
23399	:douta	=	16'h	4ace;
23400	:douta	=	16'h	29eb;
23401	:douta	=	16'h	632e;
23402	:douta	=	16'h	3a8c;
23403	:douta	=	16'h	2147;
23404	:douta	=	16'h	1905;
23405	:douta	=	16'h	10c5;
23406	:douta	=	16'h	2947;
23407	:douta	=	16'h	5b0e;
23408	:douta	=	16'h	39ea;
23409	:douta	=	16'h	1083;
23410	:douta	=	16'h	10c5;
23411	:douta	=	16'h	10e5;
23412	:douta	=	16'h	18e5;
23413	:douta	=	16'h	18e5;
23414	:douta	=	16'h	18e5;
23415	:douta	=	16'h	18c4;
23416	:douta	=	16'h	2106;
23417	:douta	=	16'h	18e5;
23418	:douta	=	16'h	18e5;
23419	:douta	=	16'h	0883;
23420	:douta	=	16'h	0863;
23421	:douta	=	16'h	73f2;
23422	:douta	=	16'h	8453;
23423	:douta	=	16'h	9492;
23424	:douta	=	16'h	a4b2;
23425	:douta	=	16'h	acf2;
23426	:douta	=	16'h	7c0f;
23427	:douta	=	16'h	634d;
23428	:douta	=	16'h	39e8;
23429	:douta	=	16'h	42ae;
23430	:douta	=	16'h	8d18;
23431	:douta	=	16'h	8d18;
23432	:douta	=	16'h	84d7;
23433	:douta	=	16'h	7cb7;
23434	:douta	=	16'h	8d38;
23435	:douta	=	16'h	9579;
23436	:douta	=	16'h	8d18;
23437	:douta	=	16'h	8d38;
23438	:douta	=	16'h	8d38;
23439	:douta	=	16'h	9579;
23440	:douta	=	16'h	9579;
23441	:douta	=	16'h	84f7;
23442	:douta	=	16'h	84b6;
23443	:douta	=	16'h	8d18;
23444	:douta	=	16'h	8d39;
23445	:douta	=	16'h	7cb6;
23446	:douta	=	16'h	6c35;
23447	:douta	=	16'h	84d7;
23448	:douta	=	16'h	8d18;
23449	:douta	=	16'h	84f8;
23450	:douta	=	16'h	8518;
23451	:douta	=	16'h	7c96;
23452	:douta	=	16'h	84f8;
23453	:douta	=	16'h	84d8;
23454	:douta	=	16'h	7435;
23455	:douta	=	16'h	5352;
23456	:douta	=	16'h	7496;
23457	:douta	=	16'h	8d39;
23458	:douta	=	16'h	84f8;
23459	:douta	=	16'h	9dbb;
23460	:douta	=	16'h	8d59;
23461	:douta	=	16'h	7496;
23462	:douta	=	16'h	84f8;
23463	:douta	=	16'h	8518;
23464	:douta	=	16'h	959a;
23465	:douta	=	16'h	8d5a;
23466	:douta	=	16'h	84f8;
23467	:douta	=	16'h	8539;
23468	:douta	=	16'h	8d5a;
23469	:douta	=	16'h	8539;
23470	:douta	=	16'h	8d59;
23471	:douta	=	16'h	7cf8;
23472	:douta	=	16'h	8518;
23473	:douta	=	16'h	84d8;
23474	:douta	=	16'h	7cb7;
23475	:douta	=	16'h	8518;
23476	:douta	=	16'h	8c52;
23477	:douta	=	16'h	7b2a;
23478	:douta	=	16'h	528c;
23479	:douta	=	16'h	18a2;
23480	:douta	=	16'h	31c9;
23481	:douta	=	16'h	8d7a;
23482	:douta	=	16'h	8d59;
23483	:douta	=	16'h	8538;
23484	:douta	=	16'h	9ddb;
23485	:douta	=	16'h	95ba;
23486	:douta	=	16'h	8539;
23487	:douta	=	16'h	8518;
23488	:douta	=	16'h	7cd8;
23489	:douta	=	16'h	8d5a;
23490	:douta	=	16'h	959b;
23491	:douta	=	16'h	9ddb;
23492	:douta	=	16'h	959a;
23493	:douta	=	16'h	8539;
23494	:douta	=	16'h	9ddb;
23495	:douta	=	16'h	95ba;
23496	:douta	=	16'h	a5db;
23497	:douta	=	16'h	ae1c;
23498	:douta	=	16'h	8519;
23499	:douta	=	16'h	8d9a;
23500	:douta	=	16'h	8d7a;
23501	:douta	=	16'h	8d59;
23502	:douta	=	16'h	8d59;
23503	:douta	=	16'h	a5db;
23504	:douta	=	16'h	a5fb;
23505	:douta	=	16'h	9dda;
23506	:douta	=	16'h	8d5a;
23507	:douta	=	16'h	957a;
23508	:douta	=	16'h	9d9b;
23509	:douta	=	16'h	8d5a;
23510	:douta	=	16'h	8519;
23511	:douta	=	16'h	7cd9;
23512	:douta	=	16'h	8d3a;
23513	:douta	=	16'h	8d3a;
23514	:douta	=	16'h	84f9;
23515	:douta	=	16'h	7497;
23516	:douta	=	16'h	7cb8;
23517	:douta	=	16'h	7cb8;
23518	:douta	=	16'h	853a;
23519	:douta	=	16'h	957b;
23520	:douta	=	16'h	95bb;
23521	:douta	=	16'h	8d5a;
23522	:douta	=	16'h	851a;
23523	:douta	=	16'h	84f9;
23524	:douta	=	16'h	62cb;
23525	:douta	=	16'h	4964;
23526	:douta	=	16'h	2903;
23527	:douta	=	16'h	10a2;
23528	:douta	=	16'h	0020;
23529	:douta	=	16'h	5bb4;
23530	:douta	=	16'h	8d39;
23531	:douta	=	16'h	4060;
23532	:douta	=	16'h	29ec;
23533	:douta	=	16'h	4b73;
23534	:douta	=	16'h	5bf5;
23535	:douta	=	16'h	84f9;
23536	:douta	=	16'h	7cd7;
23537	:douta	=	16'h	a61c;
23538	:douta	=	16'h	6c56;
23539	:douta	=	16'h	42f1;
23540	:douta	=	16'h	3af1;
23541	:douta	=	16'h	6288;
23542	:douta	=	16'h	0800;
23543	:douta	=	16'h	8d7a;
23544	:douta	=	16'h	9dba;
23545	:douta	=	16'h	955a;
23546	:douta	=	16'h	7c76;
23547	:douta	=	16'h	8497;
23548	:douta	=	16'h	6436;
23549	:douta	=	16'h	74b8;
23550	:douta	=	16'h	6c15;
23551	:douta	=	16'h	0020;
23552	:douta	=	16'h	3966;
23553	:douta	=	16'h	3165;
23554	:douta	=	16'h	3165;
23555	:douta	=	16'h	1063;
23556	:douta	=	16'h	4333;
23557	:douta	=	16'h	3b95;
23558	:douta	=	16'h	2a2e;
23559	:douta	=	16'h	3270;
23560	:douta	=	16'h	2a8f;
23561	:douta	=	16'h	3b12;
23562	:douta	=	16'h	4332;
23563	:douta	=	16'h	6c36;
23564	:douta	=	16'h	7456;
23565	:douta	=	16'h	7c97;
23566	:douta	=	16'h	7456;
23567	:douta	=	16'h	6bb3;
23568	:douta	=	16'h	7c55;
23569	:douta	=	16'h	8cb6;
23570	:douta	=	16'h	7413;
23571	:douta	=	16'h	9c52;
23572	:douta	=	16'h	ddb0;
23573	:douta	=	16'h	e613;
23574	:douta	=	16'h	e654;
23575	:douta	=	16'h	ee96;
23576	:douta	=	16'h	ee95;
23577	:douta	=	16'h	ee75;
23578	:douta	=	16'h	de33;
23579	:douta	=	16'h	ddf2;
23580	:douta	=	16'h	cd6f;
23581	:douta	=	16'h	bced;
23582	:douta	=	16'h	bcee;
23583	:douta	=	16'h	7b28;
23584	:douta	=	16'h	72c7;
23585	:douta	=	16'h	ac8c;
23586	:douta	=	16'h	bcee;
23587	:douta	=	16'h	bcef;
23588	:douta	=	16'h	d612;
23589	:douta	=	16'h	de33;
23590	:douta	=	16'h	ddf3;
23591	:douta	=	16'h	de34;
23592	:douta	=	16'h	cd91;
23593	:douta	=	16'h	ee95;
23594	:douta	=	16'h	eed7;
23595	:douta	=	16'h	ddf3;
23596	:douta	=	16'h	ee95;
23597	:douta	=	16'h	f6f8;
23598	:douta	=	16'h	e675;
23599	:douta	=	16'h	eeb5;
23600	:douta	=	16'h	e654;
23601	:douta	=	16'h	ddf3;
23602	:douta	=	16'h	e613;
23603	:douta	=	16'h	d5d1;
23604	:douta	=	16'h	d591;
23605	:douta	=	16'h	bcef;
23606	:douta	=	16'h	a40f;
23607	:douta	=	16'h	940e;
23608	:douta	=	16'h	7b90;
23609	:douta	=	16'h	734f;
23610	:douta	=	16'h	6b0c;
23611	:douta	=	16'h	6b2c;
23612	:douta	=	16'h	6b0c;
23613	:douta	=	16'h	62ab;
23614	:douta	=	16'h	49e9;
23615	:douta	=	16'h	8306;
23616	:douta	=	16'h	b44b;
23617	:douta	=	16'h	b46b;
23618	:douta	=	16'h	c4ed;
23619	:douta	=	16'h	d54f;
23620	:douta	=	16'h	ddf2;
23621	:douta	=	16'h	e634;
23622	:douta	=	16'h	e654;
23623	:douta	=	16'h	e654;
23624	:douta	=	16'h	ee95;
23625	:douta	=	16'h	e613;
23626	:douta	=	16'h	e654;
23627	:douta	=	16'h	ee75;
23628	:douta	=	16'h	ee54;
23629	:douta	=	16'h	e634;
23630	:douta	=	16'h	ddf3;
23631	:douta	=	16'h	d571;
23632	:douta	=	16'h	d591;
23633	:douta	=	16'h	b4b1;
23634	:douta	=	16'h	ac91;
23635	:douta	=	16'h	9431;
23636	:douta	=	16'h	a471;
23637	:douta	=	16'h	9c51;
23638	:douta	=	16'h	8c31;
23639	:douta	=	16'h	9432;
23640	:douta	=	16'h	83f1;
23641	:douta	=	16'h	8c13;
23642	:douta	=	16'h	7c12;
23643	:douta	=	16'h	73d1;
23644	:douta	=	16'h	73b0;
23645	:douta	=	16'h	736f;
23646	:douta	=	16'h	736f;
23647	:douta	=	16'h	6b2e;
23648	:douta	=	16'h	5aee;
23649	:douta	=	16'h	4208;
23650	:douta	=	16'h	7a87;
23651	:douta	=	16'h	9368;
23652	:douta	=	16'h	d56e;
23653	:douta	=	16'h	ddd2;
23654	:douta	=	16'h	9c4f;
23655	:douta	=	16'h	4ace;
23656	:douta	=	16'h	322b;
23657	:douta	=	16'h	734f;
23658	:douta	=	16'h	4aee;
23659	:douta	=	16'h	2168;
23660	:douta	=	16'h	10e5;
23661	:douta	=	16'h	1926;
23662	:douta	=	16'h	10c5;
23663	:douta	=	16'h	2988;
23664	:douta	=	16'h	5ace;
23665	:douta	=	16'h	2126;
23666	:douta	=	16'h	0062;
23667	:douta	=	16'h	18e5;
23668	:douta	=	16'h	18e5;
23669	:douta	=	16'h	1926;
23670	:douta	=	16'h	18e5;
23671	:douta	=	16'h	18e5;
23672	:douta	=	16'h	10e4;
23673	:douta	=	16'h	10c5;
23674	:douta	=	16'h	10c4;
23675	:douta	=	16'h	1905;
23676	:douta	=	16'h	0022;
23677	:douta	=	16'h	7bf3;
23678	:douta	=	16'h	4b31;
23679	:douta	=	16'h	5b70;
23680	:douta	=	16'h	4a6c;
23681	:douta	=	16'h	a4b1;
23682	:douta	=	16'h	4a6a;
23683	:douta	=	16'h	8c70;
23684	:douta	=	16'h	7b8e;
23685	:douta	=	16'h	4249;
23686	:douta	=	16'h	2189;
23687	:douta	=	16'h	a61c;
23688	:douta	=	16'h	8d18;
23689	:douta	=	16'h	9539;
23690	:douta	=	16'h	8518;
23691	:douta	=	16'h	84d7;
23692	:douta	=	16'h	8d39;
23693	:douta	=	16'h	8d58;
23694	:douta	=	16'h	8d38;
23695	:douta	=	16'h	9579;
23696	:douta	=	16'h	8d38;
23697	:douta	=	16'h	8d17;
23698	:douta	=	16'h	8cd7;
23699	:douta	=	16'h	8496;
23700	:douta	=	16'h	84f7;
23701	:douta	=	16'h	8d38;
23702	:douta	=	16'h	8d18;
23703	:douta	=	16'h	7476;
23704	:douta	=	16'h	7c96;
23705	:douta	=	16'h	7cb7;
23706	:douta	=	16'h	84d7;
23707	:douta	=	16'h	84f8;
23708	:douta	=	16'h	84d7;
23709	:douta	=	16'h	8d18;
23710	:douta	=	16'h	84b7;
23711	:douta	=	16'h	7c76;
23712	:douta	=	16'h	6c35;
23713	:douta	=	16'h	63d4;
23714	:douta	=	16'h	6c35;
23715	:douta	=	16'h	84f8;
23716	:douta	=	16'h	8518;
23717	:douta	=	16'h	8d39;
23718	:douta	=	16'h	7cd7;
23719	:douta	=	16'h	7476;
23720	:douta	=	16'h	8518;
23721	:douta	=	16'h	84d8;
23722	:douta	=	16'h	84f9;
23723	:douta	=	16'h	8d39;
23724	:douta	=	16'h	8539;
23725	:douta	=	16'h	84d8;
23726	:douta	=	16'h	8539;
23727	:douta	=	16'h	8d7a;
23728	:douta	=	16'h	8539;
23729	:douta	=	16'h	8d59;
23730	:douta	=	16'h	7cf8;
23731	:douta	=	16'h	8518;
23732	:douta	=	16'h	8c73;
23733	:douta	=	16'h	832b;
23734	:douta	=	16'h	52ad;
23735	:douta	=	16'h	1861;
23736	:douta	=	16'h	39e9;
23737	:douta	=	16'h	8d7a;
23738	:douta	=	16'h	8539;
23739	:douta	=	16'h	8d5a;
23740	:douta	=	16'h	8519;
23741	:douta	=	16'h	8518;
23742	:douta	=	16'h	9dbb;
23743	:douta	=	16'h	959a;
23744	:douta	=	16'h	84f9;
23745	:douta	=	16'h	8519;
23746	:douta	=	16'h	8d59;
23747	:douta	=	16'h	959a;
23748	:douta	=	16'h	8d7a;
23749	:douta	=	16'h	9dbb;
23750	:douta	=	16'h	8d59;
23751	:douta	=	16'h	8d7a;
23752	:douta	=	16'h	9d9a;
23753	:douta	=	16'h	ae1c;
23754	:douta	=	16'h	7cd9;
23755	:douta	=	16'h	9ddb;
23756	:douta	=	16'h	959a;
23757	:douta	=	16'h	959a;
23758	:douta	=	16'h	959a;
23759	:douta	=	16'h	9ddb;
23760	:douta	=	16'h	957a;
23761	:douta	=	16'h	9ddb;
23762	:douta	=	16'h	95bb;
23763	:douta	=	16'h	957a;
23764	:douta	=	16'h	9d9a;
23765	:douta	=	16'h	957a;
23766	:douta	=	16'h	959a;
23767	:douta	=	16'h	8d59;
23768	:douta	=	16'h	8519;
23769	:douta	=	16'h	959b;
23770	:douta	=	16'h	959a;
23771	:douta	=	16'h	95bb;
23772	:douta	=	16'h	8519;
23773	:douta	=	16'h	84f9;
23774	:douta	=	16'h	6c37;
23775	:douta	=	16'h	957b;
23776	:douta	=	16'h	8d7b;
23777	:douta	=	16'h	7d3b;
23778	:douta	=	16'h	74b8;
23779	:douta	=	16'h	6b2e;
23780	:douta	=	16'h	6244;
23781	:douta	=	16'h	6246;
23782	:douta	=	16'h	3124;
23783	:douta	=	16'h	18c3;
23784	:douta	=	16'h	0882;
23785	:douta	=	16'h	29cb;
23786	:douta	=	16'h	6c57;
23787	:douta	=	16'h	942e;
23788	:douta	=	16'h	3880;
23789	:douta	=	16'h	74fa;
23790	:douta	=	16'h	6416;
23791	:douta	=	16'h	4311;
23792	:douta	=	16'h	5bb4;
23793	:douta	=	16'h	6c35;
23794	:douta	=	16'h	ae3d;
23795	:douta	=	16'h	6c15;
23796	:douta	=	16'h	95dd;
23797	:douta	=	16'h	1800;
23798	:douta	=	16'h	29a9;
23799	:douta	=	16'h	4b32;
23800	:douta	=	16'h	b65c;
23801	:douta	=	16'h	8d39;
23802	:douta	=	16'h	9dbb;
23803	:douta	=	16'h	9dbb;
23804	:douta	=	16'h	6436;
23805	:douta	=	16'h	7c77;
23806	:douta	=	16'h	6415;
23807	:douta	=	16'h	0000;
23808	:douta	=	16'h	3966;
23809	:douta	=	16'h	3966;
23810	:douta	=	16'h	3145;
23811	:douta	=	16'h	20c3;
23812	:douta	=	16'h	29ec;
23813	:douta	=	16'h	32d2;
23814	:douta	=	16'h	3290;
23815	:douta	=	16'h	3290;
23816	:douta	=	16'h	3b12;
23817	:douta	=	16'h	5bf6;
23818	:douta	=	16'h	53b4;
23819	:douta	=	16'h	4b32;
23820	:douta	=	16'h	5b93;
23821	:douta	=	16'h	3a8f;
23822	:douta	=	16'h	6c36;
23823	:douta	=	16'h	7414;
23824	:douta	=	16'h	7435;
23825	:douta	=	16'h	8cf7;
23826	:douta	=	16'h	7c34;
23827	:douta	=	16'h	a578;
23828	:douta	=	16'h	bd55;
23829	:douta	=	16'h	de34;
23830	:douta	=	16'h	e695;
23831	:douta	=	16'h	ee96;
23832	:douta	=	16'h	d5d2;
23833	:douta	=	16'h	ddf3;
23834	:douta	=	16'h	ddf3;
23835	:douta	=	16'h	d591;
23836	:douta	=	16'h	bcef;
23837	:douta	=	16'h	ac6c;
23838	:douta	=	16'h	7ae8;
23839	:douta	=	16'h	b48d;
23840	:douta	=	16'h	b4ee;
23841	:douta	=	16'h	b4ad;
23842	:douta	=	16'h	c54f;
23843	:douta	=	16'h	c530;
23844	:douta	=	16'h	de34;
23845	:douta	=	16'h	e654;
23846	:douta	=	16'h	de14;
23847	:douta	=	16'h	e675;
23848	:douta	=	16'h	e655;
23849	:douta	=	16'h	e634;
23850	:douta	=	16'h	eeb7;
23851	:douta	=	16'h	eeb7;
23852	:douta	=	16'h	cd2e;
23853	:douta	=	16'h	d571;
23854	:douta	=	16'h	f6f7;
23855	:douta	=	16'h	ee95;
23856	:douta	=	16'h	e633;
23857	:douta	=	16'h	d5b1;
23858	:douta	=	16'h	d591;
23859	:douta	=	16'h	cd50;
23860	:douta	=	16'h	bccf;
23861	:douta	=	16'h	a46f;
23862	:douta	=	16'h	83cf;
23863	:douta	=	16'h	7b6f;
23864	:douta	=	16'h	734e;
23865	:douta	=	16'h	730e;
23866	:douta	=	16'h	62cb;
23867	:douta	=	16'h	62ab;
23868	:douta	=	16'h	524a;
23869	:douta	=	16'h	51c4;
23870	:douta	=	16'h	9b48;
23871	:douta	=	16'h	ac0b;
23872	:douta	=	16'h	bc8b;
23873	:douta	=	16'h	c50d;
23874	:douta	=	16'h	e5f2;
23875	:douta	=	16'h	e634;
23876	:douta	=	16'h	e674;
23877	:douta	=	16'h	e654;
23878	:douta	=	16'h	e674;
23879	:douta	=	16'h	ee95;
23880	:douta	=	16'h	ee75;
23881	:douta	=	16'h	e655;
23882	:douta	=	16'h	ee95;
23883	:douta	=	16'h	e654;
23884	:douta	=	16'h	ddf3;
23885	:douta	=	16'h	ddd2;
23886	:douta	=	16'h	d5b2;
23887	:douta	=	16'h	bcd1;
23888	:douta	=	16'h	bcf1;
23889	:douta	=	16'h	acb2;
23890	:douta	=	16'h	acb1;
23891	:douta	=	16'h	9c71;
23892	:douta	=	16'h	9c92;
23893	:douta	=	16'h	9472;
23894	:douta	=	16'h	8c32;
23895	:douta	=	16'h	8412;
23896	:douta	=	16'h	7bd1;
23897	:douta	=	16'h	7bd1;
23898	:douta	=	16'h	7370;
23899	:douta	=	16'h	734e;
23900	:douta	=	16'h	6aed;
23901	:douta	=	16'h	62ed;
23902	:douta	=	16'h	6aed;
23903	:douta	=	16'h	49e8;
23904	:douta	=	16'h	9307;
23905	:douta	=	16'h	b42b;
23906	:douta	=	16'h	d50e;
23907	:douta	=	16'h	e633;
23908	:douta	=	16'h	eeb6;
23909	:douta	=	16'h	cd71;
23910	:douta	=	16'h	ac90;
23911	:douta	=	16'h	6b70;
23912	:douta	=	16'h	52ef;
23913	:douta	=	16'h	83d0;
23914	:douta	=	16'h	73b1;
23915	:douta	=	16'h	31eb;
23916	:douta	=	16'h	29a9;
23917	:douta	=	16'h	39ea;
23918	:douta	=	16'h	2988;
23919	:douta	=	16'h	18e5;
23920	:douta	=	16'h	18e5;
23921	:douta	=	16'h	1927;
23922	:douta	=	16'h	5b2f;
23923	:douta	=	16'h	10e6;
23924	:douta	=	16'h	18e5;
23925	:douta	=	16'h	18e5;
23926	:douta	=	16'h	18e5;
23927	:douta	=	16'h	1905;
23928	:douta	=	16'h	18e5;
23929	:douta	=	16'h	1905;
23930	:douta	=	16'h	18e5;
23931	:douta	=	16'h	10e4;
23932	:douta	=	16'h	10c5;
23933	:douta	=	16'h	08a4;
23934	:douta	=	16'h	2946;
23935	:douta	=	16'h	6bb1;
23936	:douta	=	16'h	6c13;
23937	:douta	=	16'h	6c33;
23938	:douta	=	16'h	83ee;
23939	:douta	=	16'h	8c30;
23940	:douta	=	16'h	ad33;
23941	:douta	=	16'h	a512;
23942	:douta	=	16'h	6b6c;
23943	:douta	=	16'h	2967;
23944	:douta	=	16'h	5b92;
23945	:douta	=	16'h	9dfc;
23946	:douta	=	16'h	9579;
23947	:douta	=	16'h	8d18;
23948	:douta	=	16'h	84f8;
23949	:douta	=	16'h	9559;
23950	:douta	=	16'h	84f8;
23951	:douta	=	16'h	84f8;
23952	:douta	=	16'h	8d18;
23953	:douta	=	16'h	8d38;
23954	:douta	=	16'h	84b6;
23955	:douta	=	16'h	9538;
23956	:douta	=	16'h	84d7;
23957	:douta	=	16'h	84d7;
23958	:douta	=	16'h	84d7;
23959	:douta	=	16'h	7cb7;
23960	:douta	=	16'h	8d39;
23961	:douta	=	16'h	8d39;
23962	:douta	=	16'h	9559;
23963	:douta	=	16'h	8d59;
23964	:douta	=	16'h	8d18;
23965	:douta	=	16'h	84f8;
23966	:douta	=	16'h	84f8;
23967	:douta	=	16'h	84f8;
23968	:douta	=	16'h	7476;
23969	:douta	=	16'h	8cd8;
23970	:douta	=	16'h	8d18;
23971	:douta	=	16'h	6c15;
23972	:douta	=	16'h	6c35;
23973	:douta	=	16'h	7c96;
23974	:douta	=	16'h	63d4;
23975	:douta	=	16'h	8d19;
23976	:douta	=	16'h	7c97;
23977	:douta	=	16'h	7cd7;
23978	:douta	=	16'h	8539;
23979	:douta	=	16'h	7cf8;
23980	:douta	=	16'h	8519;
23981	:douta	=	16'h	8d7a;
23982	:douta	=	16'h	959b;
23983	:douta	=	16'h	8539;
23984	:douta	=	16'h	84f8;
23985	:douta	=	16'h	8d3a;
23986	:douta	=	16'h	8539;
23987	:douta	=	16'h	8d5a;
23988	:douta	=	16'h	8c53;
23989	:douta	=	16'h	6246;
23990	:douta	=	16'h	5a6b;
23991	:douta	=	16'h	0820;
23992	:douta	=	16'h	4a6c;
23993	:douta	=	16'h	8519;
23994	:douta	=	16'h	8d59;
23995	:douta	=	16'h	9559;
23996	:douta	=	16'h	8d59;
23997	:douta	=	16'h	955a;
23998	:douta	=	16'h	8d39;
23999	:douta	=	16'h	8d59;
24000	:douta	=	16'h	8d39;
24001	:douta	=	16'h	957a;
24002	:douta	=	16'h	959a;
24003	:douta	=	16'h	84d8;
24004	:douta	=	16'h	8d59;
24005	:douta	=	16'h	8d39;
24006	:douta	=	16'h	8519;
24007	:douta	=	16'h	84f9;
24008	:douta	=	16'h	9ddb;
24009	:douta	=	16'h	9dbb;
24010	:douta	=	16'h	a5db;
24011	:douta	=	16'h	8d7a;
24012	:douta	=	16'h	8d5a;
24013	:douta	=	16'h	8d7a;
24014	:douta	=	16'h	8d7a;
24015	:douta	=	16'h	9dbb;
24016	:douta	=	16'h	959a;
24017	:douta	=	16'h	8d7a;
24018	:douta	=	16'h	7d18;
24019	:douta	=	16'h	8d7a;
24020	:douta	=	16'h	9d9b;
24021	:douta	=	16'h	9dba;
24022	:douta	=	16'h	8d7a;
24023	:douta	=	16'h	9ddb;
24024	:douta	=	16'h	9dbb;
24025	:douta	=	16'h	84f9;
24026	:douta	=	16'h	957b;
24027	:douta	=	16'h	959a;
24028	:douta	=	16'h	8d5a;
24029	:douta	=	16'h	959b;
24030	:douta	=	16'h	ae5e;
24031	:douta	=	16'h	a61d;
24032	:douta	=	16'h	9d38;
24033	:douta	=	16'h	5aad;
24034	:douta	=	16'h	424d;
24035	:douta	=	16'h	8ddf;
24036	:douta	=	16'h	6203;
24037	:douta	=	16'h	7ac8;
24038	:douta	=	16'h	4985;
24039	:douta	=	16'h	3123;
24040	:douta	=	16'h	0882;
24041	:douta	=	16'h	0000;
24042	:douta	=	16'h	3a8d;
24043	:douta	=	16'h	4374;
24044	:douta	=	16'h	6477;
24045	:douta	=	16'h	2840;
24046	:douta	=	16'h	4353;
24047	:douta	=	16'h	5392;
24048	:douta	=	16'h	9579;
24049	:douta	=	16'h	959a;
24050	:douta	=	16'h	7cd7;
24051	:douta	=	16'h	7498;
24052	:douta	=	16'h	7436;
24053	:douta	=	16'h	18a2;
24054	:douta	=	16'h	5c16;
24055	:douta	=	16'h	a5db;
24056	:douta	=	16'h	6c56;
24057	:douta	=	16'h	9d9b;
24058	:douta	=	16'h	7cb8;
24059	:douta	=	16'h	6c77;
24060	:douta	=	16'h	7476;
24061	:douta	=	16'h	84f8;
24062	:douta	=	16'h	a5db;
24063	:douta	=	16'h	0000;
24064	:douta	=	16'h	3966;
24065	:douta	=	16'h	3166;
24066	:douta	=	16'h	3146;
24067	:douta	=	16'h	18c4;
24068	:douta	=	16'h	29eb;
24069	:douta	=	16'h	4354;
24070	:douta	=	16'h	220d;
24071	:douta	=	16'h	4312;
24072	:douta	=	16'h	3290;
24073	:douta	=	16'h	32b0;
24074	:douta	=	16'h	4332;
24075	:douta	=	16'h	6416;
24076	:douta	=	16'h	6c36;
24077	:douta	=	16'h	5353;
24078	:douta	=	16'h	7cd9;
24079	:douta	=	16'h	63b3;
24080	:douta	=	16'h	4acf;
24081	:douta	=	16'h	6bd3;
24082	:douta	=	16'h	7413;
24083	:douta	=	16'h	73d1;
24084	:douta	=	16'h	8c75;
24085	:douta	=	16'h	e632;
24086	:douta	=	16'h	ee96;
24087	:douta	=	16'h	ee75;
24088	:douta	=	16'h	de13;
24089	:douta	=	16'h	cd70;
24090	:douta	=	16'h	d5d1;
24091	:douta	=	16'h	cd71;
24092	:douta	=	16'h	b4ad;
24093	:douta	=	16'h	8329;
24094	:douta	=	16'h	7b07;
24095	:douta	=	16'h	bcee;
24096	:douta	=	16'h	bcee;
24097	:douta	=	16'h	bd0f;
24098	:douta	=	16'h	c52f;
24099	:douta	=	16'h	cd71;
24100	:douta	=	16'h	e655;
24101	:douta	=	16'h	e676;
24102	:douta	=	16'h	de13;
24103	:douta	=	16'h	e696;
24104	:douta	=	16'h	e696;
24105	:douta	=	16'h	e654;
24106	:douta	=	16'h	e675;
24107	:douta	=	16'h	ee96;
24108	:douta	=	16'h	ddd2;
24109	:douta	=	16'h	c4ee;
24110	:douta	=	16'h	ee95;
24111	:douta	=	16'h	eed6;
24112	:douta	=	16'h	ddf2;
24113	:douta	=	16'h	d591;
24114	:douta	=	16'h	cd70;
24115	:douta	=	16'h	bcf0;
24116	:douta	=	16'h	ac8f;
24117	:douta	=	16'h	9410;
24118	:douta	=	16'h	8bf0;
24119	:douta	=	16'h	7b8f;
24120	:douta	=	16'h	6b2e;
24121	:douta	=	16'h	6aec;
24122	:douta	=	16'h	6b0c;
24123	:douta	=	16'h	5a6a;
24124	:douta	=	16'h	3125;
24125	:douta	=	16'h	a389;
24126	:douta	=	16'h	abea;
24127	:douta	=	16'h	bc8c;
24128	:douta	=	16'h	cd2d;
24129	:douta	=	16'h	d58f;
24130	:douta	=	16'h	e654;
24131	:douta	=	16'h	ee95;
24132	:douta	=	16'h	e675;
24133	:douta	=	16'h	ee95;
24134	:douta	=	16'h	e674;
24135	:douta	=	16'h	ee75;
24136	:douta	=	16'h	ee95;
24137	:douta	=	16'h	e654;
24138	:douta	=	16'h	e633;
24139	:douta	=	16'h	ee75;
24140	:douta	=	16'h	d5b3;
24141	:douta	=	16'h	cd72;
24142	:douta	=	16'h	c552;
24143	:douta	=	16'h	bd12;
24144	:douta	=	16'h	bd11;
24145	:douta	=	16'h	acb3;
24146	:douta	=	16'h	a492;
24147	:douta	=	16'h	9c93;
24148	:douta	=	16'h	9472;
24149	:douta	=	16'h	9452;
24150	:douta	=	16'h	8432;
24151	:douta	=	16'h	8432;
24152	:douta	=	16'h	7391;
24153	:douta	=	16'h	6b4f;
24154	:douta	=	16'h	6b2e;
24155	:douta	=	16'h	630e;
24156	:douta	=	16'h	62ec;
24157	:douta	=	16'h	6aed;
24158	:douta	=	16'h	5a6a;
24159	:douta	=	16'h	6226;
24160	:douta	=	16'h	b46b;
24161	:douta	=	16'h	bc8d;
24162	:douta	=	16'h	ddd0;
24163	:douta	=	16'h	e633;
24164	:douta	=	16'h	e634;
24165	:douta	=	16'h	d591;
24166	:douta	=	16'h	bcf0;
24167	:douta	=	16'h	7391;
24168	:douta	=	16'h	6330;
24169	:douta	=	16'h	9431;
24170	:douta	=	16'h	8412;
24171	:douta	=	16'h	3a2c;
24172	:douta	=	16'h	31ca;
24173	:douta	=	16'h	3a0a;
24174	:douta	=	16'h	3a2c;
24175	:douta	=	16'h	2989;
24176	:douta	=	16'h	2127;
24177	:douta	=	16'h	1084;
24178	:douta	=	16'h	0863;
24179	:douta	=	16'h	5b51;
24180	:douta	=	16'h	0842;
24181	:douta	=	16'h	18e5;
24182	:douta	=	16'h	10c5;
24183	:douta	=	16'h	10c4;
24184	:douta	=	16'h	18e5;
24185	:douta	=	16'h	1906;
24186	:douta	=	16'h	18e4;
24187	:douta	=	16'h	10a4;
24188	:douta	=	16'h	18e5;
24189	:douta	=	16'h	1905;
24190	:douta	=	16'h	0001;
24191	:douta	=	16'h	0862;
24192	:douta	=	16'h	7c74;
24193	:douta	=	16'h	7475;
24194	:douta	=	16'h	42cf;
24195	:douta	=	16'h	424a;
24196	:douta	=	16'h	52ac;
24197	:douta	=	16'h	7bef;
24198	:douta	=	16'h	2988;
24199	:douta	=	16'h	7bae;
24200	:douta	=	16'h	29ca;
24201	:douta	=	16'h	5b50;
24202	:douta	=	16'h	ae3d;
24203	:douta	=	16'h	ae3d;
24204	:douta	=	16'h	7cf8;
24205	:douta	=	16'h	8d18;
24206	:douta	=	16'h	9579;
24207	:douta	=	16'h	8d59;
24208	:douta	=	16'h	8d38;
24209	:douta	=	16'h	84d6;
24210	:douta	=	16'h	8d18;
24211	:douta	=	16'h	9538;
24212	:douta	=	16'h	84f7;
24213	:douta	=	16'h	84d7;
24214	:douta	=	16'h	a5fb;
24215	:douta	=	16'h	7476;
24216	:douta	=	16'h	7cb7;
24217	:douta	=	16'h	84f8;
24218	:douta	=	16'h	84f8;
24219	:douta	=	16'h	959a;
24220	:douta	=	16'h	7cb7;
24221	:douta	=	16'h	84d7;
24222	:douta	=	16'h	9579;
24223	:douta	=	16'h	a59a;
24224	:douta	=	16'h	7c96;
24225	:douta	=	16'h	84b7;
24226	:douta	=	16'h	84d7;
24227	:douta	=	16'h	84d7;
24228	:douta	=	16'h	7435;
24229	:douta	=	16'h	7c96;
24230	:douta	=	16'h	7c96;
24231	:douta	=	16'h	7476;
24232	:douta	=	16'h	6c15;
24233	:douta	=	16'h	63b3;
24234	:douta	=	16'h	84d8;
24235	:douta	=	16'h	8519;
24236	:douta	=	16'h	8d7b;
24237	:douta	=	16'h	7cb8;
24238	:douta	=	16'h	7cb7;
24239	:douta	=	16'h	8d5a;
24240	:douta	=	16'h	8d5a;
24241	:douta	=	16'h	84f9;
24242	:douta	=	16'h	84f9;
24243	:douta	=	16'h	8d39;
24244	:douta	=	16'h	8d18;
24245	:douta	=	16'h	628a;
24246	:douta	=	16'h	5208;
24247	:douta	=	16'h	3146;
24248	:douta	=	16'h	7455;
24249	:douta	=	16'h	7cf8;
24250	:douta	=	16'h	84f8;
24251	:douta	=	16'h	8539;
24252	:douta	=	16'h	8d59;
24253	:douta	=	16'h	8519;
24254	:douta	=	16'h	957a;
24255	:douta	=	16'h	9559;
24256	:douta	=	16'h	8d39;
24257	:douta	=	16'h	8518;
24258	:douta	=	16'h	959a;
24259	:douta	=	16'h	8519;
24260	:douta	=	16'h	74b8;
24261	:douta	=	16'h	9dbb;
24262	:douta	=	16'h	8d59;
24263	:douta	=	16'h	8d5a;
24264	:douta	=	16'h	8d19;
24265	:douta	=	16'h	957a;
24266	:douta	=	16'h	a61c;
24267	:douta	=	16'h	9dba;
24268	:douta	=	16'h	9ddb;
24269	:douta	=	16'h	8d59;
24270	:douta	=	16'h	8539;
24271	:douta	=	16'h	959a;
24272	:douta	=	16'h	957a;
24273	:douta	=	16'h	8d7a;
24274	:douta	=	16'h	959a;
24275	:douta	=	16'h	957a;
24276	:douta	=	16'h	9dbb;
24277	:douta	=	16'h	8d5a;
24278	:douta	=	16'h	8d3a;
24279	:douta	=	16'h	9ddb;
24280	:douta	=	16'h	9ddb;
24281	:douta	=	16'h	959a;
24282	:douta	=	16'h	959a;
24283	:douta	=	16'h	8d5a;
24284	:douta	=	16'h	8559;
24285	:douta	=	16'h	8d3a;
24286	:douta	=	16'h	8dbc;
24287	:douta	=	16'h	ad57;
24288	:douta	=	16'h	7b6e;
24289	:douta	=	16'h	3b13;
24290	:douta	=	16'h	5417;
24291	:douta	=	16'h	6498;
24292	:douta	=	16'h	6b2c;
24293	:douta	=	16'h	7a65;
24294	:douta	=	16'h	51e4;
24295	:douta	=	16'h	4144;
24296	:douta	=	16'h	1083;
24297	:douta	=	16'h	1061;
24298	:douta	=	16'h	0000;
24299	:douta	=	16'h	7cda;
24300	:douta	=	16'h	74fa;
24301	:douta	=	16'h	8308;
24302	:douta	=	16'h	4b53;
24303	:douta	=	16'h	84f8;
24304	:douta	=	16'h	6c35;
24305	:douta	=	16'h	7c97;
24306	:douta	=	16'h	8d18;
24307	:douta	=	16'h	74ba;
24308	:douta	=	16'h	7390;
24309	:douta	=	16'h	320c;
24310	:douta	=	16'h	855a;
24311	:douta	=	16'h	6415;
24312	:douta	=	16'h	7497;
24313	:douta	=	16'h	84b8;
24314	:douta	=	16'h	7cb8;
24315	:douta	=	16'h	7c98;
24316	:douta	=	16'h	b65d;
24317	:douta	=	16'h	74d9;
24318	:douta	=	16'h	4aef;
24319	:douta	=	16'h	0821;
24320	:douta	=	16'h	3985;
24321	:douta	=	16'h	3966;
24322	:douta	=	16'h	3145;
24323	:douta	=	16'h	3146;
24324	:douta	=	16'h	29a9;
24325	:douta	=	16'h	3af1;
24326	:douta	=	16'h	21ed;
24327	:douta	=	16'h	32b0;
24328	:douta	=	16'h	32d1;
24329	:douta	=	16'h	5394;
24330	:douta	=	16'h	63f6;
24331	:douta	=	16'h	3aaf;
24332	:douta	=	16'h	4af0;
24333	:douta	=	16'h	6c56;
24334	:douta	=	16'h	7477;
24335	:douta	=	16'h	42af;
24336	:douta	=	16'h	5330;
24337	:douta	=	16'h	7414;
24338	:douta	=	16'h	6bd3;
24339	:douta	=	16'h	a557;
24340	:douta	=	16'h	ad98;
24341	:douta	=	16'h	d593;
24342	:douta	=	16'h	ee73;
24343	:douta	=	16'h	ee75;
24344	:douta	=	16'h	e654;
24345	:douta	=	16'h	d5d2;
24346	:douta	=	16'h	c550;
24347	:douta	=	16'h	c50e;
24348	:douta	=	16'h	8b6a;
24349	:douta	=	16'h	ac6c;
24350	:douta	=	16'h	bcee;
24351	:douta	=	16'h	bd0f;
24352	:douta	=	16'h	bd0e;
24353	:douta	=	16'h	d5d2;
24354	:douta	=	16'h	cd90;
24355	:douta	=	16'h	e634;
24356	:douta	=	16'h	de54;
24357	:douta	=	16'h	ee96;
24358	:douta	=	16'h	de14;
24359	:douta	=	16'h	eeb7;
24360	:douta	=	16'h	e655;
24361	:douta	=	16'h	f6d8;
24362	:douta	=	16'h	eeb6;
24363	:douta	=	16'h	ee75;
24364	:douta	=	16'h	e635;
24365	:douta	=	16'h	e634;
24366	:douta	=	16'h	ac2d;
24367	:douta	=	16'h	ac2d;
24368	:douta	=	16'h	ee94;
24369	:douta	=	16'h	c550;
24370	:douta	=	16'h	bcf0;
24371	:douta	=	16'h	ac70;
24372	:douta	=	16'h	9c50;
24373	:douta	=	16'h	8bf0;
24374	:douta	=	16'h	7b8f;
24375	:douta	=	16'h	6b4d;
24376	:douta	=	16'h	62cc;
24377	:douta	=	16'h	628b;
24378	:douta	=	16'h	4a09;
24379	:douta	=	16'h	6206;
24380	:douta	=	16'h	c4ab;
24381	:douta	=	16'h	ac2b;
24382	:douta	=	16'h	bc8b;
24383	:douta	=	16'h	cd2e;
24384	:douta	=	16'h	e633;
24385	:douta	=	16'h	e634;
24386	:douta	=	16'h	ee75;
24387	:douta	=	16'h	e654;
24388	:douta	=	16'h	eeb6;
24389	:douta	=	16'h	ee95;
24390	:douta	=	16'h	ee74;
24391	:douta	=	16'h	de13;
24392	:douta	=	16'h	ddf3;
24393	:douta	=	16'h	d5b2;
24394	:douta	=	16'h	bcf1;
24395	:douta	=	16'h	cd52;
24396	:douta	=	16'h	cd72;
24397	:douta	=	16'h	bd12;
24398	:douta	=	16'h	acd2;
24399	:douta	=	16'h	b4f2;
24400	:douta	=	16'h	a4b3;
24401	:douta	=	16'h	9cb3;
24402	:douta	=	16'h	9c94;
24403	:douta	=	16'h	9473;
24404	:douta	=	16'h	8433;
24405	:douta	=	16'h	8433;
24406	:douta	=	16'h	73b1;
24407	:douta	=	16'h	736f;
24408	:douta	=	16'h	6b2f;
24409	:douta	=	16'h	630e;
24410	:douta	=	16'h	6b0d;
24411	:douta	=	16'h	6b0e;
24412	:douta	=	16'h	62ad;
24413	:douta	=	16'h	6227;
24414	:douta	=	16'h	8b28;
24415	:douta	=	16'h	c46c;
24416	:douta	=	16'h	cd6e;
24417	:douta	=	16'h	d590;
24418	:douta	=	16'h	de11;
24419	:douta	=	16'h	de12;
24420	:douta	=	16'h	e612;
24421	:douta	=	16'h	ddf2;
24422	:douta	=	16'h	cd71;
24423	:douta	=	16'h	8c10;
24424	:douta	=	16'h	7bd0;
24425	:douta	=	16'h	9432;
24426	:douta	=	16'h	9474;
24427	:douta	=	16'h	5b91;
24428	:douta	=	16'h	3a6c;
24429	:douta	=	16'h	4aae;
24430	:douta	=	16'h	324c;
24431	:douta	=	16'h	324d;
24432	:douta	=	16'h	322b;
24433	:douta	=	16'h	29c9;
24434	:douta	=	16'h	1947;
24435	:douta	=	16'h	08a4;
24436	:douta	=	16'h	5b51;
24437	:douta	=	16'h	428d;
24438	:douta	=	16'h	10a4;
24439	:douta	=	16'h	18e5;
24440	:douta	=	16'h	10c5;
24441	:douta	=	16'h	10e4;
24442	:douta	=	16'h	18c5;
24443	:douta	=	16'h	10e4;
24444	:douta	=	16'h	10c5;
24445	:douta	=	16'h	1905;
24446	:douta	=	16'h	10e5;
24447	:douta	=	16'h	1906;
24448	:douta	=	16'h	0042;
24449	:douta	=	16'h	0000;
24450	:douta	=	16'h	7c54;
24451	:douta	=	16'h	31ea;
24452	:douta	=	16'h	0000;
24453	:douta	=	16'h	0885;
24454	:douta	=	16'h	52ed;
24455	:douta	=	16'h	4a6a;
24456	:douta	=	16'h	73f3;
24457	:douta	=	16'h	4209;
24458	:douta	=	16'h	41c8;
24459	:douta	=	16'h	2169;
24460	:douta	=	16'h	9d9a;
24461	:douta	=	16'h	959a;
24462	:douta	=	16'h	9d79;
24463	:douta	=	16'h	8d18;
24464	:douta	=	16'h	9559;
24465	:douta	=	16'h	8d18;
24466	:douta	=	16'h	84d6;
24467	:douta	=	16'h	7c96;
24468	:douta	=	16'h	8d18;
24469	:douta	=	16'h	84d7;
24470	:douta	=	16'h	84b7;
24471	:douta	=	16'h	84d7;
24472	:douta	=	16'h	7476;
24473	:douta	=	16'h	9579;
24474	:douta	=	16'h	9579;
24475	:douta	=	16'h	7c76;
24476	:douta	=	16'h	8d38;
24477	:douta	=	16'h	84d7;
24478	:douta	=	16'h	8d38;
24479	:douta	=	16'h	8d18;
24480	:douta	=	16'h	9579;
24481	:douta	=	16'h	8d59;
24482	:douta	=	16'h	9559;
24483	:douta	=	16'h	8d39;
24484	:douta	=	16'h	9559;
24485	:douta	=	16'h	8d39;
24486	:douta	=	16'h	84d7;
24487	:douta	=	16'h	7cb7;
24488	:douta	=	16'h	9d9a;
24489	:douta	=	16'h	8d39;
24490	:douta	=	16'h	6391;
24491	:douta	=	16'h	63b2;
24492	:douta	=	16'h	6bd2;
24493	:douta	=	16'h	7cb7;
24494	:douta	=	16'h	7cb7;
24495	:douta	=	16'h	8d7a;
24496	:douta	=	16'h	7cb8;
24497	:douta	=	16'h	8539;
24498	:douta	=	16'h	7cd8;
24499	:douta	=	16'h	8519;
24500	:douta	=	16'h	8539;
24501	:douta	=	16'h	8d5b;
24502	:douta	=	16'h	857b;
24503	:douta	=	16'h	95bc;
24504	:douta	=	16'h	7cd8;
24505	:douta	=	16'h	959a;
24506	:douta	=	16'h	95bb;
24507	:douta	=	16'h	74b8;
24508	:douta	=	16'h	84f9;
24509	:douta	=	16'h	8519;
24510	:douta	=	16'h	84d8;
24511	:douta	=	16'h	957a;
24512	:douta	=	16'h	8d59;
24513	:douta	=	16'h	957a;
24514	:douta	=	16'h	8d19;
24515	:douta	=	16'h	8d19;
24516	:douta	=	16'h	8519;
24517	:douta	=	16'h	9dbb;
24518	:douta	=	16'h	959a;
24519	:douta	=	16'h	957a;
24520	:douta	=	16'h	959a;
24521	:douta	=	16'h	8d7a;
24522	:douta	=	16'h	8d5a;
24523	:douta	=	16'h	a5db;
24524	:douta	=	16'h	957a;
24525	:douta	=	16'h	a5db;
24526	:douta	=	16'h	a5fc;
24527	:douta	=	16'h	a5db;
24528	:douta	=	16'h	9dbb;
24529	:douta	=	16'h	a5db;
24530	:douta	=	16'h	9dda;
24531	:douta	=	16'h	959a;
24532	:douta	=	16'h	959a;
24533	:douta	=	16'h	a5fb;
24534	:douta	=	16'h	b65c;
24535	:douta	=	16'h	959a;
24536	:douta	=	16'h	8d7a;
24537	:douta	=	16'h	959a;
24538	:douta	=	16'h	957a;
24539	:douta	=	16'h	a5dc;
24540	:douta	=	16'h	9dfc;
24541	:douta	=	16'h	8c95;
24542	:douta	=	16'h	5b0e;
24543	:douta	=	16'h	5c38;
24544	:douta	=	16'h	5c79;
24545	:douta	=	16'h	857c;
24546	:douta	=	16'h	5c16;
24547	:douta	=	16'h	5373;
24548	:douta	=	16'h	6cba;
24549	:douta	=	16'h	630c;
24550	:douta	=	16'h	7b08;
24551	:douta	=	16'h	6245;
24552	:douta	=	16'h	20e3;
24553	:douta	=	16'h	0842;
24554	:douta	=	16'h	0862;
24555	:douta	=	16'h	5331;
24556	:douta	=	16'h	857c;
24557	:douta	=	16'h	6458;
24558	:douta	=	16'h	61c3;
24559	:douta	=	16'h	10a5;
24560	:douta	=	16'h	8518;
24561	:douta	=	16'h	7cd7;
24562	:douta	=	16'h	7456;
24563	:douta	=	16'h	7c32;
24564	:douta	=	16'h	3040;
24565	:douta	=	16'h	7498;
24566	:douta	=	16'h	21ec;
24567	:douta	=	16'h	5352;
24568	:douta	=	16'h	63d3;
24569	:douta	=	16'h	6415;
24570	:douta	=	16'h	be5c;
24571	:douta	=	16'h	84d8;
24572	:douta	=	16'h	6c78;
24573	:douta	=	16'h	0000;
24574	:douta	=	16'h	29a8;
24575	:douta	=	16'h	4acd;
24576	:douta	=	16'h	3965;
24577	:douta	=	16'h	3966;
24578	:douta	=	16'h	3165;
24579	:douta	=	16'h	2926;
24580	:douta	=	16'h	3a4d;
24581	:douta	=	16'h	3ad1;
24582	:douta	=	16'h	324f;
24583	:douta	=	16'h	3af1;
24584	:douta	=	16'h	53d6;
24585	:douta	=	16'h	32b0;
24586	:douta	=	16'h	4b73;
24587	:douta	=	16'h	4b32;
24588	:douta	=	16'h	63f4;
24589	:douta	=	16'h	7457;
24590	:douta	=	16'h	7cb8;
24591	:douta	=	16'h	5331;
24592	:douta	=	16'h	5351;
24593	:douta	=	16'h	6bf4;
24594	:douta	=	16'h	5b72;
24595	:douta	=	16'h	8c73;
24596	:douta	=	16'h	9d16;
24597	:douta	=	16'h	9452;
24598	:douta	=	16'h	ddd1;
24599	:douta	=	16'h	e675;
24600	:douta	=	16'h	ddf3;
24601	:douta	=	16'h	c52f;
24602	:douta	=	16'h	a42c;
24603	:douta	=	16'h	a44c;
24604	:douta	=	16'h	8348;
24605	:douta	=	16'h	bd0e;
24606	:douta	=	16'h	bcee;
24607	:douta	=	16'h	bd0f;
24608	:douta	=	16'h	c50e;
24609	:douta	=	16'h	de13;
24610	:douta	=	16'h	d5d2;
24611	:douta	=	16'h	e675;
24612	:douta	=	16'h	de54;
24613	:douta	=	16'h	e696;
24614	:douta	=	16'h	e655;
24615	:douta	=	16'h	eeb7;
24616	:douta	=	16'h	e655;
24617	:douta	=	16'h	eed8;
24618	:douta	=	16'h	ee96;
24619	:douta	=	16'h	ee75;
24620	:douta	=	16'h	ddf3;
24621	:douta	=	16'h	de13;
24622	:douta	=	16'h	cd50;
24623	:douta	=	16'h	9c0d;
24624	:douta	=	16'h	d591;
24625	:douta	=	16'h	cd70;
24626	:douta	=	16'h	ac50;
24627	:douta	=	16'h	9c70;
24628	:douta	=	16'h	9c50;
24629	:douta	=	16'h	83cf;
24630	:douta	=	16'h	736d;
24631	:douta	=	16'h	6b2c;
24632	:douta	=	16'h	62cc;
24633	:douta	=	16'h	62cc;
24634	:douta	=	16'h	2905;
24635	:douta	=	16'h	b42a;
24636	:douta	=	16'h	cd2d;
24637	:douta	=	16'h	b46b;
24638	:douta	=	16'h	c4ed;
24639	:douta	=	16'h	cd4f;
24640	:douta	=	16'h	e654;
24641	:douta	=	16'h	e634;
24642	:douta	=	16'h	f6b6;
24643	:douta	=	16'h	ee96;
24644	:douta	=	16'h	e654;
24645	:douta	=	16'h	e654;
24646	:douta	=	16'h	e654;
24647	:douta	=	16'h	ddb1;
24648	:douta	=	16'h	ddb1;
24649	:douta	=	16'h	ddd2;
24650	:douta	=	16'h	bd12;
24651	:douta	=	16'h	ac91;
24652	:douta	=	16'h	d5b2;
24653	:douta	=	16'h	b4f1;
24654	:douta	=	16'h	9c92;
24655	:douta	=	16'h	acd3;
24656	:douta	=	16'h	a4d3;
24657	:douta	=	16'h	9c73;
24658	:douta	=	16'h	9473;
24659	:douta	=	16'h	8c53;
24660	:douta	=	16'h	8412;
24661	:douta	=	16'h	7bf2;
24662	:douta	=	16'h	7390;
24663	:douta	=	16'h	736f;
24664	:douta	=	16'h	732e;
24665	:douta	=	16'h	6b2e;
24666	:douta	=	16'h	632e;
24667	:douta	=	16'h	5229;
24668	:douta	=	16'h	6228;
24669	:douta	=	16'h	abca;
24670	:douta	=	16'h	b3eb;
24671	:douta	=	16'h	cd0e;
24672	:douta	=	16'h	ddd1;
24673	:douta	=	16'h	ddf2;
24674	:douta	=	16'h	e654;
24675	:douta	=	16'h	e634;
24676	:douta	=	16'h	e613;
24677	:douta	=	16'h	ddf2;
24678	:douta	=	16'h	cd71;
24679	:douta	=	16'h	8c10;
24680	:douta	=	16'h	83f1;
24681	:douta	=	16'h	8c11;
24682	:douta	=	16'h	8c32;
24683	:douta	=	16'h	7433;
24684	:douta	=	16'h	3a6d;
24685	:douta	=	16'h	52ef;
24686	:douta	=	16'h	426d;
24687	:douta	=	16'h	322c;
24688	:douta	=	16'h	2a0b;
24689	:douta	=	16'h	29eb;
24690	:douta	=	16'h	21a9;
24691	:douta	=	16'h	2127;
24692	:douta	=	16'h	2107;
24693	:douta	=	16'h	5b30;
24694	:douta	=	16'h	10c4;
24695	:douta	=	16'h	1063;
24696	:douta	=	16'h	10c4;
24697	:douta	=	16'h	10a4;
24698	:douta	=	16'h	10c5;
24699	:douta	=	16'h	10c5;
24700	:douta	=	16'h	10e4;
24701	:douta	=	16'h	18e5;
24702	:douta	=	16'h	18e4;
24703	:douta	=	16'h	10a4;
24704	:douta	=	16'h	2147;
24705	:douta	=	16'h	18e4;
24706	:douta	=	16'h	10e5;
24707	:douta	=	16'h	2167;
24708	:douta	=	16'h	0842;
24709	:douta	=	16'h	10e5;
24710	:douta	=	16'h	10c4;
24711	:douta	=	16'h	0883;
24712	:douta	=	16'h	9cf5;
24713	:douta	=	16'h	a4b1;
24714	:douta	=	16'h	b573;
24715	:douta	=	16'h	9c90;
24716	:douta	=	16'h	29aa;
24717	:douta	=	16'h	959a;
24718	:douta	=	16'h	a5db;
24719	:douta	=	16'h	a5da;
24720	:douta	=	16'h	a5ba;
24721	:douta	=	16'h	957a;
24722	:douta	=	16'h	9559;
24723	:douta	=	16'h	8d18;
24724	:douta	=	16'h	9559;
24725	:douta	=	16'h	8d38;
24726	:douta	=	16'h	84d7;
24727	:douta	=	16'h	84d7;
24728	:douta	=	16'h	7c96;
24729	:douta	=	16'h	8d18;
24730	:douta	=	16'h	8d59;
24731	:douta	=	16'h	8d18;
24732	:douta	=	16'h	7cb7;
24733	:douta	=	16'h	84f8;
24734	:douta	=	16'h	9dba;
24735	:douta	=	16'h	9dba;
24736	:douta	=	16'h	7cb6;
24737	:douta	=	16'h	957a;
24738	:douta	=	16'h	9559;
24739	:douta	=	16'h	8d39;
24740	:douta	=	16'h	84f8;
24741	:douta	=	16'h	957a;
24742	:douta	=	16'h	8d18;
24743	:douta	=	16'h	84b7;
24744	:douta	=	16'h	7476;
24745	:douta	=	16'h	8d18;
24746	:douta	=	16'h	7c55;
24747	:douta	=	16'h	6bb3;
24748	:douta	=	16'h	7434;
24749	:douta	=	16'h	84b7;
24750	:douta	=	16'h	6bd4;
24751	:douta	=	16'h	5b93;
24752	:douta	=	16'h	7cb7;
24753	:douta	=	16'h	8d39;
24754	:douta	=	16'h	7d18;
24755	:douta	=	16'h	8519;
24756	:douta	=	16'h	7cf8;
24757	:douta	=	16'h	8519;
24758	:douta	=	16'h	8539;
24759	:douta	=	16'h	8d5b;
24760	:douta	=	16'h	851a;
24761	:douta	=	16'h	7cd8;
24762	:douta	=	16'h	8539;
24763	:douta	=	16'h	84f8;
24764	:douta	=	16'h	95bb;
24765	:douta	=	16'h	957a;
24766	:douta	=	16'h	8539;
24767	:douta	=	16'h	84f8;
24768	:douta	=	16'h	84f8;
24769	:douta	=	16'h	8d39;
24770	:douta	=	16'h	8d59;
24771	:douta	=	16'h	9d9a;
24772	:douta	=	16'h	8518;
24773	:douta	=	16'h	7cd7;
24774	:douta	=	16'h	959a;
24775	:douta	=	16'h	9dbb;
24776	:douta	=	16'h	8d59;
24777	:douta	=	16'h	957a;
24778	:douta	=	16'h	8d5a;
24779	:douta	=	16'h	959a;
24780	:douta	=	16'h	9dbb;
24781	:douta	=	16'h	8518;
24782	:douta	=	16'h	959a;
24783	:douta	=	16'h	adfc;
24784	:douta	=	16'h	9d9a;
24785	:douta	=	16'h	9559;
24786	:douta	=	16'h	959a;
24787	:douta	=	16'h	9dbb;
24788	:douta	=	16'h	8d5a;
24789	:douta	=	16'h	959b;
24790	:douta	=	16'h	8d5a;
24791	:douta	=	16'h	ae3c;
24792	:douta	=	16'h	b67d;
24793	:douta	=	16'h	a5fb;
24794	:douta	=	16'h	a61d;
24795	:douta	=	16'h	a61c;
24796	:douta	=	16'h	632e;
24797	:douta	=	16'h	6b2f;
24798	:douta	=	16'h	4bf7;
24799	:douta	=	16'h	6478;
24800	:douta	=	16'h	5c57;
24801	:douta	=	16'h	6c99;
24802	:douta	=	16'h	53f5;
24803	:douta	=	16'h	6498;
24804	:douta	=	16'h	5c78;
24805	:douta	=	16'h	4b0f;
24806	:douta	=	16'h	8308;
24807	:douta	=	16'h	72a6;
24808	:douta	=	16'h	2923;
24809	:douta	=	16'h	0863;
24810	:douta	=	16'h	0862;
24811	:douta	=	16'h	1926;
24812	:douta	=	16'h	4bd4;
24813	:douta	=	16'h	959b;
24814	:douta	=	16'h	a535;
24815	:douta	=	16'h	4060;
24816	:douta	=	16'h	7d3c;
24817	:douta	=	16'h	4b52;
24818	:douta	=	16'h	63d4;
24819	:douta	=	16'h	734b;
24820	:douta	=	16'h	1800;
24821	:douta	=	16'h	7c97;
24822	:douta	=	16'h	5bb3;
24823	:douta	=	16'h	5bb4;
24824	:douta	=	16'h	4b32;
24825	:douta	=	16'h	3ab0;
24826	:douta	=	16'h	6bd3;
24827	:douta	=	16'h	7455;
24828	:douta	=	16'h	5310;
24829	:douta	=	16'h	18e5;
24830	:douta	=	16'h	7433;
24831	:douta	=	16'h	5b8f;
24832	:douta	=	16'h	3104;
24833	:douta	=	16'h	3966;
24834	:douta	=	16'h	3966;
24835	:douta	=	16'h	2925;
24836	:douta	=	16'h	2126;
24837	:douta	=	16'h	3a6e;
24838	:douta	=	16'h	4353;
24839	:douta	=	16'h	42f1;
24840	:douta	=	16'h	3af1;
24841	:douta	=	16'h	32b0;
24842	:douta	=	16'h	4b12;
24843	:douta	=	16'h	6436;
24844	:douta	=	16'h	5bf5;
24845	:douta	=	16'h	7456;
24846	:douta	=	16'h	6c15;
24847	:douta	=	16'h	5b93;
24848	:douta	=	16'h	7414;
24849	:douta	=	16'h	8cb6;
24850	:douta	=	16'h	73f4;
24851	:douta	=	16'h	9d16;
24852	:douta	=	16'h	9494;
24853	:douta	=	16'h	6bb1;
24854	:douta	=	16'h	ad15;
24855	:douta	=	16'h	e653;
24856	:douta	=	16'h	7b4c;
24857	:douta	=	16'h	ac8f;
24858	:douta	=	16'h	9beb;
24859	:douta	=	16'h	9389;
24860	:douta	=	16'h	c50f;
24861	:douta	=	16'h	cd50;
24862	:douta	=	16'h	c570;
24863	:douta	=	16'h	cd90;
24864	:douta	=	16'h	c56f;
24865	:douta	=	16'h	e634;
24866	:douta	=	16'h	e655;
24867	:douta	=	16'h	eeb7;
24868	:douta	=	16'h	eeb7;
24869	:douta	=	16'h	e675;
24870	:douta	=	16'h	eeb7;
24871	:douta	=	16'h	eeb7;
24872	:douta	=	16'h	ee96;
24873	:douta	=	16'h	e675;
24874	:douta	=	16'h	eeb7;
24875	:douta	=	16'h	ddf3;
24876	:douta	=	16'h	de13;
24877	:douta	=	16'h	d5d2;
24878	:douta	=	16'h	cd72;
24879	:douta	=	16'h	d591;
24880	:douta	=	16'h	a450;
24881	:douta	=	16'h	a450;
24882	:douta	=	16'h	c551;
24883	:douta	=	16'h	8c10;
24884	:douta	=	16'h	736f;
24885	:douta	=	16'h	736e;
24886	:douta	=	16'h	6b2c;
24887	:douta	=	16'h	6b0c;
24888	:douta	=	16'h	5a8b;
24889	:douta	=	16'h	3966;
24890	:douta	=	16'h	bc6a;
24891	:douta	=	16'h	b48c;
24892	:douta	=	16'h	cd0e;
24893	:douta	=	16'h	d5b0;
24894	:douta	=	16'h	e5f3;
24895	:douta	=	16'h	e634;
24896	:douta	=	16'h	ee54;
24897	:douta	=	16'h	ee76;
24898	:douta	=	16'h	ee95;
24899	:douta	=	16'h	e634;
24900	:douta	=	16'h	e634;
24901	:douta	=	16'h	de13;
24902	:douta	=	16'h	ddd1;
24903	:douta	=	16'h	d5d1;
24904	:douta	=	16'h	d5d1;
24905	:douta	=	16'h	cd71;
24906	:douta	=	16'h	c531;
24907	:douta	=	16'h	acb1;
24908	:douta	=	16'h	9431;
24909	:douta	=	16'h	c552;
24910	:douta	=	16'h	a4b2;
24911	:douta	=	16'h	9473;
24912	:douta	=	16'h	9cb3;
24913	:douta	=	16'h	9c93;
24914	:douta	=	16'h	9c94;
24915	:douta	=	16'h	8432;
24916	:douta	=	16'h	83f1;
24917	:douta	=	16'h	7390;
24918	:douta	=	16'h	6b2e;
24919	:douta	=	16'h	6b0e;
24920	:douta	=	16'h	736f;
24921	:douta	=	16'h	6b2e;
24922	:douta	=	16'h	51a6;
24923	:douta	=	16'h	8b48;
24924	:douta	=	16'h	9b8a;
24925	:douta	=	16'h	c4eb;
24926	:douta	=	16'h	d54e;
24927	:douta	=	16'h	ddf2;
24928	:douta	=	16'h	e654;
24929	:douta	=	16'h	e654;
24930	:douta	=	16'h	e634;
24931	:douta	=	16'h	e674;
24932	:douta	=	16'h	de12;
24933	:douta	=	16'h	d571;
24934	:douta	=	16'h	c510;
24935	:douta	=	16'h	9c51;
24936	:douta	=	16'h	9451;
24937	:douta	=	16'h	83f1;
24938	:douta	=	16'h	8433;
24939	:douta	=	16'h	8c54;
24940	:douta	=	16'h	6bf3;
24941	:douta	=	16'h	5b51;
24942	:douta	=	16'h	5330;
24943	:douta	=	16'h	3a8d;
24944	:douta	=	16'h	3a6d;
24945	:douta	=	16'h	322b;
24946	:douta	=	16'h	322b;
24947	:douta	=	16'h	2168;
24948	:douta	=	16'h	18e5;
24949	:douta	=	16'h	10c3;
24950	:douta	=	16'h	31ea;
24951	:douta	=	16'h	5330;
24952	:douta	=	16'h	0042;
24953	:douta	=	16'h	18e5;
24954	:douta	=	16'h	18c4;
24955	:douta	=	16'h	1905;
24956	:douta	=	16'h	18e5;
24957	:douta	=	16'h	10e4;
24958	:douta	=	16'h	10a4;
24959	:douta	=	16'h	10c4;
24960	:douta	=	16'h	18e5;
24961	:douta	=	16'h	10c5;
24962	:douta	=	16'h	1926;
24963	:douta	=	16'h	0021;
24964	:douta	=	16'h	0863;
24965	:douta	=	16'h	2146;
24966	:douta	=	16'h	1905;
24967	:douta	=	16'h	1105;
24968	:douta	=	16'h	0003;
24969	:douta	=	16'h	3188;
24970	:douta	=	16'h	ad32;
24971	:douta	=	16'h	3a28;
24972	:douta	=	16'h	9450;
24973	:douta	=	16'h	31c8;
24974	:douta	=	16'h	31c9;
24975	:douta	=	16'h	7435;
24976	:douta	=	16'h	9d9a;
24977	:douta	=	16'h	84d7;
24978	:douta	=	16'h	9559;
24979	:douta	=	16'h	a5da;
24980	:douta	=	16'h	9579;
24981	:douta	=	16'h	9559;
24982	:douta	=	16'h	9d9a;
24983	:douta	=	16'h	8d59;
24984	:douta	=	16'h	7cb7;
24985	:douta	=	16'h	8d18;
24986	:douta	=	16'h	8d39;
24987	:douta	=	16'h	8cd8;
24988	:douta	=	16'h	7cb7;
24989	:douta	=	16'h	6c14;
24990	:douta	=	16'h	84f8;
24991	:douta	=	16'h	84f8;
24992	:douta	=	16'h	9559;
24993	:douta	=	16'h	84d7;
24994	:douta	=	16'h	6c55;
24995	:douta	=	16'h	63d4;
24996	:douta	=	16'h	7476;
24997	:douta	=	16'h	9d9a;
24998	:douta	=	16'h	8d39;
24999	:douta	=	16'h	8d59;
25000	:douta	=	16'h	8d39;
25001	:douta	=	16'h	8d39;
25002	:douta	=	16'h	8d18;
25003	:douta	=	16'h	84f7;
25004	:douta	=	16'h	7c76;
25005	:douta	=	16'h	7c56;
25006	:douta	=	16'h	84d7;
25007	:douta	=	16'h	8d59;
25008	:douta	=	16'h	8518;
25009	:douta	=	16'h	8d39;
25010	:douta	=	16'h	5b93;
25011	:douta	=	16'h	7c77;
25012	:douta	=	16'h	8519;
25013	:douta	=	16'h	8519;
25014	:douta	=	16'h	8519;
25015	:douta	=	16'h	8539;
25016	:douta	=	16'h	8519;
25017	:douta	=	16'h	8d39;
25018	:douta	=	16'h	8d39;
25019	:douta	=	16'h	8539;
25020	:douta	=	16'h	8539;
25021	:douta	=	16'h	7cd8;
25022	:douta	=	16'h	7cd8;
25023	:douta	=	16'h	8d5a;
25024	:douta	=	16'h	8d59;
25025	:douta	=	16'h	8d59;
25026	:douta	=	16'h	8d18;
25027	:douta	=	16'h	84f8;
25028	:douta	=	16'h	957a;
25029	:douta	=	16'h	8d3a;
25030	:douta	=	16'h	955a;
25031	:douta	=	16'h	84f8;
25032	:douta	=	16'h	84f9;
25033	:douta	=	16'h	8518;
25034	:douta	=	16'h	9dbb;
25035	:douta	=	16'h	957a;
25036	:douta	=	16'h	8539;
25037	:douta	=	16'h	8d5a;
25038	:douta	=	16'h	957a;
25039	:douta	=	16'h	959a;
25040	:douta	=	16'h	95ba;
25041	:douta	=	16'h	8539;
25042	:douta	=	16'h	9dba;
25043	:douta	=	16'h	9d9a;
25044	:douta	=	16'h	ae1b;
25045	:douta	=	16'h	a5db;
25046	:douta	=	16'h	a5fb;
25047	:douta	=	16'h	95dc;
25048	:douta	=	16'h	959c;
25049	:douta	=	16'h	6b70;
25050	:douta	=	16'h	39ea;
25051	:douta	=	16'h	4b32;
25052	:douta	=	16'h	7dbe;
25053	:douta	=	16'h	4bf7;
25054	:douta	=	16'h	5c37;
25055	:douta	=	16'h	4bb5;
25056	:douta	=	16'h	53d6;
25057	:douta	=	16'h	53b5;
25058	:douta	=	16'h	53f6;
25059	:douta	=	16'h	6cba;
25060	:douta	=	16'h	4c16;
25061	:douta	=	16'h	7d5c;
25062	:douta	=	16'h	72a6;
25063	:douta	=	16'h	8328;
25064	:douta	=	16'h	51c5;
25065	:douta	=	16'h	20c2;
25066	:douta	=	16'h	0862;
25067	:douta	=	16'h	0820;
25068	:douta	=	16'h	0884;
25069	:douta	=	16'h	74d9;
25070	:douta	=	16'h	857b;
25071	:douta	=	16'h	7d5b;
25072	:douta	=	16'h	3060;
25073	:douta	=	16'h	2a8e;
25074	:douta	=	16'h	74da;
25075	:douta	=	16'h	2000;
25076	:douta	=	16'h	42cf;
25077	:douta	=	16'h	955a;
25078	:douta	=	16'h	6415;
25079	:douta	=	16'h	7455;
25080	:douta	=	16'h	84f8;
25081	:douta	=	16'h	957a;
25082	:douta	=	16'h	8517;
25083	:douta	=	16'h	6bf3;
25084	:douta	=	16'h	6baf;
25085	:douta	=	16'h	bdb5;
25086	:douta	=	16'h	bdb5;
25087	:douta	=	16'h	deba;
25088	:douta	=	16'h	3945;
25089	:douta	=	16'h	4187;
25090	:douta	=	16'h	3966;
25091	:douta	=	16'h	2945;
25092	:douta	=	16'h	1083;
25093	:douta	=	16'h	3a0b;
25094	:douta	=	16'h	5bf7;
25095	:douta	=	16'h	32b0;
25096	:douta	=	16'h	4333;
25097	:douta	=	16'h	3ad1;
25098	:douta	=	16'h	5373;
25099	:douta	=	16'h	5c15;
25100	:douta	=	16'h	5bd4;
25101	:douta	=	16'h	6c56;
25102	:douta	=	16'h	7498;
25103	:douta	=	16'h	5351;
25104	:douta	=	16'h	5b92;
25105	:douta	=	16'h	6c14;
25106	:douta	=	16'h	5b72;
25107	:douta	=	16'h	9d36;
25108	:douta	=	16'h	8cb4;
25109	:douta	=	16'h	8432;
25110	:douta	=	16'h	ad57;
25111	:douta	=	16'h	ee95;
25112	:douta	=	16'h	836c;
25113	:douta	=	16'h	5247;
25114	:douta	=	16'h	ac6c;
25115	:douta	=	16'h	bcee;
25116	:douta	=	16'h	c530;
25117	:douta	=	16'h	cdb1;
25118	:douta	=	16'h	cd91;
25119	:douta	=	16'h	d5b1;
25120	:douta	=	16'h	cdb1;
25121	:douta	=	16'h	e655;
25122	:douta	=	16'h	ee96;
25123	:douta	=	16'h	eeb7;
25124	:douta	=	16'h	ee96;
25125	:douta	=	16'h	ee96;
25126	:douta	=	16'h	e675;
25127	:douta	=	16'h	eeb7;
25128	:douta	=	16'h	ee97;
25129	:douta	=	16'h	de34;
25130	:douta	=	16'h	ee96;
25131	:douta	=	16'h	d613;
25132	:douta	=	16'h	d5d2;
25133	:douta	=	16'h	d5d2;
25134	:douta	=	16'h	bd30;
25135	:douta	=	16'h	bd30;
25136	:douta	=	16'h	b4f1;
25137	:douta	=	16'h	8bf0;
25138	:douta	=	16'h	a430;
25139	:douta	=	16'h	a4b1;
25140	:douta	=	16'h	7baf;
25141	:douta	=	16'h	6b2c;
25142	:douta	=	16'h	62eb;
25143	:douta	=	16'h	6b0d;
25144	:douta	=	16'h	3125;
25145	:douta	=	16'h	7a65;
25146	:douta	=	16'h	bcab;
25147	:douta	=	16'h	c4cc;
25148	:douta	=	16'h	c4ec;
25149	:douta	=	16'h	d5b1;
25150	:douta	=	16'h	ddd2;
25151	:douta	=	16'h	de14;
25152	:douta	=	16'h	ee95;
25153	:douta	=	16'h	e634;
25154	:douta	=	16'h	eeb7;
25155	:douta	=	16'h	e654;
25156	:douta	=	16'h	e614;
25157	:douta	=	16'h	de12;
25158	:douta	=	16'h	ddf2;
25159	:douta	=	16'h	cd30;
25160	:douta	=	16'h	cd50;
25161	:douta	=	16'h	c530;
25162	:douta	=	16'h	bd11;
25163	:douta	=	16'h	bcf1;
25164	:douta	=	16'h	8bf1;
25165	:douta	=	16'h	9452;
25166	:douta	=	16'h	bd53;
25167	:douta	=	16'h	8c52;
25168	:douta	=	16'h	9473;
25169	:douta	=	16'h	9c94;
25170	:douta	=	16'h	8c53;
25171	:douta	=	16'h	7bf1;
25172	:douta	=	16'h	7bd0;
25173	:douta	=	16'h	734f;
25174	:douta	=	16'h	732e;
25175	:douta	=	16'h	630e;
25176	:douta	=	16'h	6b0d;
25177	:douta	=	16'h	4a08;
25178	:douta	=	16'h	7aa7;
25179	:douta	=	16'h	ac09;
25180	:douta	=	16'h	b46b;
25181	:douta	=	16'h	c4cc;
25182	:douta	=	16'h	ddaf;
25183	:douta	=	16'h	e612;
25184	:douta	=	16'h	e654;
25185	:douta	=	16'h	e634;
25186	:douta	=	16'h	e613;
25187	:douta	=	16'h	de13;
25188	:douta	=	16'h	ddd1;
25189	:douta	=	16'h	cd30;
25190	:douta	=	16'h	c511;
25191	:douta	=	16'h	a470;
25192	:douta	=	16'h	a491;
25193	:douta	=	16'h	8c12;
25194	:douta	=	16'h	8453;
25195	:douta	=	16'h	8454;
25196	:douta	=	16'h	7c34;
25197	:douta	=	16'h	6bf3;
25198	:douta	=	16'h	5b71;
25199	:douta	=	16'h	42cf;
25200	:douta	=	16'h	42ae;
25201	:douta	=	16'h	3a4c;
25202	:douta	=	16'h	3a2c;
25203	:douta	=	16'h	322c;
25204	:douta	=	16'h	2167;
25205	:douta	=	16'h	1947;
25206	:douta	=	16'h	08a3;
25207	:douta	=	16'h	29a9;
25208	:douta	=	16'h	2167;
25209	:douta	=	16'h	1905;
25210	:douta	=	16'h	18e5;
25211	:douta	=	16'h	18e5;
25212	:douta	=	16'h	10e4;
25213	:douta	=	16'h	10a4;
25214	:douta	=	16'h	10c5;
25215	:douta	=	16'h	18e4;
25216	:douta	=	16'h	10c5;
25217	:douta	=	16'h	18e5;
25218	:douta	=	16'h	10c4;
25219	:douta	=	16'h	2126;
25220	:douta	=	16'h	0883;
25221	:douta	=	16'h	10a4;
25222	:douta	=	16'h	1926;
25223	:douta	=	16'h	1905;
25224	:douta	=	16'h	10a4;
25225	:douta	=	16'h	0864;
25226	:douta	=	16'h	d655;
25227	:douta	=	16'h	944e;
25228	:douta	=	16'h	c5f4;
25229	:douta	=	16'h	9450;
25230	:douta	=	16'h	39e8;
25231	:douta	=	16'h	630d;
25232	:douta	=	16'h	428d;
25233	:douta	=	16'h	8d59;
25234	:douta	=	16'h	8d39;
25235	:douta	=	16'h	84d7;
25236	:douta	=	16'h	9579;
25237	:douta	=	16'h	957a;
25238	:douta	=	16'h	9dba;
25239	:douta	=	16'h	9d9a;
25240	:douta	=	16'h	84f8;
25241	:douta	=	16'h	8d39;
25242	:douta	=	16'h	7455;
25243	:douta	=	16'h	9d9a;
25244	:douta	=	16'h	8d38;
25245	:douta	=	16'h	9559;
25246	:douta	=	16'h	84d7;
25247	:douta	=	16'h	84f7;
25248	:douta	=	16'h	8d38;
25249	:douta	=	16'h	84b7;
25250	:douta	=	16'h	84f8;
25251	:douta	=	16'h	7c96;
25252	:douta	=	16'h	7455;
25253	:douta	=	16'h	7cb7;
25254	:douta	=	16'h	9559;
25255	:douta	=	16'h	9559;
25256	:douta	=	16'h	8d39;
25257	:douta	=	16'h	9559;
25258	:douta	=	16'h	7cb7;
25259	:douta	=	16'h	7496;
25260	:douta	=	16'h	8d59;
25261	:douta	=	16'h	7435;
25262	:douta	=	16'h	7c75;
25263	:douta	=	16'h	8d39;
25264	:douta	=	16'h	7c97;
25265	:douta	=	16'h	9d9a;
25266	:douta	=	16'h	7496;
25267	:douta	=	16'h	7477;
25268	:douta	=	16'h	7c77;
25269	:douta	=	16'h	74b7;
25270	:douta	=	16'h	8519;
25271	:douta	=	16'h	8d3a;
25272	:douta	=	16'h	8519;
25273	:douta	=	16'h	8539;
25274	:douta	=	16'h	8519;
25275	:douta	=	16'h	8539;
25276	:douta	=	16'h	8d3a;
25277	:douta	=	16'h	957b;
25278	:douta	=	16'h	8539;
25279	:douta	=	16'h	8519;
25280	:douta	=	16'h	7497;
25281	:douta	=	16'h	8d7a;
25282	:douta	=	16'h	959a;
25283	:douta	=	16'h	959a;
25284	:douta	=	16'h	8d7a;
25285	:douta	=	16'h	8518;
25286	:douta	=	16'h	7cb7;
25287	:douta	=	16'h	8519;
25288	:douta	=	16'h	8519;
25289	:douta	=	16'h	7cd8;
25290	:douta	=	16'h	8d39;
25291	:douta	=	16'h	959a;
25292	:douta	=	16'h	959b;
25293	:douta	=	16'h	95bb;
25294	:douta	=	16'h	9ddb;
25295	:douta	=	16'h	8559;
25296	:douta	=	16'h	959b;
25297	:douta	=	16'h	8d7a;
25298	:douta	=	16'h	959a;
25299	:douta	=	16'h	8d18;
25300	:douta	=	16'h	9d9a;
25301	:douta	=	16'h	b69e;
25302	:douta	=	16'h	ae7e;
25303	:douta	=	16'h	8474;
25304	:douta	=	16'h	62ec;
25305	:douta	=	16'h	530f;
25306	:douta	=	16'h	6cb9;
25307	:douta	=	16'h	53f6;
25308	:douta	=	16'h	6457;
25309	:douta	=	16'h	6436;
25310	:douta	=	16'h	5c37;
25311	:douta	=	16'h	74fb;
25312	:douta	=	16'h	4bd6;
25313	:douta	=	16'h	4394;
25314	:douta	=	16'h	4374;
25315	:douta	=	16'h	5c17;
25316	:douta	=	16'h	64b8;
25317	:douta	=	16'h	6cd9;
25318	:douta	=	16'h	62cc;
25319	:douta	=	16'h	7ac5;
25320	:douta	=	16'h	6a44;
25321	:douta	=	16'h	20c2;
25322	:douta	=	16'h	1082;
25323	:douta	=	16'h	1063;
25324	:douta	=	16'h	0000;
25325	:douta	=	16'h	6c77;
25326	:douta	=	16'h	7477;
25327	:douta	=	16'h	53f5;
25328	:douta	=	16'h	7aeb;
25329	:douta	=	16'h	3880;
25330	:douta	=	16'h	85bd;
25331	:douta	=	16'h	1882;
25332	:douta	=	16'h	6478;
25333	:douta	=	16'h	6c35;
25334	:douta	=	16'h	6435;
25335	:douta	=	16'h	7497;
25336	:douta	=	16'h	9dba;
25337	:douta	=	16'h	6c35;
25338	:douta	=	16'h	5b2e;
25339	:douta	=	16'h	8472;
25340	:douta	=	16'h	9d14;
25341	:douta	=	16'h	deda;
25342	:douta	=	16'h	c638;
25343	:douta	=	16'h	a5d8;
25344	:douta	=	16'h	526b;
25345	:douta	=	16'h	3966;
25346	:douta	=	16'h	3966;
25347	:douta	=	16'h	3145;
25348	:douta	=	16'h	1882;
25349	:douta	=	16'h	31a8;
25350	:douta	=	16'h	4332;
25351	:douta	=	16'h	4333;
25352	:douta	=	16'h	3ad1;
25353	:douta	=	16'h	3ad1;
25354	:douta	=	16'h	2a4f;
25355	:douta	=	16'h	5bb4;
25356	:douta	=	16'h	6436;
25357	:douta	=	16'h	7c98;
25358	:douta	=	16'h	63f5;
25359	:douta	=	16'h	6c35;
25360	:douta	=	16'h	6bf4;
25361	:douta	=	16'h	6bd3;
25362	:douta	=	16'h	6bd3;
25363	:douta	=	16'h	8433;
25364	:douta	=	16'h	9cb5;
25365	:douta	=	16'h	94d5;
25366	:douta	=	16'h	8c73;
25367	:douta	=	16'h	b5b8;
25368	:douta	=	16'h	c551;
25369	:douta	=	16'h	a40b;
25370	:douta	=	16'h	c54f;
25371	:douta	=	16'h	c530;
25372	:douta	=	16'h	c551;
25373	:douta	=	16'h	d5f3;
25374	:douta	=	16'h	d5d2;
25375	:douta	=	16'h	de15;
25376	:douta	=	16'h	de14;
25377	:douta	=	16'h	eeb6;
25378	:douta	=	16'h	eed7;
25379	:douta	=	16'h	eeb6;
25380	:douta	=	16'h	ee96;
25381	:douta	=	16'h	eeb6;
25382	:douta	=	16'h	ee96;
25383	:douta	=	16'h	d591;
25384	:douta	=	16'h	de34;
25385	:douta	=	16'h	e675;
25386	:douta	=	16'h	de13;
25387	:douta	=	16'h	d5b2;
25388	:douta	=	16'h	bd11;
25389	:douta	=	16'h	bcf1;
25390	:douta	=	16'h	a4b1;
25391	:douta	=	16'h	9450;
25392	:douta	=	16'h	9450;
25393	:douta	=	16'h	8c10;
25394	:douta	=	16'h	7b8f;
25395	:douta	=	16'h	838e;
25396	:douta	=	16'h	7baf;
25397	:douta	=	16'h	736d;
25398	:douta	=	16'h	528a;
25399	:douta	=	16'h	3945;
25400	:douta	=	16'h	bc6a;
25401	:douta	=	16'h	bccc;
25402	:douta	=	16'h	c50e;
25403	:douta	=	16'h	d570;
25404	:douta	=	16'h	d56f;
25405	:douta	=	16'h	ee54;
25406	:douta	=	16'h	e674;
25407	:douta	=	16'h	ee74;
25408	:douta	=	16'h	ee75;
25409	:douta	=	16'h	ddf2;
25410	:douta	=	16'h	e674;
25411	:douta	=	16'h	f6b6;
25412	:douta	=	16'h	ddd2;
25413	:douta	=	16'h	d5b2;
25414	:douta	=	16'h	dd91;
25415	:douta	=	16'h	cd71;
25416	:douta	=	16'h	b4cf;
25417	:douta	=	16'h	b4d1;
25418	:douta	=	16'h	b4f2;
25419	:douta	=	16'h	a491;
25420	:douta	=	16'h	9c72;
25421	:douta	=	16'h	9453;
25422	:douta	=	16'h	8412;
25423	:douta	=	16'h	a4b4;
25424	:douta	=	16'h	83f1;
25425	:douta	=	16'h	7bf1;
25426	:douta	=	16'h	8c52;
25427	:douta	=	16'h	7bd1;
25428	:douta	=	16'h	6b2e;
25429	:douta	=	16'h	6b2e;
25430	:douta	=	16'h	632e;
25431	:douta	=	16'h	4a4a;
25432	:douta	=	16'h	59a5;
25433	:douta	=	16'h	9329;
25434	:douta	=	16'h	a3ea;
25435	:douta	=	16'h	c4cc;
25436	:douta	=	16'h	dd90;
25437	:douta	=	16'h	e632;
25438	:douta	=	16'h	e653;
25439	:douta	=	16'h	e654;
25440	:douta	=	16'h	e634;
25441	:douta	=	16'h	e633;
25442	:douta	=	16'h	ddf3;
25443	:douta	=	16'h	ddd3;
25444	:douta	=	16'h	d591;
25445	:douta	=	16'h	c4f0;
25446	:douta	=	16'h	b4af;
25447	:douta	=	16'h	a491;
25448	:douta	=	16'h	ac92;
25449	:douta	=	16'h	9432;
25450	:douta	=	16'h	8433;
25451	:douta	=	16'h	7c13;
25452	:douta	=	16'h	7c34;
25453	:douta	=	16'h	8454;
25454	:douta	=	16'h	73f3;
25455	:douta	=	16'h	5bb2;
25456	:douta	=	16'h	5b71;
25457	:douta	=	16'h	4aef;
25458	:douta	=	16'h	4aef;
25459	:douta	=	16'h	3a6d;
25460	:douta	=	16'h	324d;
25461	:douta	=	16'h	3a4e;
25462	:douta	=	16'h	3a8e;
25463	:douta	=	16'h	3aae;
25464	:douta	=	16'h	21ca;
25465	:douta	=	16'h	322b;
25466	:douta	=	16'h	10a4;
25467	:douta	=	16'h	10e5;
25468	:douta	=	16'h	10c4;
25469	:douta	=	16'h	10c4;
25470	:douta	=	16'h	10c4;
25471	:douta	=	16'h	10c4;
25472	:douta	=	16'h	10c4;
25473	:douta	=	16'h	18c4;
25474	:douta	=	16'h	10c5;
25475	:douta	=	16'h	18e5;
25476	:douta	=	16'h	1905;
25477	:douta	=	16'h	2126;
25478	:douta	=	16'h	10c5;
25479	:douta	=	16'h	0883;
25480	:douta	=	16'h	10a5;
25481	:douta	=	16'h	424a;
25482	:douta	=	16'h	63b3;
25483	:douta	=	16'h	7412;
25484	:douta	=	16'h	52cd;
25485	:douta	=	16'h	3166;
25486	:douta	=	16'h	736c;
25487	:douta	=	16'h	52cb;
25488	:douta	=	16'h	7bef;
25489	:douta	=	16'h	6b4d;
25490	:douta	=	16'h	5aec;
25491	:douta	=	16'h	6391;
25492	:douta	=	16'h	84d8;
25493	:douta	=	16'h	8d39;
25494	:douta	=	16'h	84d8;
25495	:douta	=	16'h	8497;
25496	:douta	=	16'h	84f7;
25497	:douta	=	16'h	8d39;
25498	:douta	=	16'h	84d7;
25499	:douta	=	16'h	8d18;
25500	:douta	=	16'h	a5da;
25501	:douta	=	16'h	9dba;
25502	:douta	=	16'h	9d99;
25503	:douta	=	16'h	8cf7;
25504	:douta	=	16'h	84b6;
25505	:douta	=	16'h	84b6;
25506	:douta	=	16'h	8cf7;
25507	:douta	=	16'h	84b7;
25508	:douta	=	16'h	7c96;
25509	:douta	=	16'h	959a;
25510	:douta	=	16'h	84d7;
25511	:douta	=	16'h	84d7;
25512	:douta	=	16'h	7c96;
25513	:douta	=	16'h	84d7;
25514	:douta	=	16'h	7476;
25515	:douta	=	16'h	8d39;
25516	:douta	=	16'h	8d39;
25517	:douta	=	16'h	8d39;
25518	:douta	=	16'h	7cd7;
25519	:douta	=	16'h	a5db;
25520	:douta	=	16'h	a5db;
25521	:douta	=	16'h	6c55;
25522	:douta	=	16'h	7476;
25523	:douta	=	16'h	7c96;
25524	:douta	=	16'h	8d18;
25525	:douta	=	16'h	957a;
25526	:douta	=	16'h	84f8;
25527	:douta	=	16'h	7476;
25528	:douta	=	16'h	7456;
25529	:douta	=	16'h	7cd8;
25530	:douta	=	16'h	8519;
25531	:douta	=	16'h	8519;
25532	:douta	=	16'h	7cd8;
25533	:douta	=	16'h	7cd8;
25534	:douta	=	16'h	7cf9;
25535	:douta	=	16'h	8d5a;
25536	:douta	=	16'h	8d5a;
25537	:douta	=	16'h	8539;
25538	:douta	=	16'h	8519;
25539	:douta	=	16'h	8519;
25540	:douta	=	16'h	7cf9;
25541	:douta	=	16'h	7cb8;
25542	:douta	=	16'h	957b;
25543	:douta	=	16'h	959b;
25544	:douta	=	16'h	84f9;
25545	:douta	=	16'h	8d5a;
25546	:douta	=	16'h	8d3a;
25547	:douta	=	16'h	74b8;
25548	:douta	=	16'h	6457;
25549	:douta	=	16'h	8d3a;
25550	:douta	=	16'h	957a;
25551	:douta	=	16'h	959b;
25552	:douta	=	16'h	959a;
25553	:douta	=	16'h	9ddb;
25554	:douta	=	16'h	959c;
25555	:douta	=	16'h	8d9c;
25556	:douta	=	16'h	8cf6;
25557	:douta	=	16'h	428d;
25558	:douta	=	16'h	3a4c;
25559	:douta	=	16'h	3b12;
25560	:douta	=	16'h	4c16;
25561	:douta	=	16'h	6456;
25562	:douta	=	16'h	6cf9;
25563	:douta	=	16'h	74b9;
25564	:douta	=	16'h	5c37;
25565	:douta	=	16'h	6cda;
25566	:douta	=	16'h	753b;
25567	:douta	=	16'h	3b13;
25568	:douta	=	16'h	4374;
25569	:douta	=	16'h	4353;
25570	:douta	=	16'h	4b95;
25571	:douta	=	16'h	4395;
25572	:douta	=	16'h	7d5b;
25573	:douta	=	16'h	4bf6;
25574	:douta	=	16'h	651c;
25575	:douta	=	16'h	732c;
25576	:douta	=	16'h	8329;
25577	:douta	=	16'h	4144;
25578	:douta	=	16'h	28e3;
25579	:douta	=	16'h	0882;
25580	:douta	=	16'h	0862;
25581	:douta	=	16'h	29ca;
25582	:douta	=	16'h	5c16;
25583	:douta	=	16'h	6436;
25584	:douta	=	16'h	5418;
25585	:douta	=	16'h	6cd9;
25586	:douta	=	16'h	40c0;
25587	:douta	=	16'h	5c57;
25588	:douta	=	16'h	7498;
25589	:douta	=	16'h	5bf6;
25590	:douta	=	16'h	8d18;
25591	:douta	=	16'h	63b1;
25592	:douta	=	16'h	73f0;
25593	:douta	=	16'h	a535;
25594	:douta	=	16'h	bdd6;
25595	:douta	=	16'h	add7;
25596	:douta	=	16'h	8cb3;
25597	:douta	=	16'h	4aaa;
25598	:douta	=	16'h	39a6;
25599	:douta	=	16'h	1840;
25600	:douta	=	16'h	5b0e;
25601	:douta	=	16'h	3966;
25602	:douta	=	16'h	3986;
25603	:douta	=	16'h	3146;
25604	:douta	=	16'h	1883;
25605	:douta	=	16'h	3188;
25606	:douta	=	16'h	326e;
25607	:douta	=	16'h	3ad1;
25608	:douta	=	16'h	4b53;
25609	:douta	=	16'h	4353;
25610	:douta	=	16'h	3290;
25611	:douta	=	16'h	5bd5;
25612	:douta	=	16'h	7477;
25613	:douta	=	16'h	5bb4;
25614	:douta	=	16'h	7455;
25615	:douta	=	16'h	63f4;
25616	:douta	=	16'h	8475;
25617	:douta	=	16'h	73f4;
25618	:douta	=	16'h	7c75;
25619	:douta	=	16'h	73f2;
25620	:douta	=	16'h	ad77;
25621	:douta	=	16'h	6bb1;
25622	:douta	=	16'h	6bb1;
25623	:douta	=	16'h	c63a;
25624	:douta	=	16'h	c572;
25625	:douta	=	16'h	bcee;
25626	:douta	=	16'h	c570;
25627	:douta	=	16'h	cd90;
25628	:douta	=	16'h	cdb2;
25629	:douta	=	16'h	d614;
25630	:douta	=	16'h	d5d3;
25631	:douta	=	16'h	e656;
25632	:douta	=	16'h	e655;
25633	:douta	=	16'h	eeb7;
25634	:douta	=	16'h	eed7;
25635	:douta	=	16'h	eed7;
25636	:douta	=	16'h	ee96;
25637	:douta	=	16'h	e696;
25638	:douta	=	16'h	eeb6;
25639	:douta	=	16'h	d5d2;
25640	:douta	=	16'h	c54f;
25641	:douta	=	16'h	eeb6;
25642	:douta	=	16'h	e674;
25643	:douta	=	16'h	c551;
25644	:douta	=	16'h	a4b1;
25645	:douta	=	16'h	a471;
25646	:douta	=	16'h	a4b1;
25647	:douta	=	16'h	9c51;
25648	:douta	=	16'h	7baf;
25649	:douta	=	16'h	8c10;
25650	:douta	=	16'h	8c10;
25651	:douta	=	16'h	7b6e;
25652	:douta	=	16'h	734d;
25653	:douta	=	16'h	730d;
25654	:douta	=	16'h	41a5;
25655	:douta	=	16'h	8ae8;
25656	:douta	=	16'h	bcec;
25657	:douta	=	16'h	b4ac;
25658	:douta	=	16'h	cd4f;
25659	:douta	=	16'h	ddd2;
25660	:douta	=	16'h	d5b1;
25661	:douta	=	16'h	eeb6;
25662	:douta	=	16'h	ee95;
25663	:douta	=	16'h	e674;
25664	:douta	=	16'h	e654;
25665	:douta	=	16'h	e634;
25666	:douta	=	16'h	ddf3;
25667	:douta	=	16'h	ee95;
25668	:douta	=	16'h	de13;
25669	:douta	=	16'h	cd71;
25670	:douta	=	16'h	cd31;
25671	:douta	=	16'h	cd31;
25672	:douta	=	16'h	bd10;
25673	:douta	=	16'h	ac91;
25674	:douta	=	16'h	a4b2;
25675	:douta	=	16'h	acb2;
25676	:douta	=	16'h	9c93;
25677	:douta	=	16'h	9452;
25678	:douta	=	16'h	7bf2;
25679	:douta	=	16'h	9cb3;
25680	:douta	=	16'h	9cb4;
25681	:douta	=	16'h	632e;
25682	:douta	=	16'h	7bd0;
25683	:douta	=	16'h	8412;
25684	:douta	=	16'h	734f;
25685	:douta	=	16'h	6b2f;
25686	:douta	=	16'h	41e8;
25687	:douta	=	16'h	28c3;
25688	:douta	=	16'h	9348;
25689	:douta	=	16'h	a40a;
25690	:douta	=	16'h	bc8b;
25691	:douta	=	16'h	ddaf;
25692	:douta	=	16'h	ddf2;
25693	:douta	=	16'h	e654;
25694	:douta	=	16'h	ee54;
25695	:douta	=	16'h	e633;
25696	:douta	=	16'h	e633;
25697	:douta	=	16'h	e633;
25698	:douta	=	16'h	ddf2;
25699	:douta	=	16'h	ddd3;
25700	:douta	=	16'h	d570;
25701	:douta	=	16'h	c510;
25702	:douta	=	16'h	b4b0;
25703	:douta	=	16'h	acb1;
25704	:douta	=	16'h	a491;
25705	:douta	=	16'h	9453;
25706	:douta	=	16'h	8c53;
25707	:douta	=	16'h	7c13;
25708	:douta	=	16'h	7c34;
25709	:douta	=	16'h	7c34;
25710	:douta	=	16'h	7414;
25711	:douta	=	16'h	5b92;
25712	:douta	=	16'h	5b71;
25713	:douta	=	16'h	5b51;
25714	:douta	=	16'h	5330;
25715	:douta	=	16'h	42ae;
25716	:douta	=	16'h	3a6d;
25717	:douta	=	16'h	3a8d;
25718	:douta	=	16'h	42ae;
25719	:douta	=	16'h	3a6d;
25720	:douta	=	16'h	21c9;
25721	:douta	=	16'h	5b71;
25722	:douta	=	16'h	4b0e;
25723	:douta	=	16'h	0862;
25724	:douta	=	16'h	1084;
25725	:douta	=	16'h	10c5;
25726	:douta	=	16'h	18e5;
25727	:douta	=	16'h	18e5;
25728	:douta	=	16'h	18e5;
25729	:douta	=	16'h	2126;
25730	:douta	=	16'h	1905;
25731	:douta	=	16'h	1906;
25732	:douta	=	16'h	1905;
25733	:douta	=	16'h	10e5;
25734	:douta	=	16'h	1906;
25735	:douta	=	16'h	0883;
25736	:douta	=	16'h	0062;
25737	:douta	=	16'h	2146;
25738	:douta	=	16'h	324c;
25739	:douta	=	16'h	42b0;
25740	:douta	=	16'h	7433;
25741	:douta	=	16'h	7bce;
25742	:douta	=	16'h	ded7;
25743	:douta	=	16'h	738f;
25744	:douta	=	16'h	6b2c;
25745	:douta	=	16'h	8c31;
25746	:douta	=	16'h	4229;
25747	:douta	=	16'h	3187;
25748	:douta	=	16'h	5aeb;
25749	:douta	=	16'h	5b0f;
25750	:douta	=	16'h	7cb7;
25751	:douta	=	16'h	8539;
25752	:douta	=	16'h	adfb;
25753	:douta	=	16'h	9dba;
25754	:douta	=	16'h	9559;
25755	:douta	=	16'h	7456;
25756	:douta	=	16'h	84f7;
25757	:douta	=	16'h	8d58;
25758	:douta	=	16'h	9559;
25759	:douta	=	16'h	84b7;
25760	:douta	=	16'h	84b7;
25761	:douta	=	16'h	7c76;
25762	:douta	=	16'h	84b7;
25763	:douta	=	16'h	8d18;
25764	:douta	=	16'h	8d38;
25765	:douta	=	16'h	84d7;
25766	:douta	=	16'h	7cb7;
25767	:douta	=	16'h	957a;
25768	:douta	=	16'h	6c35;
25769	:douta	=	16'h	8d18;
25770	:douta	=	16'h	6c55;
25771	:douta	=	16'h	63f4;
25772	:douta	=	16'h	8d39;
25773	:douta	=	16'h	9559;
25774	:douta	=	16'h	8d39;
25775	:douta	=	16'h	8d39;
25776	:douta	=	16'h	8d39;
25777	:douta	=	16'h	a5fb;
25778	:douta	=	16'h	6c55;
25779	:douta	=	16'h	7cb7;
25780	:douta	=	16'h	9559;
25781	:douta	=	16'h	84f8;
25782	:douta	=	16'h	6c14;
25783	:douta	=	16'h	8d39;
25784	:douta	=	16'h	9559;
25785	:douta	=	16'h	84d8;
25786	:douta	=	16'h	7455;
25787	:douta	=	16'h	7cb7;
25788	:douta	=	16'h	8d7a;
25789	:douta	=	16'h	959b;
25790	:douta	=	16'h	7497;
25791	:douta	=	16'h	7cd8;
25792	:douta	=	16'h	84f9;
25793	:douta	=	16'h	959b;
25794	:douta	=	16'h	8d7a;
25795	:douta	=	16'h	8d5a;
25796	:douta	=	16'h	8d5a;
25797	:douta	=	16'h	8519;
25798	:douta	=	16'h	8519;
25799	:douta	=	16'h	8d59;
25800	:douta	=	16'h	8d39;
25801	:douta	=	16'h	8d39;
25802	:douta	=	16'h	8d7a;
25803	:douta	=	16'h	957a;
25804	:douta	=	16'h	7cb8;
25805	:douta	=	16'h	6c76;
25806	:douta	=	16'h	74d7;
25807	:douta	=	16'h	9ddb;
25808	:douta	=	16'h	9e1d;
25809	:douta	=	16'h	8d7a;
25810	:douta	=	16'h	7c95;
25811	:douta	=	16'h	6bb1;
25812	:douta	=	16'h	42ae;
25813	:douta	=	16'h	5417;
25814	:douta	=	16'h	3312;
25815	:douta	=	16'h	4394;
25816	:douta	=	16'h	3b11;
25817	:douta	=	16'h	3b33;
25818	:douta	=	16'h	6c99;
25819	:douta	=	16'h	4393;
25820	:douta	=	16'h	6479;
25821	:douta	=	16'h	5bf7;
25822	:douta	=	16'h	6cda;
25823	:douta	=	16'h	4374;
25824	:douta	=	16'h	5c37;
25825	:douta	=	16'h	5c78;
25826	:douta	=	16'h	4b94;
25827	:douta	=	16'h	6cda;
25828	:douta	=	16'h	4354;
25829	:douta	=	16'h	3af3;
25830	:douta	=	16'h	4bd7;
25831	:douta	=	16'h	63f5;
25832	:douta	=	16'h	8b69;
25833	:douta	=	16'h	51c4;
25834	:douta	=	16'h	3123;
25835	:douta	=	16'h	1082;
25836	:douta	=	16'h	0862;
25837	:douta	=	16'h	0000;
25838	:douta	=	16'h	6c99;
25839	:douta	=	16'h	5bf5;
25840	:douta	=	16'h	74f9;
25841	:douta	=	16'h	64ba;
25842	:douta	=	16'h	4942;
25843	:douta	=	16'h	5c37;
25844	:douta	=	16'h	751b;
25845	:douta	=	16'h	7476;
25846	:douta	=	16'h	8493;
25847	:douta	=	16'h	94f3;
25848	:douta	=	16'h	bdd6;
25849	:douta	=	16'h	ce18;
25850	:douta	=	16'h	a576;
25851	:douta	=	16'h	6bcf;
25852	:douta	=	16'h	5aaa;
25853	:douta	=	16'h	1040;
25854	:douta	=	16'h	1881;
25855	:douta	=	16'h	3124;
25856	:douta	=	16'h	6413;
25857	:douta	=	16'h	3986;
25858	:douta	=	16'h	3966;
25859	:douta	=	16'h	3145;
25860	:douta	=	16'h	20c3;
25861	:douta	=	16'h	20e4;
25862	:douta	=	16'h	322d;
25863	:douta	=	16'h	3af1;
25864	:douta	=	16'h	32b0;
25865	:douta	=	16'h	4353;
25866	:douta	=	16'h	2a90;
25867	:douta	=	16'h	5394;
25868	:douta	=	16'h	5c15;
25869	:douta	=	16'h	6c14;
25870	:douta	=	16'h	84d7;
25871	:douta	=	16'h	8d18;
25872	:douta	=	16'h	5b51;
25873	:douta	=	16'h	8454;
25874	:douta	=	16'h	7c55;
25875	:douta	=	16'h	94b5;
25876	:douta	=	16'h	a516;
25877	:douta	=	16'h	94b4;
25878	:douta	=	16'h	7c12;
25879	:douta	=	16'h	c619;
25880	:douta	=	16'h	bdb7;
25881	:douta	=	16'h	cd92;
25882	:douta	=	16'h	d5d2;
25883	:douta	=	16'h	d613;
25884	:douta	=	16'h	d613;
25885	:douta	=	16'h	de55;
25886	:douta	=	16'h	de14;
25887	:douta	=	16'h	eeb7;
25888	:douta	=	16'h	eeb7;
25889	:douta	=	16'h	eeb7;
25890	:douta	=	16'h	eeb7;
25891	:douta	=	16'h	eeb6;
25892	:douta	=	16'h	ee96;
25893	:douta	=	16'h	ee96;
25894	:douta	=	16'h	e675;
25895	:douta	=	16'h	de35;
25896	:douta	=	16'h	e655;
25897	:douta	=	16'h	bcf0;
25898	:douta	=	16'h	c552;
25899	:douta	=	16'h	cd91;
25900	:douta	=	16'h	9451;
25901	:douta	=	16'h	8c31;
25902	:douta	=	16'h	7bb0;
25903	:douta	=	16'h	7b90;
25904	:douta	=	16'h	83f0;
25905	:douta	=	16'h	83b0;
25906	:douta	=	16'h	7b8f;
25907	:douta	=	16'h	7b6e;
25908	:douta	=	16'h	7b4e;
25909	:douta	=	16'h	5207;
25910	:douta	=	16'h	c4cd;
25911	:douta	=	16'h	b4cd;
25912	:douta	=	16'h	bccd;
25913	:douta	=	16'h	d570;
25914	:douta	=	16'h	ddd1;
25915	:douta	=	16'h	e654;
25916	:douta	=	16'h	ee95;
25917	:douta	=	16'h	e654;
25918	:douta	=	16'h	e634;
25919	:douta	=	16'h	e654;
25920	:douta	=	16'h	e634;
25921	:douta	=	16'h	e634;
25922	:douta	=	16'h	ddd2;
25923	:douta	=	16'h	ddd2;
25924	:douta	=	16'h	e613;
25925	:douta	=	16'h	cd72;
25926	:douta	=	16'h	c531;
25927	:douta	=	16'h	acb2;
25928	:douta	=	16'h	acb2;
25929	:douta	=	16'h	b512;
25930	:douta	=	16'h	9cb3;
25931	:douta	=	16'h	9473;
25932	:douta	=	16'h	9432;
25933	:douta	=	16'h	9452;
25934	:douta	=	16'h	8432;
25935	:douta	=	16'h	6b6f;
25936	:douta	=	16'h	736f;
25937	:douta	=	16'h	7bd1;
25938	:douta	=	16'h	6b2e;
25939	:douta	=	16'h	73b0;
25940	:douta	=	16'h	62cc;
25941	:douta	=	16'h	5a27;
25942	:douta	=	16'h	8b08;
25943	:douta	=	16'h	a3e9;
25944	:douta	=	16'h	d52f;
25945	:douta	=	16'h	ddb1;
25946	:douta	=	16'h	e5f2;
25947	:douta	=	16'h	e654;
25948	:douta	=	16'h	ee74;
25949	:douta	=	16'h	de12;
25950	:douta	=	16'h	e612;
25951	:douta	=	16'h	ee54;
25952	:douta	=	16'h	e633;
25953	:douta	=	16'h	e633;
25954	:douta	=	16'h	ddd2;
25955	:douta	=	16'h	d5b1;
25956	:douta	=	16'h	c52f;
25957	:douta	=	16'h	c510;
25958	:douta	=	16'h	bcf0;
25959	:douta	=	16'h	a470;
25960	:douta	=	16'h	9c51;
25961	:douta	=	16'h	9432;
25962	:douta	=	16'h	9473;
25963	:douta	=	16'h	8c74;
25964	:douta	=	16'h	7c34;
25965	:douta	=	16'h	7c13;
25966	:douta	=	16'h	73f3;
25967	:douta	=	16'h	73f3;
25968	:douta	=	16'h	73f3;
25969	:douta	=	16'h	6392;
25970	:douta	=	16'h	5b51;
25971	:douta	=	16'h	530f;
25972	:douta	=	16'h	4b10;
25973	:douta	=	16'h	4acf;
25974	:douta	=	16'h	3a8e;
25975	:douta	=	16'h	3a6d;
25976	:douta	=	16'h	21a9;
25977	:douta	=	16'h	5330;
25978	:douta	=	16'h	2a0b;
25979	:douta	=	16'h	3a2c;
25980	:douta	=	16'h	4aef;
25981	:douta	=	16'h	1926;
25982	:douta	=	16'h	1906;
25983	:douta	=	16'h	1906;
25984	:douta	=	16'h	1906;
25985	:douta	=	16'h	10e5;
25986	:douta	=	16'h	10e5;
25987	:douta	=	16'h	2146;
25988	:douta	=	16'h	1926;
25989	:douta	=	16'h	1906;
25990	:douta	=	16'h	1926;
25991	:douta	=	16'h	10e4;
25992	:douta	=	16'h	2127;
25993	:douta	=	16'h	1083;
25994	:douta	=	16'h	0000;
25995	:douta	=	16'h	0041;
25996	:douta	=	16'h	0062;
25997	:douta	=	16'h	5b52;
25998	:douta	=	16'h	5352;
25999	:douta	=	16'h	0001;
26000	:douta	=	16'h	0022;
26001	:douta	=	16'h	29a8;
26002	:douta	=	16'h	a511;
26003	:douta	=	16'h	7b8d;
26004	:douta	=	16'h	7b8c;
26005	:douta	=	16'h	8c4f;
26006	:douta	=	16'h	62ea;
26007	:douta	=	16'h	7b6d;
26008	:douta	=	16'h	526a;
26009	:douta	=	16'h	324d;
26010	:douta	=	16'h	324c;
26011	:douta	=	16'h	8d18;
26012	:douta	=	16'h	a5db;
26013	:douta	=	16'h	9d9a;
26014	:douta	=	16'h	7cb6;
26015	:douta	=	16'h	8d38;
26016	:douta	=	16'h	84f7;
26017	:douta	=	16'h	8d38;
26018	:douta	=	16'h	7c96;
26019	:douta	=	16'h	8d18;
26020	:douta	=	16'h	8517;
26021	:douta	=	16'h	8d39;
26022	:douta	=	16'h	84d7;
26023	:douta	=	16'h	8d18;
26024	:douta	=	16'h	8d38;
26025	:douta	=	16'h	8d58;
26026	:douta	=	16'h	7c96;
26027	:douta	=	16'h	84d7;
26028	:douta	=	16'h	84d7;
26029	:douta	=	16'h	84d7;
26030	:douta	=	16'h	84f8;
26031	:douta	=	16'h	8d19;
26032	:douta	=	16'h	8d18;
26033	:douta	=	16'h	8d18;
26034	:douta	=	16'h	84f8;
26035	:douta	=	16'h	8d39;
26036	:douta	=	16'h	957a;
26037	:douta	=	16'h	8d39;
26038	:douta	=	16'h	9ddb;
26039	:douta	=	16'h	8d18;
26040	:douta	=	16'h	7c76;
26041	:douta	=	16'h	5392;
26042	:douta	=	16'h	7cb7;
26043	:douta	=	16'h	7476;
26044	:douta	=	16'h	a5fc;
26045	:douta	=	16'h	7456;
26046	:douta	=	16'h	7cd7;
26047	:douta	=	16'h	8d39;
26048	:douta	=	16'h	9d9a;
26049	:douta	=	16'h	8519;
26050	:douta	=	16'h	8d39;
26051	:douta	=	16'h	8519;
26052	:douta	=	16'h	8519;
26053	:douta	=	16'h	8519;
26054	:douta	=	16'h	7cd8;
26055	:douta	=	16'h	8539;
26056	:douta	=	16'h	8539;
26057	:douta	=	16'h	7cf9;
26058	:douta	=	16'h	8d7a;
26059	:douta	=	16'h	857b;
26060	:douta	=	16'h	95bc;
26061	:douta	=	16'h	8d39;
26062	:douta	=	16'h	6c34;
26063	:douta	=	16'h	528c;
26064	:douta	=	16'h	5a49;
26065	:douta	=	16'h	732d;
26066	:douta	=	16'h	09ac;
26067	:douta	=	16'h	1230;
26068	:douta	=	16'h	2a4e;
26069	:douta	=	16'h	5459;
26070	:douta	=	16'h	43b5;
26071	:douta	=	16'h	3b53;
26072	:douta	=	16'h	43d5;
26073	:douta	=	16'h	4bd6;
26074	:douta	=	16'h	3b13;
26075	:douta	=	16'h	53d6;
26076	:douta	=	16'h	6cb9;
26077	:douta	=	16'h	5416;
26078	:douta	=	16'h	5c58;
26079	:douta	=	16'h	5c37;
26080	:douta	=	16'h	751a;
26081	:douta	=	16'h	53d6;
26082	:douta	=	16'h	5c16;
26083	:douta	=	16'h	4bb5;
26084	:douta	=	16'h	53f6;
26085	:douta	=	16'h	5416;
26086	:douta	=	16'h	649a;
26087	:douta	=	16'h	5c9a;
26088	:douta	=	16'h	7aa6;
26089	:douta	=	16'h	72c6;
26090	:douta	=	16'h	5a04;
26091	:douta	=	16'h	20e3;
26092	:douta	=	16'h	1083;
26093	:douta	=	16'h	0861;
26094	:douta	=	16'h	4b31;
26095	:douta	=	16'h	7d7d;
26096	:douta	=	16'h	53d6;
26097	:douta	=	16'h	6436;
26098	:douta	=	16'h	1083;
26099	:douta	=	16'h	8c0e;
26100	:douta	=	16'h	8450;
26101	:douta	=	16'h	ce15;
26102	:douta	=	16'h	e6b7;
26103	:douta	=	16'h	b5d5;
26104	:douta	=	16'h	5b2c;
26105	:douta	=	16'h	39c6;
26106	:douta	=	16'h	28a1;
26107	:douta	=	16'h	28c2;
26108	:douta	=	16'h	3123;
26109	:douta	=	16'h	3944;
26110	:douta	=	16'h	3944;
26111	:douta	=	16'h	3964;
26112	:douta	=	16'h	6413;
26113	:douta	=	16'h	3945;
26114	:douta	=	16'h	41a6;
26115	:douta	=	16'h	3945;
26116	:douta	=	16'h	20e4;
26117	:douta	=	16'h	18c3;
26118	:douta	=	16'h	3a6e;
26119	:douta	=	16'h	53d6;
26120	:douta	=	16'h	3ad0;
26121	:douta	=	16'h	53d5;
26122	:douta	=	16'h	4353;
26123	:douta	=	16'h	4b74;
26124	:douta	=	16'h	5bf5;
26125	:douta	=	16'h	4b32;
26126	:douta	=	16'h	63d4;
26127	:douta	=	16'h	63f4;
26128	:douta	=	16'h	6352;
26129	:douta	=	16'h	8495;
26130	:douta	=	16'h	7434;
26131	:douta	=	16'h	8454;
26132	:douta	=	16'h	a516;
26133	:douta	=	16'h	94b4;
26134	:douta	=	16'h	9cf5;
26135	:douta	=	16'h	bdd9;
26136	:douta	=	16'h	9d37;
26137	:douta	=	16'h	cdd6;
26138	:douta	=	16'h	d5f3;
26139	:douta	=	16'h	de14;
26140	:douta	=	16'h	de34;
26141	:douta	=	16'h	e676;
26142	:douta	=	16'h	de34;
26143	:douta	=	16'h	eed7;
26144	:douta	=	16'h	eed7;
26145	:douta	=	16'h	eed7;
26146	:douta	=	16'h	eeb7;
26147	:douta	=	16'h	eeb7;
26148	:douta	=	16'h	eeb6;
26149	:douta	=	16'h	e675;
26150	:douta	=	16'h	e655;
26151	:douta	=	16'h	de13;
26152	:douta	=	16'h	ddf3;
26153	:douta	=	16'h	cd91;
26154	:douta	=	16'h	b4d0;
26155	:douta	=	16'h	acd1;
26156	:douta	=	16'h	a491;
26157	:douta	=	16'h	8c30;
26158	:douta	=	16'h	83d1;
26159	:douta	=	16'h	7bd0;
26160	:douta	=	16'h	6b4f;
26161	:douta	=	16'h	734e;
26162	:douta	=	16'h	736e;
26163	:douta	=	16'h	734d;
26164	:douta	=	16'h	628a;
26165	:douta	=	16'h	8b49;
26166	:douta	=	16'h	b4ac;
26167	:douta	=	16'h	bcce;
26168	:douta	=	16'h	cd4e;
26169	:douta	=	16'h	ddd1;
26170	:douta	=	16'h	e633;
26171	:douta	=	16'h	e654;
26172	:douta	=	16'h	e634;
26173	:douta	=	16'h	e654;
26174	:douta	=	16'h	e653;
26175	:douta	=	16'h	e654;
26176	:douta	=	16'h	e613;
26177	:douta	=	16'h	de13;
26178	:douta	=	16'h	d592;
26179	:douta	=	16'h	d591;
26180	:douta	=	16'h	ddf2;
26181	:douta	=	16'h	c531;
26182	:douta	=	16'h	c531;
26183	:douta	=	16'h	acb2;
26184	:douta	=	16'h	a4b2;
26185	:douta	=	16'h	a4b2;
26186	:douta	=	16'h	a4d3;
26187	:douta	=	16'h	9c93;
26188	:douta	=	16'h	8c32;
26189	:douta	=	16'h	7bd1;
26190	:douta	=	16'h	8412;
26191	:douta	=	16'h	73b0;
26192	:douta	=	16'h	734f;
26193	:douta	=	16'h	736f;
26194	:douta	=	16'h	6b4f;
26195	:douta	=	16'h	5aec;
26196	:douta	=	16'h	59e5;
26197	:douta	=	16'h	7266;
26198	:douta	=	16'h	ac2a;
26199	:douta	=	16'h	c4eb;
26200	:douta	=	16'h	e5d2;
26201	:douta	=	16'h	e653;
26202	:douta	=	16'h	e653;
26203	:douta	=	16'h	ee75;
26204	:douta	=	16'h	ee74;
26205	:douta	=	16'h	e653;
26206	:douta	=	16'h	e613;
26207	:douta	=	16'h	ee74;
26208	:douta	=	16'h	e633;
26209	:douta	=	16'h	e612;
26210	:douta	=	16'h	ddd1;
26211	:douta	=	16'h	cd50;
26212	:douta	=	16'h	c4f0;
26213	:douta	=	16'h	bcb0;
26214	:douta	=	16'h	b4b0;
26215	:douta	=	16'h	9c51;
26216	:douta	=	16'h	9452;
26217	:douta	=	16'h	8c12;
26218	:douta	=	16'h	8c73;
26219	:douta	=	16'h	8453;
26220	:douta	=	16'h	8c95;
26221	:douta	=	16'h	8455;
26222	:douta	=	16'h	73f3;
26223	:douta	=	16'h	73d2;
26224	:douta	=	16'h	7413;
26225	:douta	=	16'h	73f3;
26226	:douta	=	16'h	6bf3;
26227	:douta	=	16'h	5370;
26228	:douta	=	16'h	5b72;
26229	:douta	=	16'h	5330;
26230	:douta	=	16'h	4b10;
26231	:douta	=	16'h	4b31;
26232	:douta	=	16'h	31ea;
26233	:douta	=	16'h	4acf;
26234	:douta	=	16'h	42ae;
26235	:douta	=	16'h	0884;
26236	:douta	=	16'h	1926;
26237	:douta	=	16'h	29eb;
26238	:douta	=	16'h	0842;
26239	:douta	=	16'h	0862;
26240	:douta	=	16'h	1084;
26241	:douta	=	16'h	10a3;
26242	:douta	=	16'h	10a4;
26243	:douta	=	16'h	1905;
26244	:douta	=	16'h	1926;
26245	:douta	=	16'h	1905;
26246	:douta	=	16'h	1905;
26247	:douta	=	16'h	1926;
26248	:douta	=	16'h	1905;
26249	:douta	=	16'h	1946;
26250	:douta	=	16'h	0000;
26251	:douta	=	16'h	0000;
26252	:douta	=	16'h	0001;
26253	:douta	=	16'h	7cf9;
26254	:douta	=	16'h	84b7;
26255	:douta	=	16'h	0021;
26256	:douta	=	16'h	10e5;
26257	:douta	=	16'h	10e5;
26258	:douta	=	16'h	1106;
26259	:douta	=	16'h	31c8;
26260	:douta	=	16'h	8bed;
26261	:douta	=	16'h	9470;
26262	:douta	=	16'h	5248;
26263	:douta	=	16'h	946f;
26264	:douta	=	16'h	ad31;
26265	:douta	=	16'h	6b4b;
26266	:douta	=	16'h	83ce;
26267	:douta	=	16'h	3a2a;
26268	:douta	=	16'h	5b92;
26269	:douta	=	16'h	6c15;
26270	:douta	=	16'h	9dba;
26271	:douta	=	16'h	9d9a;
26272	:douta	=	16'h	8d17;
26273	:douta	=	16'h	84d7;
26274	:douta	=	16'h	8d18;
26275	:douta	=	16'h	84f8;
26276	:douta	=	16'h	8d59;
26277	:douta	=	16'h	9559;
26278	:douta	=	16'h	7cb7;
26279	:douta	=	16'h	7c97;
26280	:douta	=	16'h	8d39;
26281	:douta	=	16'h	8d18;
26282	:douta	=	16'h	9dbb;
26283	:douta	=	16'h	8d39;
26284	:douta	=	16'h	7476;
26285	:douta	=	16'h	84d7;
26286	:douta	=	16'h	84d7;
26287	:douta	=	16'h	7456;
26288	:douta	=	16'h	6c14;
26289	:douta	=	16'h	6c14;
26290	:douta	=	16'h	8d59;
26291	:douta	=	16'h	9dbb;
26292	:douta	=	16'h	84d8;
26293	:douta	=	16'h	8519;
26294	:douta	=	16'h	9d9a;
26295	:douta	=	16'h	9dba;
26296	:douta	=	16'h	9d9a;
26297	:douta	=	16'h	84f7;
26298	:douta	=	16'h	7497;
26299	:douta	=	16'h	6c15;
26300	:douta	=	16'h	5392;
26301	:douta	=	16'h	7cb7;
26302	:douta	=	16'h	8d39;
26303	:douta	=	16'h	8519;
26304	:douta	=	16'h	8518;
26305	:douta	=	16'h	957b;
26306	:douta	=	16'h	9dbb;
26307	:douta	=	16'h	959a;
26308	:douta	=	16'h	959a;
26309	:douta	=	16'h	8d5a;
26310	:douta	=	16'h	84f9;
26311	:douta	=	16'h	7cf9;
26312	:douta	=	16'h	8d39;
26313	:douta	=	16'h	957a;
26314	:douta	=	16'h	95dd;
26315	:douta	=	16'h	7476;
26316	:douta	=	16'h	5b92;
26317	:douta	=	16'h	5aed;
26318	:douta	=	16'h	5207;
26319	:douta	=	16'h	72a9;
26320	:douta	=	16'h	6248;
26321	:douta	=	16'h	6248;
26322	:douta	=	16'h	62ec;
26323	:douta	=	16'h	3a2c;
26324	:douta	=	16'h	224e;
26325	:douta	=	16'h	220c;
26326	:douta	=	16'h	2a6f;
26327	:douta	=	16'h	4c17;
26328	:douta	=	16'h	5438;
26329	:douta	=	16'h	4374;
26330	:douta	=	16'h	3b54;
26331	:douta	=	16'h	4b94;
26332	:douta	=	16'h	4bb4;
26333	:douta	=	16'h	4394;
26334	:douta	=	16'h	5c58;
26335	:douta	=	16'h	53b6;
26336	:douta	=	16'h	4b95;
26337	:douta	=	16'h	4b94;
26338	:douta	=	16'h	6457;
26339	:douta	=	16'h	53f6;
26340	:douta	=	16'h	53b6;
26341	:douta	=	16'h	4b95;
26342	:douta	=	16'h	3b33;
26343	:douta	=	16'h	5c17;
26344	:douta	=	16'h	6b0c;
26345	:douta	=	16'h	7b29;
26346	:douta	=	16'h	6a65;
26347	:douta	=	16'h	3144;
26348	:douta	=	16'h	20a2;
26349	:douta	=	16'h	0062;
26350	:douta	=	16'h	1926;
26351	:douta	=	16'h	5c58;
26352	:douta	=	16'h	649a;
26353	:douta	=	16'h	4af0;
26354	:douta	=	16'h	6bd0;
26355	:douta	=	16'h	bdd4;
26356	:douta	=	16'h	deb7;
26357	:douta	=	16'h	d657;
26358	:douta	=	16'h	ad52;
26359	:douta	=	16'h	5aa8;
26360	:douta	=	16'h	28c2;
26361	:douta	=	16'h	2881;
26362	:douta	=	16'h	3944;
26363	:douta	=	16'h	3964;
26364	:douta	=	16'h	4164;
26365	:douta	=	16'h	4185;
26366	:douta	=	16'h	3964;
26367	:douta	=	16'h	49a6;
26368	:douta	=	16'h	6390;
26369	:douta	=	16'h	3124;
26370	:douta	=	16'h	3986;
26371	:douta	=	16'h	3965;
26372	:douta	=	16'h	2904;
26373	:douta	=	16'h	1882;
26374	:douta	=	16'h	424b;
26375	:douta	=	16'h	2a4e;
26376	:douta	=	16'h	4353;
26377	:douta	=	16'h	4b95;
26378	:douta	=	16'h	4374;
26379	:douta	=	16'h	3ad1;
26380	:douta	=	16'h	6457;
26381	:douta	=	16'h	6c56;
26382	:douta	=	16'h	7476;
26383	:douta	=	16'h	6c15;
26384	:douta	=	16'h	63d3;
26385	:douta	=	16'h	73f3;
26386	:douta	=	16'h	8496;
26387	:douta	=	16'h	73f3;
26388	:douta	=	16'h	8c74;
26389	:douta	=	16'h	7c12;
26390	:douta	=	16'h	8433;
26391	:douta	=	16'h	ad77;
26392	:douta	=	16'h	c638;
26393	:douta	=	16'h	9d16;
26394	:douta	=	16'h	e613;
26395	:douta	=	16'h	ee95;
26396	:douta	=	16'h	e676;
26397	:douta	=	16'h	e696;
26398	:douta	=	16'h	e696;
26399	:douta	=	16'h	eed8;
26400	:douta	=	16'h	eed8;
26401	:douta	=	16'h	eed7;
26402	:douta	=	16'h	eed7;
26403	:douta	=	16'h	ee96;
26404	:douta	=	16'h	eeb7;
26405	:douta	=	16'h	ee96;
26406	:douta	=	16'h	e634;
26407	:douta	=	16'h	de13;
26408	:douta	=	16'h	d5b2;
26409	:douta	=	16'h	c551;
26410	:douta	=	16'h	bd31;
26411	:douta	=	16'h	8c10;
26412	:douta	=	16'h	7bd1;
26413	:douta	=	16'h	83f1;
26414	:douta	=	16'h	7bb0;
26415	:douta	=	16'h	7390;
26416	:douta	=	16'h	7bb0;
26417	:douta	=	16'h	734f;
26418	:douta	=	16'h	6b0d;
26419	:douta	=	16'h	4985;
26420	:douta	=	16'h	8328;
26421	:douta	=	16'h	ac4c;
26422	:douta	=	16'h	bcac;
26423	:douta	=	16'h	d570;
26424	:douta	=	16'h	e634;
26425	:douta	=	16'h	e675;
26426	:douta	=	16'h	ee75;
26427	:douta	=	16'h	e633;
26428	:douta	=	16'h	ddb1;
26429	:douta	=	16'h	ee75;
26430	:douta	=	16'h	e654;
26431	:douta	=	16'h	de13;
26432	:douta	=	16'h	d5b1;
26433	:douta	=	16'h	d591;
26434	:douta	=	16'h	cd71;
26435	:douta	=	16'h	c530;
26436	:douta	=	16'h	bd11;
26437	:douta	=	16'h	c531;
26438	:douta	=	16'h	b4f1;
26439	:douta	=	16'h	a4b2;
26440	:douta	=	16'h	a4b2;
26441	:douta	=	16'h	9453;
26442	:douta	=	16'h	8c12;
26443	:douta	=	16'h	9472;
26444	:douta	=	16'h	8412;
26445	:douta	=	16'h	83f1;
26446	:douta	=	16'h	732e;
26447	:douta	=	16'h	7bb0;
26448	:douta	=	16'h	7bb0;
26449	:douta	=	16'h	734f;
26450	:douta	=	16'h	4a28;
26451	:douta	=	16'h	7a87;
26452	:douta	=	16'h	9b8a;
26453	:douta	=	16'h	a3ca;
26454	:douta	=	16'h	cd2d;
26455	:douta	=	16'h	ddd1;
26456	:douta	=	16'h	e654;
26457	:douta	=	16'h	e654;
26458	:douta	=	16'h	ee74;
26459	:douta	=	16'h	ee74;
26460	:douta	=	16'h	ee74;
26461	:douta	=	16'h	ee54;
26462	:douta	=	16'h	e653;
26463	:douta	=	16'h	e632;
26464	:douta	=	16'h	ddd0;
26465	:douta	=	16'h	ddb0;
26466	:douta	=	16'h	cd30;
26467	:douta	=	16'h	bd0f;
26468	:douta	=	16'h	b48f;
26469	:douta	=	16'h	a450;
26470	:douta	=	16'h	a470;
26471	:douta	=	16'h	9451;
26472	:douta	=	16'h	8c11;
26473	:douta	=	16'h	9432;
26474	:douta	=	16'h	8c32;
26475	:douta	=	16'h	8c94;
26476	:douta	=	16'h	8454;
26477	:douta	=	16'h	8474;
26478	:douta	=	16'h	8474;
26479	:douta	=	16'h	8475;
26480	:douta	=	16'h	7c13;
26481	:douta	=	16'h	7413;
26482	:douta	=	16'h	73f3;
26483	:douta	=	16'h	63b2;
26484	:douta	=	16'h	5b50;
26485	:douta	=	16'h	5b30;
26486	:douta	=	16'h	3a2c;
26487	:douta	=	16'h	7b2d;
26488	:douta	=	16'h	4ace;
26489	:douta	=	16'h	428d;
26490	:douta	=	16'h	4ace;
26491	:douta	=	16'h	3a8d;
26492	:douta	=	16'h	2167;
26493	:douta	=	16'h	10c4;
26494	:douta	=	16'h	428d;
26495	:douta	=	16'h	4acf;
26496	:douta	=	16'h	0883;
26497	:douta	=	16'h	0863;
26498	:douta	=	16'h	10c4;
26499	:douta	=	16'h	18e5;
26500	:douta	=	16'h	10e5;
26501	:douta	=	16'h	10e4;
26502	:douta	=	16'h	10c4;
26503	:douta	=	16'h	10c4;
26504	:douta	=	16'h	10e5;
26505	:douta	=	16'h	10e5;
26506	:douta	=	16'h	1926;
26507	:douta	=	16'h	1926;
26508	:douta	=	16'h	0000;
26509	:douta	=	16'h	0000;
26510	:douta	=	16'h	0000;
26511	:douta	=	16'h	1905;
26512	:douta	=	16'h	2126;
26513	:douta	=	16'h	2147;
26514	:douta	=	16'h	1946;
26515	:douta	=	16'h	1926;
26516	:douta	=	16'h	3a08;
26517	:douta	=	16'h	5aec;
26518	:douta	=	16'h	bd51;
26519	:douta	=	16'h	ad11;
26520	:douta	=	16'h	7bad;
26521	:douta	=	16'h	a4b0;
26522	:douta	=	16'h	4248;
26523	:douta	=	16'h	62eb;
26524	:douta	=	16'h	9c8f;
26525	:douta	=	16'h	7b8c;
26526	:douta	=	16'h	6b0b;
26527	:douta	=	16'h	4208;
26528	:douta	=	16'h	428d;
26529	:douta	=	16'h	530e;
26530	:douta	=	16'h	5b51;
26531	:douta	=	16'h	7476;
26532	:douta	=	16'h	9559;
26533	:douta	=	16'h	8d59;
26534	:douta	=	16'h	8d39;
26535	:douta	=	16'h	8d18;
26536	:douta	=	16'h	8cf8;
26537	:douta	=	16'h	8518;
26538	:douta	=	16'h	8d39;
26539	:douta	=	16'h	9559;
26540	:douta	=	16'h	8d18;
26541	:douta	=	16'h	84d7;
26542	:douta	=	16'h	7cb7;
26543	:douta	=	16'h	8d39;
26544	:douta	=	16'h	9dbb;
26545	:douta	=	16'h	84f8;
26546	:douta	=	16'h	7cb7;
26547	:douta	=	16'h	6c76;
26548	:douta	=	16'h	959a;
26549	:douta	=	16'h	8518;
26550	:douta	=	16'h	7cb7;
26551	:douta	=	16'h	8d39;
26552	:douta	=	16'h	8d39;
26553	:douta	=	16'h	84f8;
26554	:douta	=	16'h	9559;
26555	:douta	=	16'h	84f8;
26556	:douta	=	16'h	9ddc;
26557	:douta	=	16'h	957a;
26558	:douta	=	16'h	6435;
26559	:douta	=	16'h	5371;
26560	:douta	=	16'h	5b52;
26561	:douta	=	16'h	74b6;
26562	:douta	=	16'h	7cf8;
26563	:douta	=	16'h	8539;
26564	:douta	=	16'h	74b7;
26565	:douta	=	16'h	8d59;
26566	:douta	=	16'h	7cb7;
26567	:douta	=	16'h	7496;
26568	:douta	=	16'h	63b3;
26569	:douta	=	16'h	42cf;
26570	:douta	=	16'h	3a2d;
26571	:douta	=	16'h	4310;
26572	:douta	=	16'h	5bb4;
26573	:douta	=	16'h	42d0;
26574	:douta	=	16'h	4b11;
26575	:douta	=	16'h	62ed;
26576	:douta	=	16'h	72a8;
26577	:douta	=	16'h	72a9;
26578	:douta	=	16'h	6248;
26579	:douta	=	16'h	6248;
26580	:douta	=	16'h	5a8a;
26581	:douta	=	16'h	3ad0;
26582	:douta	=	16'h	11cd;
26583	:douta	=	16'h	4395;
26584	:douta	=	16'h	2ab0;
26585	:douta	=	16'h	3b95;
26586	:douta	=	16'h	43d6;
26587	:douta	=	16'h	3b33;
26588	:douta	=	16'h	4bd6;
26589	:douta	=	16'h	3b74;
26590	:douta	=	16'h	4bb5;
26591	:douta	=	16'h	4374;
26592	:douta	=	16'h	4b75;
26593	:douta	=	16'h	6cba;
26594	:douta	=	16'h	6458;
26595	:douta	=	16'h	53d6;
26596	:douta	=	16'h	6479;
26597	:douta	=	16'h	4334;
26598	:douta	=	16'h	7d7c;
26599	:douta	=	16'h	5c37;
26600	:douta	=	16'h	5c78;
26601	:douta	=	16'h	8b26;
26602	:douta	=	16'h	8348;
26603	:douta	=	16'h	51c4;
26604	:douta	=	16'h	3144;
26605	:douta	=	16'h	0882;
26606	:douta	=	16'h	0000;
26607	:douta	=	16'h	08e5;
26608	:douta	=	16'h	94d3;
26609	:douta	=	16'h	b593;
26610	:douta	=	16'h	de75;
26611	:douta	=	16'h	ad10;
26612	:douta	=	16'h	6b4a;
26613	:douta	=	16'h	3964;
26614	:douta	=	16'h	30c2;
26615	:douta	=	16'h	3944;
26616	:douta	=	16'h	3944;
26617	:douta	=	16'h	4164;
26618	:douta	=	16'h	4185;
26619	:douta	=	16'h	41a5;
26620	:douta	=	16'h	4985;
26621	:douta	=	16'h	3985;
26622	:douta	=	16'h	41a5;
26623	:douta	=	16'h	49c7;
26624	:douta	=	16'h	5b0e;
26625	:douta	=	16'h	3924;
26626	:douta	=	16'h	3966;
26627	:douta	=	16'h	3945;
26628	:douta	=	16'h	2904;
26629	:douta	=	16'h	18a3;
26630	:douta	=	16'h	4a6c;
26631	:douta	=	16'h	21ca;
26632	:douta	=	16'h	4b95;
26633	:douta	=	16'h	3b53;
26634	:douta	=	16'h	53d6;
26635	:douta	=	16'h	4333;
26636	:douta	=	16'h	5c16;
26637	:douta	=	16'h	74b8;
26638	:douta	=	16'h	7455;
26639	:douta	=	16'h	7c97;
26640	:douta	=	16'h	6bf4;
26641	:douta	=	16'h	73f4;
26642	:douta	=	16'h	7c75;
26643	:douta	=	16'h	73f4;
26644	:douta	=	16'h	94b5;
26645	:douta	=	16'h	8c74;
26646	:douta	=	16'h	8c74;
26647	:douta	=	16'h	bdd8;
26648	:douta	=	16'h	c618;
26649	:douta	=	16'h	ad97;
26650	:douta	=	16'h	bd13;
26651	:douta	=	16'h	ee94;
26652	:douta	=	16'h	e696;
26653	:douta	=	16'h	eeb7;
26654	:douta	=	16'h	e696;
26655	:douta	=	16'h	eed8;
26656	:douta	=	16'h	eed8;
26657	:douta	=	16'h	eeb7;
26658	:douta	=	16'h	eeb7;
26659	:douta	=	16'h	eeb7;
26660	:douta	=	16'h	ee96;
26661	:douta	=	16'h	e696;
26662	:douta	=	16'h	e634;
26663	:douta	=	16'h	d5f3;
26664	:douta	=	16'h	cdb2;
26665	:douta	=	16'h	b4d2;
26666	:douta	=	16'h	a4b1;
26667	:douta	=	16'h	9c71;
26668	:douta	=	16'h	83f1;
26669	:douta	=	16'h	7bd1;
26670	:douta	=	16'h	738f;
26671	:douta	=	16'h	736f;
26672	:douta	=	16'h	6b4e;
26673	:douta	=	16'h	630c;
26674	:douta	=	16'h	41c7;
26675	:douta	=	16'h	8b29;
26676	:douta	=	16'h	b48c;
26677	:douta	=	16'h	a44c;
26678	:douta	=	16'h	cd2e;
26679	:douta	=	16'h	de12;
26680	:douta	=	16'h	e675;
26681	:douta	=	16'h	ee96;
26682	:douta	=	16'h	e675;
26683	:douta	=	16'h	e695;
26684	:douta	=	16'h	e612;
26685	:douta	=	16'h	e633;
26686	:douta	=	16'h	e674;
26687	:douta	=	16'h	ddb1;
26688	:douta	=	16'h	d591;
26689	:douta	=	16'h	cd51;
26690	:douta	=	16'h	cd50;
26691	:douta	=	16'h	c530;
26692	:douta	=	16'h	acb1;
26693	:douta	=	16'h	bcf1;
26694	:douta	=	16'h	b4d2;
26695	:douta	=	16'h	acb2;
26696	:douta	=	16'h	a493;
26697	:douta	=	16'h	8c32;
26698	:douta	=	16'h	8c12;
26699	:douta	=	16'h	8c11;
26700	:douta	=	16'h	8c12;
26701	:douta	=	16'h	83d1;
26702	:douta	=	16'h	734e;
26703	:douta	=	16'h	730e;
26704	:douta	=	16'h	6b6f;
26705	:douta	=	16'h	49a5;
26706	:douta	=	16'h	4963;
26707	:douta	=	16'h	abeb;
26708	:douta	=	16'h	ac4a;
26709	:douta	=	16'h	bcac;
26710	:douta	=	16'h	dd8f;
26711	:douta	=	16'h	e653;
26712	:douta	=	16'h	ee95;
26713	:douta	=	16'h	ee75;
26714	:douta	=	16'h	e674;
26715	:douta	=	16'h	ee54;
26716	:douta	=	16'h	ee74;
26717	:douta	=	16'h	ee54;
26718	:douta	=	16'h	e653;
26719	:douta	=	16'h	ddf2;
26720	:douta	=	16'h	d58f;
26721	:douta	=	16'h	cd4f;
26722	:douta	=	16'h	bccf;
26723	:douta	=	16'h	b4af;
26724	:douta	=	16'h	a430;
26725	:douta	=	16'h	9c51;
26726	:douta	=	16'h	9c51;
26727	:douta	=	16'h	9452;
26728	:douta	=	16'h	8c32;
26729	:douta	=	16'h	9452;
26730	:douta	=	16'h	8c33;
26731	:douta	=	16'h	8432;
26732	:douta	=	16'h	8453;
26733	:douta	=	16'h	8433;
26734	:douta	=	16'h	8453;
26735	:douta	=	16'h	7bf3;
26736	:douta	=	16'h	7c13;
26737	:douta	=	16'h	7c33;
26738	:douta	=	16'h	6bd2;
26739	:douta	=	16'h	5b0e;
26740	:douta	=	16'h	52ae;
26741	:douta	=	16'h	4a2a;
26742	:douta	=	16'h	9329;
26743	:douta	=	16'h	e5b2;
26744	:douta	=	16'h	5351;
26745	:douta	=	16'h	3a6c;
26746	:douta	=	16'h	4ace;
26747	:douta	=	16'h	3aad;
26748	:douta	=	16'h	1948;
26749	:douta	=	16'h	18e5;
26750	:douta	=	16'h	0884;
26751	:douta	=	16'h	2989;
26752	:douta	=	16'h	4aae;
26753	:douta	=	16'h	29e9;
26754	:douta	=	16'h	0883;
26755	:douta	=	16'h	10e5;
26756	:douta	=	16'h	10e5;
26757	:douta	=	16'h	10e5;
26758	:douta	=	16'h	10e5;
26759	:douta	=	16'h	10e5;
26760	:douta	=	16'h	10e5;
26761	:douta	=	16'h	10e5;
26762	:douta	=	16'h	10e5;
26763	:douta	=	16'h	1906;
26764	:douta	=	16'h	10c4;
26765	:douta	=	16'h	0842;
26766	:douta	=	16'h	0000;
26767	:douta	=	16'h	0042;
26768	:douta	=	16'h	0883;
26769	:douta	=	16'h	1926;
26770	:douta	=	16'h	2167;
26771	:douta	=	16'h	1947;
26772	:douta	=	16'h	08a5;
26773	:douta	=	16'h	29aa;
26774	:douta	=	16'h	738e;
26775	:douta	=	16'h	732b;
26776	:douta	=	16'h	3186;
26777	:douta	=	16'h	ad11;
26778	:douta	=	16'h	b512;
26779	:douta	=	16'h	2124;
26780	:douta	=	16'h	a4b0;
26781	:douta	=	16'h	5289;
26782	:douta	=	16'h	5aa9;
26783	:douta	=	16'h	41e8;
26784	:douta	=	16'h	8bcd;
26785	:douta	=	16'h	3166;
26786	:douta	=	16'h	4207;
26787	:douta	=	16'h	528b;
26788	:douta	=	16'h	5aed;
26789	:douta	=	16'h	5310;
26790	:douta	=	16'h	5b92;
26791	:douta	=	16'h	7476;
26792	:douta	=	16'h	7cd7;
26793	:douta	=	16'h	8518;
26794	:douta	=	16'h	959a;
26795	:douta	=	16'h	8d39;
26796	:douta	=	16'h	9559;
26797	:douta	=	16'h	8d39;
26798	:douta	=	16'h	957a;
26799	:douta	=	16'h	8518;
26800	:douta	=	16'h	8518;
26801	:douta	=	16'h	8d39;
26802	:douta	=	16'h	84d7;
26803	:douta	=	16'h	8538;
26804	:douta	=	16'h	8d18;
26805	:douta	=	16'h	8d39;
26806	:douta	=	16'h	8d59;
26807	:douta	=	16'h	7cd7;
26808	:douta	=	16'h	8d18;
26809	:douta	=	16'h	9dbb;
26810	:douta	=	16'h	8519;
26811	:douta	=	16'h	9dfc;
26812	:douta	=	16'h	a63d;
26813	:douta	=	16'h	9dfc;
26814	:douta	=	16'h	ae7e;
26815	:douta	=	16'h	a65e;
26816	:douta	=	16'h	4b73;
26817	:douta	=	16'h	08c5;
26818	:douta	=	16'h	10e6;
26819	:douta	=	16'h	634f;
26820	:douta	=	16'h	3a2b;
26821	:douta	=	16'h	322b;
26822	:douta	=	16'h	3a4c;
26823	:douta	=	16'h	2189;
26824	:douta	=	16'h	29ca;
26825	:douta	=	16'h	324d;
26826	:douta	=	16'h	4b51;
26827	:douta	=	16'h	3a8e;
26828	:douta	=	16'h	3aaf;
26829	:douta	=	16'h	5352;
26830	:douta	=	16'h	4b51;
26831	:douta	=	16'h	5bb3;
26832	:douta	=	16'h	734d;
26833	:douta	=	16'h	72a9;
26834	:douta	=	16'h	6aa9;
26835	:douta	=	16'h	6a89;
26836	:douta	=	16'h	6248;
26837	:douta	=	16'h	6b0d;
26838	:douta	=	16'h	320b;
26839	:douta	=	16'h	118a;
26840	:douta	=	16'h	21ed;
26841	:douta	=	16'h	4c59;
26842	:douta	=	16'h	3333;
26843	:douta	=	16'h	32d2;
26844	:douta	=	16'h	2af2;
26845	:douta	=	16'h	3b53;
26846	:douta	=	16'h	3b12;
26847	:douta	=	16'h	4bb5;
26848	:douta	=	16'h	5417;
26849	:douta	=	16'h	4bb5;
26850	:douta	=	16'h	5c17;
26851	:douta	=	16'h	6cb9;
26852	:douta	=	16'h	4374;
26853	:douta	=	16'h	53b4;
26854	:douta	=	16'h	7d7c;
26855	:douta	=	16'h	53f6;
26856	:douta	=	16'h	7dbf;
26857	:douta	=	16'h	82e6;
26858	:douta	=	16'h	8b69;
26859	:douta	=	16'h	6245;
26860	:douta	=	16'h	4164;
26861	:douta	=	16'h	0001;
26862	:douta	=	16'h	2146;
26863	:douta	=	16'h	73ef;
26864	:douta	=	16'h	ce13;
26865	:douta	=	16'h	e697;
26866	:douta	=	16'h	ad2e;
26867	:douta	=	16'h	41a6;
26868	:douta	=	16'h	3923;
26869	:douta	=	16'h	28e2;
26870	:douta	=	16'h	3944;
26871	:douta	=	16'h	41a5;
26872	:douta	=	16'h	4185;
26873	:douta	=	16'h	4185;
26874	:douta	=	16'h	49a6;
26875	:douta	=	16'h	49a6;
26876	:douta	=	16'h	41a6;
26877	:douta	=	16'h	41a6;
26878	:douta	=	16'h	41a7;
26879	:douta	=	16'h	4186;
26880	:douta	=	16'h	41a7;
26881	:douta	=	16'h	4a8b;
26882	:douta	=	16'h	3924;
26883	:douta	=	16'h	3965;
26884	:douta	=	16'h	2924;
26885	:douta	=	16'h	20e3;
26886	:douta	=	16'h	426d;
26887	:douta	=	16'h	29aa;
26888	:douta	=	16'h	320d;
26889	:douta	=	16'h	4b94;
26890	:douta	=	16'h	3af1;
26891	:douta	=	16'h	4354;
26892	:douta	=	16'h	2a6f;
26893	:douta	=	16'h	7cd9;
26894	:douta	=	16'h	63d4;
26895	:douta	=	16'h	5bb3;
26896	:douta	=	16'h	84f8;
26897	:douta	=	16'h	6c35;
26898	:douta	=	16'h	8496;
26899	:douta	=	16'h	8cf6;
26900	:douta	=	16'h	7c13;
26901	:douta	=	16'h	9d16;
26902	:douta	=	16'h	7c33;
26903	:douta	=	16'h	b576;
26904	:douta	=	16'h	b5b8;
26905	:douta	=	16'h	b5b8;
26906	:douta	=	16'h	9474;
26907	:douta	=	16'h	a4b2;
26908	:douta	=	16'h	eeb5;
26909	:douta	=	16'h	e696;
26910	:douta	=	16'h	eeb7;
26911	:douta	=	16'h	eeb7;
26912	:douta	=	16'h	eed7;
26913	:douta	=	16'h	eed7;
26914	:douta	=	16'h	eeb6;
26915	:douta	=	16'h	e675;
26916	:douta	=	16'h	e675;
26917	:douta	=	16'h	de55;
26918	:douta	=	16'h	ddf4;
26919	:douta	=	16'h	cd72;
26920	:douta	=	16'h	bd11;
26921	:douta	=	16'h	a491;
26922	:douta	=	16'h	9c71;
26923	:douta	=	16'h	8c11;
26924	:douta	=	16'h	7bd1;
26925	:douta	=	16'h	7bb0;
26926	:douta	=	16'h	734e;
26927	:douta	=	16'h	6b2e;
26928	:douta	=	16'h	5aab;
26929	:douta	=	16'h	49a4;
26930	:douta	=	16'h	9369;
26931	:douta	=	16'h	ac4c;
26932	:douta	=	16'h	bcce;
26933	:douta	=	16'h	cd2f;
26934	:douta	=	16'h	ee95;
26935	:douta	=	16'h	e675;
26936	:douta	=	16'h	ee96;
26937	:douta	=	16'h	eeb7;
26938	:douta	=	16'h	ee95;
26939	:douta	=	16'h	e633;
26940	:douta	=	16'h	ddf2;
26941	:douta	=	16'h	d590;
26942	:douta	=	16'h	d591;
26943	:douta	=	16'h	cd50;
26944	:douta	=	16'h	c510;
26945	:douta	=	16'h	c511;
26946	:douta	=	16'h	b4b0;
26947	:douta	=	16'h	b4b1;
26948	:douta	=	16'h	acb1;
26949	:douta	=	16'h	a492;
26950	:douta	=	16'h	9452;
26951	:douta	=	16'h	9432;
26952	:douta	=	16'h	9452;
26953	:douta	=	16'h	8c11;
26954	:douta	=	16'h	6b4e;
26955	:douta	=	16'h	6b4e;
26956	:douta	=	16'h	734e;
26957	:douta	=	16'h	7b6f;
26958	:douta	=	16'h	83f1;
26959	:douta	=	16'h	41a7;
26960	:douta	=	16'h	4124;
26961	:douta	=	16'h	9bca;
26962	:douta	=	16'h	b42c;
26963	:douta	=	16'h	c4cd;
26964	:douta	=	16'h	e612;
26965	:douta	=	16'h	eeb5;
26966	:douta	=	16'h	f6d7;
26967	:douta	=	16'h	f6d7;
26968	:douta	=	16'h	eeb6;
26969	:douta	=	16'h	f6b6;
26970	:douta	=	16'h	ee74;
26971	:douta	=	16'h	ee95;
26972	:douta	=	16'h	e653;
26973	:douta	=	16'h	e613;
26974	:douta	=	16'h	e613;
26975	:douta	=	16'h	d570;
26976	:douta	=	16'h	cd10;
26977	:douta	=	16'h	c4f1;
26978	:douta	=	16'h	ac70;
26979	:douta	=	16'h	a471;
26980	:douta	=	16'h	9c51;
26981	:douta	=	16'h	9c52;
26982	:douta	=	16'h	9c52;
26983	:douta	=	16'h	9c72;
26984	:douta	=	16'h	9432;
26985	:douta	=	16'h	8c12;
26986	:douta	=	16'h	8c32;
26987	:douta	=	16'h	8412;
26988	:douta	=	16'h	7bd1;
26989	:douta	=	16'h	7bb1;
26990	:douta	=	16'h	7bd2;
26991	:douta	=	16'h	7bf2;
26992	:douta	=	16'h	7b90;
26993	:douta	=	16'h	6b0d;
26994	:douta	=	16'h	62cd;
26995	:douta	=	16'h	5a49;
26996	:douta	=	16'h	b42a;
26997	:douta	=	16'h	ddaf;
26998	:douta	=	16'h	f6b7;
26999	:douta	=	16'h	d592;
27000	:douta	=	16'h	7c53;
27001	:douta	=	16'h	5b50;
27002	:douta	=	16'h	5b4f;
27003	:douta	=	16'h	6391;
27004	:douta	=	16'h	42cf;
27005	:douta	=	16'h	29ea;
27006	:douta	=	16'h	2168;
27007	:douta	=	16'h	2148;
27008	:douta	=	16'h	0884;
27009	:douta	=	16'h	10e5;
27010	:douta	=	16'h	4aae;
27011	:douta	=	16'h	320a;
27012	:douta	=	16'h	10a4;
27013	:douta	=	16'h	10c5;
27014	:douta	=	16'h	18e5;
27015	:douta	=	16'h	18e5;
27016	:douta	=	16'h	1905;
27017	:douta	=	16'h	1905;
27018	:douta	=	16'h	1905;
27019	:douta	=	16'h	18e5;
27020	:douta	=	16'h	10a4;
27021	:douta	=	16'h	10c4;
27022	:douta	=	16'h	1906;
27023	:douta	=	16'h	10e5;
27024	:douta	=	16'h	10c5;
27025	:douta	=	16'h	0021;
27026	:douta	=	16'h	0021;
27027	:douta	=	16'h	0884;
27028	:douta	=	16'h	2967;
27029	:douta	=	16'h	4229;
27030	:douta	=	16'h	4aef;
27031	:douta	=	16'h	4b52;
27032	:douta	=	16'h	7c54;
27033	:douta	=	16'h	2988;
27034	:douta	=	16'h	10a4;
27035	:douta	=	16'h	83ed;
27036	:douta	=	16'h	9c6e;
27037	:douta	=	16'h	83cd;
27038	:douta	=	16'h	62cb;
27039	:douta	=	16'h	83ef;
27040	:douta	=	16'h	944e;
27041	:douta	=	16'h	9c4f;
27042	:douta	=	16'h	a4b1;
27043	:douta	=	16'h	39e8;
27044	:douta	=	16'h	2946;
27045	:douta	=	16'h	ad32;
27046	:douta	=	16'h	6b4b;
27047	:douta	=	16'h	4a28;
27048	:douta	=	16'h	7b6c;
27049	:douta	=	16'h	528a;
27050	:douta	=	16'h	0884;
27051	:douta	=	16'h	29a8;
27052	:douta	=	16'h	526b;
27053	:douta	=	16'h	428c;
27054	:douta	=	16'h	426b;
27055	:douta	=	16'h	4a8c;
27056	:douta	=	16'h	4aee;
27057	:douta	=	16'h	4aae;
27058	:douta	=	16'h	5b70;
27059	:douta	=	16'h	5b2f;
27060	:douta	=	16'h	5b70;
27061	:douta	=	16'h	4aad;
27062	:douta	=	16'h	5b0f;
27063	:douta	=	16'h	52ef;
27064	:douta	=	16'h	4aad;
27065	:douta	=	16'h	31ea;
27066	:douta	=	16'h	31e9;
27067	:douta	=	16'h	18c5;
27068	:douta	=	16'h	6b2c;
27069	:douta	=	16'h	7b2b;
27070	:douta	=	16'h	7aa6;
27071	:douta	=	16'h	82e6;
27072	:douta	=	16'h	9bca;
27073	:douta	=	16'h	b42c;
27074	:douta	=	16'h	836c;
27075	:douta	=	16'h	1968;
27076	:douta	=	16'h	29eb;
27077	:douta	=	16'h	4aee;
27078	:douta	=	16'h	29ca;
27079	:douta	=	16'h	3a8d;
27080	:douta	=	16'h	324b;
27081	:douta	=	16'h	2a0b;
27082	:douta	=	16'h	2a0b;
27083	:douta	=	16'h	4310;
27084	:douta	=	16'h	3af1;
27085	:douta	=	16'h	63f3;
27086	:douta	=	16'h	6c14;
27087	:douta	=	16'h	5bd3;
27088	:douta	=	16'h	3acf;
27089	:douta	=	16'h	5372;
27090	:douta	=	16'h	52cd;
27091	:douta	=	16'h	6269;
27092	:douta	=	16'h	6a89;
27093	:douta	=	16'h	5a49;
27094	:douta	=	16'h	5a48;
27095	:douta	=	16'h	62aa;
27096	:douta	=	16'h	52ef;
27097	:douta	=	16'h	098c;
27098	:douta	=	16'h	2ab0;
27099	:douta	=	16'h	3b54;
27100	:douta	=	16'h	3313;
27101	:douta	=	16'h	32d1;
27102	:douta	=	16'h	3b54;
27103	:douta	=	16'h	32d1;
27104	:douta	=	16'h	2ad1;
27105	:douta	=	16'h	4373;
27106	:douta	=	16'h	5c58;
27107	:douta	=	16'h	3b53;
27108	:douta	=	16'h	4b95;
27109	:douta	=	16'h	6498;
27110	:douta	=	16'h	5c58;
27111	:douta	=	16'h	7d9c;
27112	:douta	=	16'h	3b12;
27113	:douta	=	16'h	5351;
27114	:douta	=	16'h	7ac6;
27115	:douta	=	16'h	8307;
27116	:douta	=	16'h	59e5;
27117	:douta	=	16'h	94d1;
27118	:douta	=	16'h	c5f3;
27119	:douta	=	16'h	bd71;
27120	:douta	=	16'h	5205;
27121	:douta	=	16'h	30e2;
27122	:douta	=	16'h	30c2;
27123	:douta	=	16'h	3964;
27124	:douta	=	16'h	3944;
27125	:douta	=	16'h	41a5;
27126	:douta	=	16'h	4185;
27127	:douta	=	16'h	41a5;
27128	:douta	=	16'h	41a6;
27129	:douta	=	16'h	41a6;
27130	:douta	=	16'h	41a6;
27131	:douta	=	16'h	4186;
27132	:douta	=	16'h	41a7;
27133	:douta	=	16'h	41a7;
27134	:douta	=	16'h	49c7;
27135	:douta	=	16'h	41c7;
27136	:douta	=	16'h	4144;
27137	:douta	=	16'h	5b4f;
27138	:douta	=	16'h	3904;
27139	:douta	=	16'h	3965;
27140	:douta	=	16'h	2924;
27141	:douta	=	16'h	2904;
27142	:douta	=	16'h	4a8d;
27143	:douta	=	16'h	42ce;
27144	:douta	=	16'h	2168;
27145	:douta	=	16'h	4334;
27146	:douta	=	16'h	19eb;
27147	:douta	=	16'h	220d;
27148	:douta	=	16'h	4353;
27149	:douta	=	16'h	5372;
27150	:douta	=	16'h	6c36;
27151	:douta	=	16'h	6c15;
27152	:douta	=	16'h	7cd8;
27153	:douta	=	16'h	7c96;
27154	:douta	=	16'h	7414;
27155	:douta	=	16'h	8cd7;
27156	:douta	=	16'h	94f6;
27157	:douta	=	16'h	a536;
27158	:douta	=	16'h	b597;
27159	:douta	=	16'h	9cd5;
27160	:douta	=	16'h	c5f8;
27161	:douta	=	16'h	c639;
27162	:douta	=	16'h	9492;
27163	:douta	=	16'h	7bf1;
27164	:douta	=	16'h	e614;
27165	:douta	=	16'h	e696;
27166	:douta	=	16'h	e6b7;
27167	:douta	=	16'h	eeb7;
27168	:douta	=	16'h	eed7;
27169	:douta	=	16'h	eed7;
27170	:douta	=	16'h	ee96;
27171	:douta	=	16'h	e675;
27172	:douta	=	16'h	e675;
27173	:douta	=	16'h	e654;
27174	:douta	=	16'h	d5d3;
27175	:douta	=	16'h	c571;
27176	:douta	=	16'h	b4f1;
27177	:douta	=	16'h	9c51;
27178	:douta	=	16'h	8c31;
27179	:douta	=	16'h	8c11;
27180	:douta	=	16'h	83f1;
27181	:douta	=	16'h	7b90;
27182	:douta	=	16'h	6b0e;
27183	:douta	=	16'h	62ed;
27184	:douta	=	16'h	3945;
27185	:douta	=	16'h	9baa;
27186	:douta	=	16'h	a46c;
27187	:douta	=	16'h	ac6c;
27188	:douta	=	16'h	bcee;
27189	:douta	=	16'h	ddd2;
27190	:douta	=	16'h	e655;
27191	:douta	=	16'h	e634;
27192	:douta	=	16'h	ee96;
27193	:douta	=	16'h	eeb7;
27194	:douta	=	16'h	e695;
27195	:douta	=	16'h	e655;
27196	:douta	=	16'h	bcef;
27197	:douta	=	16'h	e5f2;
27198	:douta	=	16'h	d550;
27199	:douta	=	16'h	cd50;
27200	:douta	=	16'h	bcd1;
27201	:douta	=	16'h	b4d1;
27202	:douta	=	16'h	acd1;
27203	:douta	=	16'h	a4b1;
27204	:douta	=	16'h	a471;
27205	:douta	=	16'h	a471;
27206	:douta	=	16'h	9452;
27207	:douta	=	16'h	83f1;
27208	:douta	=	16'h	7bd1;
27209	:douta	=	16'h	83d1;
27210	:douta	=	16'h	738f;
27211	:douta	=	16'h	734f;
27212	:douta	=	16'h	6b2d;
27213	:douta	=	16'h	732e;
27214	:douta	=	16'h	62cd;
27215	:douta	=	16'h	4985;
27216	:douta	=	16'h	82e9;
27217	:douta	=	16'h	ac2c;
27218	:douta	=	16'h	b48b;
27219	:douta	=	16'h	d54f;
27220	:douta	=	16'h	eeb6;
27221	:douta	=	16'h	eeb6;
27222	:douta	=	16'h	eeb7;
27223	:douta	=	16'h	eeb7;
27224	:douta	=	16'h	ee95;
27225	:douta	=	16'h	ee95;
27226	:douta	=	16'h	ee74;
27227	:douta	=	16'h	e654;
27228	:douta	=	16'h	e653;
27229	:douta	=	16'h	ddd2;
27230	:douta	=	16'h	ddb1;
27231	:douta	=	16'h	d530;
27232	:douta	=	16'h	b4d0;
27233	:douta	=	16'h	b4d1;
27234	:douta	=	16'h	a472;
27235	:douta	=	16'h	9c71;
27236	:douta	=	16'h	9c52;
27237	:douta	=	16'h	9452;
27238	:douta	=	16'h	9452;
27239	:douta	=	16'h	9432;
27240	:douta	=	16'h	8c32;
27241	:douta	=	16'h	83f1;
27242	:douta	=	16'h	7bd0;
27243	:douta	=	16'h	738f;
27244	:douta	=	16'h	7b90;
27245	:douta	=	16'h	7bb0;
27246	:douta	=	16'h	73b0;
27247	:douta	=	16'h	734f;
27248	:douta	=	16'h	734f;
27249	:douta	=	16'h	62ec;
27250	:douta	=	16'h	5a6b;
27251	:douta	=	16'h	7a87;
27252	:douta	=	16'h	ddd1;
27253	:douta	=	16'h	cd4e;
27254	:douta	=	16'h	d5d2;
27255	:douta	=	16'h	e614;
27256	:douta	=	16'h	9472;
27257	:douta	=	16'h	6391;
27258	:douta	=	16'h	6b90;
27259	:douta	=	16'h	73f2;
27260	:douta	=	16'h	5b71;
27261	:douta	=	16'h	42ae;
27262	:douta	=	16'h	29cb;
27263	:douta	=	16'h	29eb;
27264	:douta	=	16'h	2147;
27265	:douta	=	16'h	2147;
27266	:douta	=	16'h	0884;
27267	:douta	=	16'h	3a6d;
27268	:douta	=	16'h	326d;
27269	:douta	=	16'h	10a4;
27270	:douta	=	16'h	1083;
27271	:douta	=	16'h	18c5;
27272	:douta	=	16'h	1905;
27273	:douta	=	16'h	1905;
27274	:douta	=	16'h	1926;
27275	:douta	=	16'h	1926;
27276	:douta	=	16'h	18e5;
27277	:douta	=	16'h	10e4;
27278	:douta	=	16'h	1926;
27279	:douta	=	16'h	2127;
27280	:douta	=	16'h	2146;
27281	:douta	=	16'h	08a4;
27282	:douta	=	16'h	0042;
27283	:douta	=	16'h	0001;
27284	:douta	=	16'h	0001;
27285	:douta	=	16'h	1063;
27286	:douta	=	16'h	31c8;
27287	:douta	=	16'h	5bb3;
27288	:douta	=	16'h	5b93;
27289	:douta	=	16'h	320b;
27290	:douta	=	16'h	0000;
27291	:douta	=	16'h	1106;
27292	:douta	=	16'h	73ad;
27293	:douta	=	16'h	6b2c;
27294	:douta	=	16'h	9cb1;
27295	:douta	=	16'h	630b;
27296	:douta	=	16'h	5269;
27297	:douta	=	16'h	c5f4;
27298	:douta	=	16'h	944f;
27299	:douta	=	16'h	2126;
27300	:douta	=	16'h	7bce;
27301	:douta	=	16'h	840e;
27302	:douta	=	16'h	31a8;
27303	:douta	=	16'h	5aec;
27304	:douta	=	16'h	6b2d;
27305	:douta	=	16'h	5aec;
27306	:douta	=	16'h	a4d1;
27307	:douta	=	16'h	83ef;
27308	:douta	=	16'h	630c;
27309	:douta	=	16'h	840f;
27310	:douta	=	16'h	7b8d;
27311	:douta	=	16'h	5acb;
27312	:douta	=	16'h	3187;
27313	:douta	=	16'h	5249;
27314	:douta	=	16'h	39e7;
27315	:douta	=	16'h	31a6;
27316	:douta	=	16'h	5289;
27317	:douta	=	16'h	5aea;
27318	:douta	=	16'h	3186;
27319	:douta	=	16'h	20e4;
27320	:douta	=	16'h	1041;
27321	:douta	=	16'h	4a08;
27322	:douta	=	16'h	41e7;
27323	:douta	=	16'h	83ef;
27324	:douta	=	16'h	d54f;
27325	:douta	=	16'h	bc8d;
27326	:douta	=	16'h	ac0a;
27327	:douta	=	16'h	ac2a;
27328	:douta	=	16'h	a3ca;
27329	:douta	=	16'h	52ce;
27330	:douta	=	16'h	2a4e;
27331	:douta	=	16'h	21a9;
27332	:douta	=	16'h	3a4c;
27333	:douta	=	16'h	42ae;
27334	:douta	=	16'h	4aad;
27335	:douta	=	16'h	4b0f;
27336	:douta	=	16'h	3a6d;
27337	:douta	=	16'h	1969;
27338	:douta	=	16'h	530f;
27339	:douta	=	16'h	326e;
27340	:douta	=	16'h	328f;
27341	:douta	=	16'h	5b92;
27342	:douta	=	16'h	63d3;
27343	:douta	=	16'h	21ec;
27344	:douta	=	16'h	63b2;
27345	:douta	=	16'h	4b10;
27346	:douta	=	16'h	4310;
27347	:douta	=	16'h	6391;
27348	:douta	=	16'h	72eb;
27349	:douta	=	16'h	6288;
27350	:douta	=	16'h	6289;
27351	:douta	=	16'h	5a48;
27352	:douta	=	16'h	6268;
27353	:douta	=	16'h	4a8e;
27354	:douta	=	16'h	11cd;
27355	:douta	=	16'h	21ec;
27356	:douta	=	16'h	3333;
27357	:douta	=	16'h	3b74;
27358	:douta	=	16'h	5c7a;
27359	:douta	=	16'h	1a2e;
27360	:douta	=	16'h	3b54;
27361	:douta	=	16'h	53f6;
27362	:douta	=	16'h	6478;
27363	:douta	=	16'h	53f6;
27364	:douta	=	16'h	5c37;
27365	:douta	=	16'h	53d6;
27366	:douta	=	16'h	753b;
27367	:douta	=	16'h	6498;
27368	:douta	=	16'h	4b95;
27369	:douta	=	16'h	6479;
27370	:douta	=	16'h	62aa;
27371	:douta	=	16'h	7aca;
27372	:douta	=	16'h	52aa;
27373	:douta	=	16'h	ded7;
27374	:douta	=	16'h	83cc;
27375	:douta	=	16'h	4985;
27376	:douta	=	16'h	28c2;
27377	:douta	=	16'h	3123;
27378	:douta	=	16'h	4164;
27379	:douta	=	16'h	4164;
27380	:douta	=	16'h	4185;
27381	:douta	=	16'h	4185;
27382	:douta	=	16'h	41a6;
27383	:douta	=	16'h	49e7;
27384	:douta	=	16'h	4a08;
27385	:douta	=	16'h	49e8;
27386	:douta	=	16'h	3966;
27387	:douta	=	16'h	39a6;
27388	:douta	=	16'h	41c7;
27389	:douta	=	16'h	49e8;
27390	:douta	=	16'h	41c7;
27391	:douta	=	16'h	39a6;
27392	:douta	=	16'h	3944;
27393	:douta	=	16'h	6c34;
27394	:douta	=	16'h	41a7;
27395	:douta	=	16'h	3945;
27396	:douta	=	16'h	3145;
27397	:douta	=	16'h	2104;
27398	:douta	=	16'h	320a;
27399	:douta	=	16'h	4acf;
27400	:douta	=	16'h	21a9;
27401	:douta	=	16'h	3b33;
27402	:douta	=	16'h	3b12;
27403	:douta	=	16'h	3ad1;
27404	:douta	=	16'h	53b4;
27405	:douta	=	16'h	6c56;
27406	:douta	=	16'h	5373;
27407	:douta	=	16'h	5373;
27408	:douta	=	16'h	63f4;
27409	:douta	=	16'h	4b32;
27410	:douta	=	16'h	8518;
27411	:douta	=	16'h	4aef;
27412	:douta	=	16'h	5b30;
27413	:douta	=	16'h	adb9;
27414	:douta	=	16'h	6bd2;
27415	:douta	=	16'h	8411;
27416	:douta	=	16'h	add9;
27417	:douta	=	16'h	94f6;
27418	:douta	=	16'h	ce19;
27419	:douta	=	16'h	b5b7;
27420	:douta	=	16'h	de78;
27421	:douta	=	16'h	e654;
27422	:douta	=	16'h	e675;
27423	:douta	=	16'h	ee96;
27424	:douta	=	16'h	eeb7;
27425	:douta	=	16'h	e696;
27426	:douta	=	16'h	e696;
27427	:douta	=	16'h	e675;
27428	:douta	=	16'h	e634;
27429	:douta	=	16'h	d5b3;
27430	:douta	=	16'h	cd72;
27431	:douta	=	16'h	c531;
27432	:douta	=	16'h	acd1;
27433	:douta	=	16'h	9451;
27434	:douta	=	16'h	8c11;
27435	:douta	=	16'h	7b70;
27436	:douta	=	16'h	736e;
27437	:douta	=	16'h	732e;
27438	:douta	=	16'h	526a;
27439	:douta	=	16'h	2904;
27440	:douta	=	16'h	a3eb;
27441	:douta	=	16'h	ac2c;
27442	:douta	=	16'h	bc8d;
27443	:douta	=	16'h	d570;
27444	:douta	=	16'h	ddd2;
27445	:douta	=	16'h	e634;
27446	:douta	=	16'h	e675;
27447	:douta	=	16'h	e655;
27448	:douta	=	16'h	d591;
27449	:douta	=	16'h	eeb6;
27450	:douta	=	16'h	ee96;
27451	:douta	=	16'h	ee75;
27452	:douta	=	16'h	ee74;
27453	:douta	=	16'h	83ae;
27454	:douta	=	16'h	83ef;
27455	:douta	=	16'h	a491;
27456	:douta	=	16'h	b4b1;
27457	:douta	=	16'h	a471;
27458	:douta	=	16'h	9431;
27459	:douta	=	16'h	9432;
27460	:douta	=	16'h	83f1;
27461	:douta	=	16'h	83d1;
27462	:douta	=	16'h	83d1;
27463	:douta	=	16'h	7bd1;
27464	:douta	=	16'h	83f1;
27465	:douta	=	16'h	83f1;
27466	:douta	=	16'h	736e;
27467	:douta	=	16'h	736f;
27468	:douta	=	16'h	630e;
27469	:douta	=	16'h	41a7;
27470	:douta	=	16'h	6a46;
27471	:douta	=	16'h	a40a;
27472	:douta	=	16'h	ac0c;
27473	:douta	=	16'h	ccee;
27474	:douta	=	16'h	d590;
27475	:douta	=	16'h	ee75;
27476	:douta	=	16'h	f6d7;
27477	:douta	=	16'h	f6d7;
27478	:douta	=	16'h	f6b6;
27479	:douta	=	16'h	f6b6;
27480	:douta	=	16'h	ee95;
27481	:douta	=	16'h	e633;
27482	:douta	=	16'h	e674;
27483	:douta	=	16'h	ddd2;
27484	:douta	=	16'h	d590;
27485	:douta	=	16'h	bcf0;
27486	:douta	=	16'h	b4d0;
27487	:douta	=	16'h	b4d1;
27488	:douta	=	16'h	9c72;
27489	:douta	=	16'h	9c72;
27490	:douta	=	16'h	acb2;
27491	:douta	=	16'h	9c72;
27492	:douta	=	16'h	9432;
27493	:douta	=	16'h	9453;
27494	:douta	=	16'h	8c32;
27495	:douta	=	16'h	83f1;
27496	:douta	=	16'h	7bd1;
27497	:douta	=	16'h	7bb0;
27498	:douta	=	16'h	83d1;
27499	:douta	=	16'h	7bb0;
27500	:douta	=	16'h	6b2d;
27501	:douta	=	16'h	734d;
27502	:douta	=	16'h	732d;
27503	:douta	=	16'h	62cd;
27504	:douta	=	16'h	49e8;
27505	:douta	=	16'h	8b29;
27506	:douta	=	16'h	bc4b;
27507	:douta	=	16'h	ddb0;
27508	:douta	=	16'h	ddf3;
27509	:douta	=	16'h	ee75;
27510	:douta	=	16'h	d5b2;
27511	:douta	=	16'h	ddb2;
27512	:douta	=	16'h	9c92;
27513	:douta	=	16'h	73f3;
27514	:douta	=	16'h	6bf3;
27515	:douta	=	16'h	6bd2;
27516	:douta	=	16'h	6bd2;
27517	:douta	=	16'h	5330;
27518	:douta	=	16'h	42af;
27519	:douta	=	16'h	3a8e;
27520	:douta	=	16'h	3aae;
27521	:douta	=	16'h	328d;
27522	:douta	=	16'h	21ec;
27523	:douta	=	16'h	2168;
27524	:douta	=	16'h	10a4;
27525	:douta	=	16'h	31ca;
27526	:douta	=	16'h	3a8e;
27527	:douta	=	16'h	2168;
27528	:douta	=	16'h	10c3;
27529	:douta	=	16'h	10e5;
27530	:douta	=	16'h	18e5;
27531	:douta	=	16'h	18e6;
27532	:douta	=	16'h	10e5;
27533	:douta	=	16'h	1926;
27534	:douta	=	16'h	1906;
27535	:douta	=	16'h	1084;
27536	:douta	=	16'h	1083;
27537	:douta	=	16'h	1926;
27538	:douta	=	16'h	1926;
27539	:douta	=	16'h	1926;
27540	:douta	=	16'h	2147;
27541	:douta	=	16'h	1927;
27542	:douta	=	16'h	0000;
27543	:douta	=	16'h	0000;
27544	:douta	=	16'h	0000;
27545	:douta	=	16'h	2146;
27546	:douta	=	16'h	10c4;
27547	:douta	=	16'h	2126;
27548	:douta	=	16'h	1926;
27549	:douta	=	16'h	1906;
27550	:douta	=	16'h	0063;
27551	:douta	=	16'h	7bef;
27552	:douta	=	16'h	8c2f;
27553	:douta	=	16'h	10a4;
27554	:douta	=	16'h	31c8;
27555	:douta	=	16'h	de77;
27556	:douta	=	16'h	ad12;
27557	:douta	=	16'h	4a48;
27558	:douta	=	16'h	840f;
27559	:douta	=	16'h	2986;
27560	:douta	=	16'h	630b;
27561	:douta	=	16'h	736d;
27562	:douta	=	16'h	6b2c;
27563	:douta	=	16'h	a4d2;
27564	:douta	=	16'h	4208;
27565	:douta	=	16'h	52aa;
27566	:douta	=	16'h	6b6d;
27567	:douta	=	16'h	52cb;
27568	:douta	=	16'h	8c4f;
27569	:douta	=	16'h	39e9;
27570	:douta	=	16'h	31a7;
27571	:douta	=	16'h	5acb;
27572	:douta	=	16'h	632c;
27573	:douta	=	16'h	4229;
27574	:douta	=	16'h	39a6;
27575	:douta	=	16'h	39c7;
27576	:douta	=	16'h	62cb;
27577	:douta	=	16'h	acae;
27578	:douta	=	16'h	c56f;
27579	:douta	=	16'h	9348;
27580	:douta	=	16'h	a3ea;
27581	:douta	=	16'h	b44a;
27582	:douta	=	16'h	6aca;
27583	:douta	=	16'h	31c9;
27584	:douta	=	16'h	2a2d;
27585	:douta	=	16'h	428d;
27586	:douta	=	16'h	322b;
27587	:douta	=	16'h	42ae;
27588	:douta	=	16'h	3a6d;
27589	:douta	=	16'h	52ee;
27590	:douta	=	16'h	42ad;
27591	:douta	=	16'h	42ae;
27592	:douta	=	16'h	3a6c;
27593	:douta	=	16'h	530f;
27594	:douta	=	16'h	3aae;
27595	:douta	=	16'h	6370;
27596	:douta	=	16'h	73f2;
27597	:douta	=	16'h	6392;
27598	:douta	=	16'h	326d;
27599	:douta	=	16'h	5b91;
27600	:douta	=	16'h	42f0;
27601	:douta	=	16'h	42d0;
27602	:douta	=	16'h	5351;
27603	:douta	=	16'h	5b71;
27604	:douta	=	16'h	2a6f;
27605	:douta	=	16'h	6371;
27606	:douta	=	16'h	5aaa;
27607	:douta	=	16'h	5a48;
27608	:douta	=	16'h	5a88;
27609	:douta	=	16'h	5a08;
27610	:douta	=	16'h	6289;
27611	:douta	=	16'h	4a8d;
27612	:douta	=	16'h	19ac;
27613	:douta	=	16'h	19ee;
27614	:douta	=	16'h	2b13;
27615	:douta	=	16'h	3334;
27616	:douta	=	16'h	3b75;
27617	:douta	=	16'h	222e;
27618	:douta	=	16'h	3b12;
27619	:douta	=	16'h	4bd5;
27620	:douta	=	16'h	6cfa;
27621	:douta	=	16'h	5c16;
27622	:douta	=	16'h	4373;
27623	:douta	=	16'h	3af1;
27624	:douta	=	16'h	4bf8;
27625	:douta	=	16'h	7cb7;
27626	:douta	=	16'h	7c51;
27627	:douta	=	16'h	b573;
27628	:douta	=	16'h	836c;
27629	:douta	=	16'h	1820;
27630	:douta	=	16'h	4164;
27631	:douta	=	16'h	4985;
27632	:douta	=	16'h	4985;
27633	:douta	=	16'h	49a5;
27634	:douta	=	16'h	49a6;
27635	:douta	=	16'h	41a6;
27636	:douta	=	16'h	49c6;
27637	:douta	=	16'h	4186;
27638	:douta	=	16'h	4166;
27639	:douta	=	16'h	49e7;
27640	:douta	=	16'h	39a6;
27641	:douta	=	16'h	49c7;
27642	:douta	=	16'h	41a7;
27643	:douta	=	16'h	41c7;
27644	:douta	=	16'h	41a7;
27645	:douta	=	16'h	49c7;
27646	:douta	=	16'h	41a7;
27647	:douta	=	16'h	41a7;
27648	:douta	=	16'h	4185;
27649	:douta	=	16'h	6c13;
27650	:douta	=	16'h	526b;
27651	:douta	=	16'h	3945;
27652	:douta	=	16'h	3124;
27653	:douta	=	16'h	2104;
27654	:douta	=	16'h	320a;
27655	:douta	=	16'h	5b51;
27656	:douta	=	16'h	322b;
27657	:douta	=	16'h	4394;
27658	:douta	=	16'h	4353;
27659	:douta	=	16'h	2a0e;
27660	:douta	=	16'h	53d4;
27661	:douta	=	16'h	2a2d;
27662	:douta	=	16'h	6c77;
27663	:douta	=	16'h	5bf5;
27664	:douta	=	16'h	8539;
27665	:douta	=	16'h	7cd8;
27666	:douta	=	16'h	7c55;
27667	:douta	=	16'h	9d59;
27668	:douta	=	16'h	8cd6;
27669	:douta	=	16'h	9517;
27670	:douta	=	16'h	8495;
27671	:douta	=	16'h	630d;
27672	:douta	=	16'h	adfa;
27673	:douta	=	16'h	6bf2;
27674	:douta	=	16'h	b597;
27675	:douta	=	16'h	c65a;
27676	:douta	=	16'h	83f0;
27677	:douta	=	16'h	d5f5;
27678	:douta	=	16'h	ee75;
27679	:douta	=	16'h	e676;
27680	:douta	=	16'h	ee96;
27681	:douta	=	16'h	ee96;
27682	:douta	=	16'h	e675;
27683	:douta	=	16'h	e675;
27684	:douta	=	16'h	de15;
27685	:douta	=	16'h	cd93;
27686	:douta	=	16'h	c552;
27687	:douta	=	16'h	acb1;
27688	:douta	=	16'h	a471;
27689	:douta	=	16'h	8c11;
27690	:douta	=	16'h	83d0;
27691	:douta	=	16'h	7b90;
27692	:douta	=	16'h	7b6f;
27693	:douta	=	16'h	734f;
27694	:douta	=	16'h	2903;
27695	:douta	=	16'h	6a87;
27696	:douta	=	16'h	a46b;
27697	:douta	=	16'h	bccd;
27698	:douta	=	16'h	c52f;
27699	:douta	=	16'h	ddf2;
27700	:douta	=	16'h	e634;
27701	:douta	=	16'h	e675;
27702	:douta	=	16'h	e675;
27703	:douta	=	16'h	ee95;
27704	:douta	=	16'h	cd2f;
27705	:douta	=	16'h	e613;
27706	:douta	=	16'h	ee75;
27707	:douta	=	16'h	e675;
27708	:douta	=	16'h	e654;
27709	:douta	=	16'h	acb0;
27710	:douta	=	16'h	7bae;
27711	:douta	=	16'h	7390;
27712	:douta	=	16'h	9c72;
27713	:douta	=	16'h	a492;
27714	:douta	=	16'h	9431;
27715	:douta	=	16'h	8c31;
27716	:douta	=	16'h	8bf1;
27717	:douta	=	16'h	7bf1;
27718	:douta	=	16'h	7bf1;
27719	:douta	=	16'h	7bd0;
27720	:douta	=	16'h	7bd1;
27721	:douta	=	16'h	7bd1;
27722	:douta	=	16'h	7bb0;
27723	:douta	=	16'h	73b0;
27724	:douta	=	16'h	20c3;
27725	:douta	=	16'h	4984;
27726	:douta	=	16'h	9bab;
27727	:douta	=	16'h	bc8c;
27728	:douta	=	16'h	cd0e;
27729	:douta	=	16'h	ddf1;
27730	:douta	=	16'h	e633;
27731	:douta	=	16'h	ee96;
27732	:douta	=	16'h	eeb7;
27733	:douta	=	16'h	f6d7;
27734	:douta	=	16'h	ee96;
27735	:douta	=	16'h	ee75;
27736	:douta	=	16'h	ee95;
27737	:douta	=	16'h	e634;
27738	:douta	=	16'h	ddd2;
27739	:douta	=	16'h	d591;
27740	:douta	=	16'h	c531;
27741	:douta	=	16'h	acb1;
27742	:douta	=	16'h	9c72;
27743	:douta	=	16'h	a492;
27744	:douta	=	16'h	9c93;
27745	:douta	=	16'h	9472;
27746	:douta	=	16'h	9c93;
27747	:douta	=	16'h	a4b4;
27748	:douta	=	16'h	8c32;
27749	:douta	=	16'h	83f1;
27750	:douta	=	16'h	8412;
27751	:douta	=	16'h	7bd1;
27752	:douta	=	16'h	7bb0;
27753	:douta	=	16'h	7baf;
27754	:douta	=	16'h	7b6f;
27755	:douta	=	16'h	7b8f;
27756	:douta	=	16'h	736e;
27757	:douta	=	16'h	6b2d;
27758	:douta	=	16'h	6aec;
27759	:douta	=	16'h	832b;
27760	:douta	=	16'h	82e9;
27761	:douta	=	16'h	bc4b;
27762	:douta	=	16'h	dd90;
27763	:douta	=	16'h	ee74;
27764	:douta	=	16'h	e634;
27765	:douta	=	16'h	e634;
27766	:douta	=	16'h	d5d3;
27767	:douta	=	16'h	c532;
27768	:douta	=	16'h	9472;
27769	:douta	=	16'h	8434;
27770	:douta	=	16'h	7413;
27771	:douta	=	16'h	73f3;
27772	:douta	=	16'h	6bd2;
27773	:douta	=	16'h	63b2;
27774	:douta	=	16'h	5330;
27775	:douta	=	16'h	5351;
27776	:douta	=	16'h	42d0;
27777	:douta	=	16'h	3acf;
27778	:douta	=	16'h	324d;
27779	:douta	=	16'h	29eb;
27780	:douta	=	16'h	21a9;
27781	:douta	=	16'h	10a5;
27782	:douta	=	16'h	10c4;
27783	:douta	=	16'h	4af0;
27784	:douta	=	16'h	1906;
27785	:douta	=	16'h	0882;
27786	:douta	=	16'h	1105;
27787	:douta	=	16'h	10e5;
27788	:douta	=	16'h	1926;
27789	:douta	=	16'h	2127;
27790	:douta	=	16'h	10e5;
27791	:douta	=	16'h	10a4;
27792	:douta	=	16'h	10e6;
27793	:douta	=	16'h	1927;
27794	:douta	=	16'h	2168;
27795	:douta	=	16'h	1948;
27796	:douta	=	16'h	2168;
27797	:douta	=	16'h	2189;
27798	:douta	=	16'h	1926;
27799	:douta	=	16'h	0883;
27800	:douta	=	16'h	0000;
27801	:douta	=	16'h	0000;
27802	:douta	=	16'h	0883;
27803	:douta	=	16'h	1106;
27804	:douta	=	16'h	1926;
27805	:douta	=	16'h	1927;
27806	:douta	=	16'h	08a3;
27807	:douta	=	16'h	424d;
27808	:douta	=	16'h	8474;
27809	:douta	=	16'h	8431;
27810	:douta	=	16'h	3a09;
27811	:douta	=	16'h	4a49;
27812	:douta	=	16'h	7b8d;
27813	:douta	=	16'h	4a49;
27814	:douta	=	16'h	acf2;
27815	:douta	=	16'h	738e;
27816	:douta	=	16'h	31c7;
27817	:douta	=	16'h	632c;
27818	:douta	=	16'h	6b4c;
27819	:douta	=	16'h	8c2e;
27820	:douta	=	16'h	9cb1;
27821	:douta	=	16'h	5aeb;
27822	:douta	=	16'h	52ab;
27823	:douta	=	16'h	5aab;
27824	:douta	=	16'h	6b6c;
27825	:douta	=	16'h	73cf;
27826	:douta	=	16'h	4a8a;
27827	:douta	=	16'h	4229;
27828	:douta	=	16'h	31a6;
27829	:douta	=	16'h	2124;
27830	:douta	=	16'h	41e7;
27831	:douta	=	16'h	734b;
27832	:douta	=	16'h	bd30;
27833	:douta	=	16'h	b46c;
27834	:douta	=	16'h	9368;
27835	:douta	=	16'h	a3eb;
27836	:douta	=	16'h	a40b;
27837	:douta	=	16'h	72ea;
27838	:douta	=	16'h	1969;
27839	:douta	=	16'h	322c;
27840	:douta	=	16'h	530f;
27841	:douta	=	16'h	2189;
27842	:douta	=	16'h	4aee;
27843	:douta	=	16'h	530f;
27844	:douta	=	16'h	2a0b;
27845	:douta	=	16'h	42ad;
27846	:douta	=	16'h	4ace;
27847	:douta	=	16'h	19aa;
27848	:douta	=	16'h	5b50;
27849	:douta	=	16'h	530f;
27850	:douta	=	16'h	2a2b;
27851	:douta	=	16'h	530f;
27852	:douta	=	16'h	6b91;
27853	:douta	=	16'h	428e;
27854	:douta	=	16'h	3a8e;
27855	:douta	=	16'h	5b71;
27856	:douta	=	16'h	3aaf;
27857	:douta	=	16'h	5bb2;
27858	:douta	=	16'h	42d0;
27859	:douta	=	16'h	6c14;
27860	:douta	=	16'h	2a2c;
27861	:douta	=	16'h	6c14;
27862	:douta	=	16'h	5b92;
27863	:douta	=	16'h	6269;
27864	:douta	=	16'h	6227;
27865	:douta	=	16'h	5a48;
27866	:douta	=	16'h	5228;
27867	:douta	=	16'h	5a69;
27868	:douta	=	16'h	42af;
27869	:douta	=	16'h	196a;
27870	:douta	=	16'h	3334;
27871	:douta	=	16'h	4c18;
27872	:douta	=	16'h	3b54;
27873	:douta	=	16'h	4374;
27874	:douta	=	16'h	4bf7;
27875	:douta	=	16'h	4bf6;
27876	:douta	=	16'h	5c37;
27877	:douta	=	16'h	3af2;
27878	:douta	=	16'h	4332;
27879	:douta	=	16'h	4333;
27880	:douta	=	16'h	5418;
27881	:douta	=	16'h	b5b5;
27882	:douta	=	16'h	944f;
27883	:douta	=	16'h	51e6;
27884	:douta	=	16'h	2060;
27885	:douta	=	16'h	4985;
27886	:douta	=	16'h	49a5;
27887	:douta	=	16'h	49c6;
27888	:douta	=	16'h	49a6;
27889	:douta	=	16'h	49c6;
27890	:douta	=	16'h	49c6;
27891	:douta	=	16'h	49c7;
27892	:douta	=	16'h	49c8;
27893	:douta	=	16'h	4186;
27894	:douta	=	16'h	49c7;
27895	:douta	=	16'h	49e7;
27896	:douta	=	16'h	41c7;
27897	:douta	=	16'h	41a6;
27898	:douta	=	16'h	41a7;
27899	:douta	=	16'h	41a6;
27900	:douta	=	16'h	49e7;
27901	:douta	=	16'h	49e8;
27902	:douta	=	16'h	49c7;
27903	:douta	=	16'h	3146;
27904	:douta	=	16'h	49c6;
27905	:douta	=	16'h	5b0d;
27906	:douta	=	16'h	6391;
27907	:douta	=	16'h	3144;
27908	:douta	=	16'h	2924;
27909	:douta	=	16'h	2903;
27910	:douta	=	16'h	29a9;
27911	:douta	=	16'h	6bf3;
27912	:douta	=	16'h	2189;
27913	:douta	=	16'h	4bd6;
27914	:douta	=	16'h	326f;
27915	:douta	=	16'h	4332;
27916	:douta	=	16'h	6415;
27917	:douta	=	16'h	6416;
27918	:douta	=	16'h	6415;
27919	:douta	=	16'h	5bb4;
27920	:douta	=	16'h	7477;
27921	:douta	=	16'h	5b73;
27922	:douta	=	16'h	6bf3;
27923	:douta	=	16'h	63b2;
27924	:douta	=	16'h	6392;
27925	:douta	=	16'h	9d37;
27926	:douta	=	16'h	94d6;
27927	:douta	=	16'h	8c94;
27928	:douta	=	16'h	b5b8;
27929	:douta	=	16'h	b5d8;
27930	:douta	=	16'h	b5b7;
27931	:douta	=	16'h	b5d8;
27932	:douta	=	16'h	a4d4;
27933	:douta	=	16'h	c639;
27934	:douta	=	16'h	c5f8;
27935	:douta	=	16'h	e654;
27936	:douta	=	16'h	ee96;
27937	:douta	=	16'h	e675;
27938	:douta	=	16'h	e656;
27939	:douta	=	16'h	de34;
27940	:douta	=	16'h	cdd4;
27941	:douta	=	16'h	cdb3;
27942	:douta	=	16'h	b513;
27943	:douta	=	16'h	9471;
27944	:douta	=	16'h	8c31;
27945	:douta	=	16'h	8bf2;
27946	:douta	=	16'h	83b0;
27947	:douta	=	16'h	6b2d;
27948	:douta	=	16'h	4209;
27949	:douta	=	16'h	28e3;
27950	:douta	=	16'h	ac2c;
27951	:douta	=	16'h	ac8d;
27952	:douta	=	16'h	c52f;
27953	:douta	=	16'h	cd90;
27954	:douta	=	16'h	d5d2;
27955	:douta	=	16'h	ee75;
27956	:douta	=	16'h	ee95;
27957	:douta	=	16'h	ee95;
27958	:douta	=	16'h	ee76;
27959	:douta	=	16'h	ee96;
27960	:douta	=	16'h	e634;
27961	:douta	=	16'h	ddd2;
27962	:douta	=	16'h	d5d1;
27963	:douta	=	16'h	e655;
27964	:douta	=	16'h	e653;
27965	:douta	=	16'h	cd71;
27966	:douta	=	16'h	bd11;
27967	:douta	=	16'h	8c12;
27968	:douta	=	16'h	6370;
27969	:douta	=	16'h	5b2f;
27970	:douta	=	16'h	634f;
27971	:douta	=	16'h	7bb1;
27972	:douta	=	16'h	83d1;
27973	:douta	=	16'h	83d1;
27974	:douta	=	16'h	73b0;
27975	:douta	=	16'h	6b6f;
27976	:douta	=	16'h	632e;
27977	:douta	=	16'h	6b4f;
27978	:douta	=	16'h	1905;
27979	:douta	=	16'h	30e1;
27980	:douta	=	16'h	934a;
27981	:douta	=	16'h	abeb;
27982	:douta	=	16'h	bcab;
27983	:douta	=	16'h	de12;
27984	:douta	=	16'h	e675;
27985	:douta	=	16'h	f6d7;
27986	:douta	=	16'h	f6d7;
27987	:douta	=	16'h	eeb7;
27988	:douta	=	16'h	ee96;
27989	:douta	=	16'h	ee96;
27990	:douta	=	16'h	ee95;
27991	:douta	=	16'h	ee75;
27992	:douta	=	16'h	e654;
27993	:douta	=	16'h	e634;
27994	:douta	=	16'h	c511;
27995	:douta	=	16'h	d591;
27996	:douta	=	16'h	c532;
27997	:douta	=	16'h	9c92;
27998	:douta	=	16'h	a4b2;
27999	:douta	=	16'h	9473;
28000	:douta	=	16'h	8413;
28001	:douta	=	16'h	8432;
28002	:douta	=	16'h	8c12;
28003	:douta	=	16'h	8412;
28004	:douta	=	16'h	8c32;
28005	:douta	=	16'h	8bf1;
28006	:douta	=	16'h	83d1;
28007	:douta	=	16'h	83d0;
28008	:douta	=	16'h	7b90;
28009	:douta	=	16'h	7b6e;
28010	:douta	=	16'h	732d;
28011	:douta	=	16'h	62cb;
28012	:douta	=	16'h	6aab;
28013	:douta	=	16'h	832b;
28014	:douta	=	16'h	8b29;
28015	:douta	=	16'h	bc6b;
28016	:douta	=	16'h	e612;
28017	:douta	=	16'h	e674;
28018	:douta	=	16'h	ee95;
28019	:douta	=	16'h	ee75;
28020	:douta	=	16'h	e654;
28021	:douta	=	16'h	de13;
28022	:douta	=	16'h	c532;
28023	:douta	=	16'h	acb1;
28024	:douta	=	16'h	a4b3;
28025	:douta	=	16'h	8453;
28026	:douta	=	16'h	8454;
28027	:douta	=	16'h	7c54;
28028	:douta	=	16'h	7434;
28029	:douta	=	16'h	6bf3;
28030	:douta	=	16'h	6bd3;
28031	:douta	=	16'h	5b92;
28032	:douta	=	16'h	5372;
28033	:douta	=	16'h	5351;
28034	:douta	=	16'h	4b31;
28035	:douta	=	16'h	3ad0;
28036	:douta	=	16'h	3b10;
28037	:douta	=	16'h	2a4d;
28038	:douta	=	16'h	21ca;
28039	:douta	=	16'h	1105;
28040	:douta	=	16'h	2169;
28041	:douta	=	16'h	5311;
28042	:douta	=	16'h	31eb;
28043	:douta	=	16'h	1927;
28044	:douta	=	16'h	1927;
28045	:douta	=	16'h	21a9;
28046	:douta	=	16'h	21a9;
28047	:douta	=	16'h	2168;
28048	:douta	=	16'h	2189;
28049	:douta	=	16'h	1968;
28050	:douta	=	16'h	2147;
28051	:douta	=	16'h	1927;
28052	:douta	=	16'h	1927;
28053	:douta	=	16'h	1948;
28054	:douta	=	16'h	21a9;
28055	:douta	=	16'h	1926;
28056	:douta	=	16'h	1946;
28057	:douta	=	16'h	1926;
28058	:douta	=	16'h	10c5;
28059	:douta	=	16'h	0863;
28060	:douta	=	16'h	0000;
28061	:douta	=	16'h	0021;
28062	:douta	=	16'h	0863;
28063	:douta	=	16'h	39ca;
28064	:douta	=	16'h	6bd2;
28065	:douta	=	16'h	63d2;
28066	:douta	=	16'h	7cb6;
28067	:douta	=	16'h	0000;
28068	:douta	=	16'h	1906;
28069	:douta	=	16'h	1927;
28070	:douta	=	16'h	1106;
28071	:douta	=	16'h	0084;
28072	:douta	=	16'h	83ee;
28073	:douta	=	16'h	2124;
28074	:douta	=	16'h	39a6;
28075	:douta	=	16'h	738d;
28076	:douta	=	16'h	6b4c;
28077	:douta	=	16'h	1925;
28078	:douta	=	16'h	4228;
28079	:douta	=	16'h	634c;
28080	:douta	=	16'h	8410;
28081	:douta	=	16'h	3a29;
28082	:douta	=	16'h	10a4;
28083	:douta	=	16'h	2146;
28084	:douta	=	16'h	2166;
28085	:douta	=	16'h	39a8;
28086	:douta	=	16'h	bcce;
28087	:douta	=	16'h	9348;
28088	:douta	=	16'h	9baa;
28089	:douta	=	16'h	bc4c;
28090	:douta	=	16'h	b44b;
28091	:douta	=	16'h	31a8;
28092	:douta	=	16'h	1128;
28093	:douta	=	16'h	3a2a;
28094	:douta	=	16'h	31e9;
28095	:douta	=	16'h	426c;
28096	:douta	=	16'h	0907;
28097	:douta	=	16'h	6bd1;
28098	:douta	=	16'h	73d1;
28099	:douta	=	16'h	322b;
28100	:douta	=	16'h	6391;
28101	:douta	=	16'h	29cb;
28102	:douta	=	16'h	19aa;
28103	:douta	=	16'h	4aae;
28104	:douta	=	16'h	532f;
28105	:douta	=	16'h	3a8d;
28106	:douta	=	16'h	73d1;
28107	:douta	=	16'h	5330;
28108	:douta	=	16'h	320b;
28109	:douta	=	16'h	42ae;
28110	:douta	=	16'h	5b0e;
28111	:douta	=	16'h	4af0;
28112	:douta	=	16'h	42ee;
28113	:douta	=	16'h	4b10;
28114	:douta	=	16'h	21ec;
28115	:douta	=	16'h	326d;
28116	:douta	=	16'h	5352;
28117	:douta	=	16'h	3aaf;
28118	:douta	=	16'h	3a8e;
28119	:douta	=	16'h	42d0;
28120	:douta	=	16'h	4310;
28121	:douta	=	16'h	526b;
28122	:douta	=	16'h	5207;
28123	:douta	=	16'h	5229;
28124	:douta	=	16'h	49e8;
28125	:douta	=	16'h	5a28;
28126	:douta	=	16'h	424b;
28127	:douta	=	16'h	19cd;
28128	:douta	=	16'h	096a;
28129	:douta	=	16'h	32f2;
28130	:douta	=	16'h	43d6;
28131	:douta	=	16'h	2a6f;
28132	:douta	=	16'h	32b0;
28133	:douta	=	16'h	2a90;
28134	:douta	=	16'h	53d6;
28135	:douta	=	16'h	7c97;
28136	:douta	=	16'h	6b08;
28137	:douta	=	16'h	2881;
28138	:douta	=	16'h	3923;
28139	:douta	=	16'h	4184;
28140	:douta	=	16'h	4185;
28141	:douta	=	16'h	51e6;
28142	:douta	=	16'h	49a5;
28143	:douta	=	16'h	49a7;
28144	:douta	=	16'h	4a08;
28145	:douta	=	16'h	5208;
28146	:douta	=	16'h	4a08;
28147	:douta	=	16'h	41a6;
28148	:douta	=	16'h	4186;
28149	:douta	=	16'h	49e8;
28150	:douta	=	16'h	49c7;
28151	:douta	=	16'h	41a6;
28152	:douta	=	16'h	41a7;
28153	:douta	=	16'h	41c7;
28154	:douta	=	16'h	3987;
28155	:douta	=	16'h	3966;
28156	:douta	=	16'h	3966;
28157	:douta	=	16'h	3966;
28158	:douta	=	16'h	3966;
28159	:douta	=	16'h	3987;
28160	:douta	=	16'h	41a6;
28161	:douta	=	16'h	528b;
28162	:douta	=	16'h	6391;
28163	:douta	=	16'h	3965;
28164	:douta	=	16'h	3124;
28165	:douta	=	16'h	2904;
28166	:douta	=	16'h	2146;
28167	:douta	=	16'h	63d3;
28168	:douta	=	16'h	19a9;
28169	:douta	=	16'h	328f;
28170	:douta	=	16'h	5394;
28171	:douta	=	16'h	6416;
28172	:douta	=	16'h	4b11;
28173	:douta	=	16'h	5393;
28174	:douta	=	16'h	5393;
28175	:douta	=	16'h	4b11;
28176	:douta	=	16'h	7cb7;
28177	:douta	=	16'h	8cf9;
28178	:douta	=	16'h	6bf4;
28179	:douta	=	16'h	9517;
28180	:douta	=	16'h	9517;
28181	:douta	=	16'h	8495;
28182	:douta	=	16'h	8475;
28183	:douta	=	16'h	9d16;
28184	:douta	=	16'h	ad57;
28185	:douta	=	16'h	bdf8;
28186	:douta	=	16'h	bdf9;
28187	:douta	=	16'h	b5b8;
28188	:douta	=	16'h	a4d4;
28189	:douta	=	16'h	b5b6;
28190	:douta	=	16'h	ad57;
28191	:douta	=	16'h	d5f3;
28192	:douta	=	16'h	e654;
28193	:douta	=	16'h	e675;
28194	:douta	=	16'h	de55;
28195	:douta	=	16'h	d614;
28196	:douta	=	16'h	cd93;
28197	:douta	=	16'h	bd32;
28198	:douta	=	16'h	b4f3;
28199	:douta	=	16'h	9472;
28200	:douta	=	16'h	8c31;
28201	:douta	=	16'h	7bd0;
28202	:douta	=	16'h	7b8f;
28203	:douta	=	16'h	6b4f;
28204	:douta	=	16'h	3124;
28205	:douta	=	16'h	7aa7;
28206	:douta	=	16'h	9c4d;
28207	:douta	=	16'h	b48e;
28208	:douta	=	16'h	d5b1;
28209	:douta	=	16'h	d5d1;
28210	:douta	=	16'h	de13;
28211	:douta	=	16'h	e633;
28212	:douta	=	16'h	ee75;
28213	:douta	=	16'h	ee95;
28214	:douta	=	16'h	e675;
28215	:douta	=	16'h	e655;
28216	:douta	=	16'h	e614;
28217	:douta	=	16'h	e634;
28218	:douta	=	16'h	cd50;
28219	:douta	=	16'h	e614;
28220	:douta	=	16'h	de14;
28221	:douta	=	16'h	cd72;
28222	:douta	=	16'h	acd0;
28223	:douta	=	16'h	9471;
28224	:douta	=	16'h	8433;
28225	:douta	=	16'h	7bf2;
28226	:douta	=	16'h	5b2f;
28227	:douta	=	16'h	52ee;
28228	:douta	=	16'h	7390;
28229	:douta	=	16'h	73b1;
28230	:douta	=	16'h	7bf1;
28231	:douta	=	16'h	8c11;
28232	:douta	=	16'h	7bd0;
28233	:douta	=	16'h	62ee;
28234	:douta	=	16'h	38e2;
28235	:douta	=	16'h	82c6;
28236	:douta	=	16'h	b44a;
28237	:douta	=	16'h	ccec;
28238	:douta	=	16'h	e5b0;
28239	:douta	=	16'h	ee75;
28240	:douta	=	16'h	ee95;
28241	:douta	=	16'h	f6b6;
28242	:douta	=	16'h	eeb7;
28243	:douta	=	16'h	ee96;
28244	:douta	=	16'h	e655;
28245	:douta	=	16'h	e634;
28246	:douta	=	16'h	e654;
28247	:douta	=	16'h	e654;
28248	:douta	=	16'h	ddf3;
28249	:douta	=	16'h	ddd2;
28250	:douta	=	16'h	c512;
28251	:douta	=	16'h	c532;
28252	:douta	=	16'h	cd52;
28253	:douta	=	16'h	a4b2;
28254	:douta	=	16'h	9c92;
28255	:douta	=	16'h	8c53;
28256	:douta	=	16'h	8412;
28257	:douta	=	16'h	8412;
28258	:douta	=	16'h	83f1;
28259	:douta	=	16'h	8412;
28260	:douta	=	16'h	8c32;
28261	:douta	=	16'h	83d0;
28262	:douta	=	16'h	83b0;
28263	:douta	=	16'h	7baf;
28264	:douta	=	16'h	7b4e;
28265	:douta	=	16'h	7b6e;
28266	:douta	=	16'h	6b0d;
28267	:douta	=	16'h	628b;
28268	:douta	=	16'h	b46b;
28269	:douta	=	16'h	d54d;
28270	:douta	=	16'h	e5f2;
28271	:douta	=	16'h	d5d2;
28272	:douta	=	16'h	ee95;
28273	:douta	=	16'h	ee96;
28274	:douta	=	16'h	ee75;
28275	:douta	=	16'h	e654;
28276	:douta	=	16'h	ddf3;
28277	:douta	=	16'h	d5d3;
28278	:douta	=	16'h	bd11;
28279	:douta	=	16'h	a492;
28280	:douta	=	16'h	9c93;
28281	:douta	=	16'h	8c94;
28282	:douta	=	16'h	8c74;
28283	:douta	=	16'h	7c54;
28284	:douta	=	16'h	7433;
28285	:douta	=	16'h	7413;
28286	:douta	=	16'h	6bf4;
28287	:douta	=	16'h	63d3;
28288	:douta	=	16'h	5b93;
28289	:douta	=	16'h	5b92;
28290	:douta	=	16'h	4b31;
28291	:douta	=	16'h	3ad0;
28292	:douta	=	16'h	42f0;
28293	:douta	=	16'h	42cf;
28294	:douta	=	16'h	3a6e;
28295	:douta	=	16'h	29ea;
28296	:douta	=	16'h	10e7;
28297	:douta	=	16'h	1928;
28298	:douta	=	16'h	4b10;
28299	:douta	=	16'h	4b31;
28300	:douta	=	16'h	1969;
28301	:douta	=	16'h	29aa;
28302	:douta	=	16'h	2189;
28303	:douta	=	16'h	1926;
28304	:douta	=	16'h	1906;
28305	:douta	=	16'h	1906;
28306	:douta	=	16'h	1105;
28307	:douta	=	16'h	1905;
28308	:douta	=	16'h	1106;
28309	:douta	=	16'h	2147;
28310	:douta	=	16'h	29a9;
28311	:douta	=	16'h	1946;
28312	:douta	=	16'h	1926;
28313	:douta	=	16'h	1907;
28314	:douta	=	16'h	1926;
28315	:douta	=	16'h	2127;
28316	:douta	=	16'h	10a4;
28317	:douta	=	16'h	0883;
28318	:douta	=	16'h	0042;
28319	:douta	=	16'h	0000;
28320	:douta	=	16'h	1063;
28321	:douta	=	16'h	42ad;
28322	:douta	=	16'h	7413;
28323	:douta	=	16'h	0021;
28324	:douta	=	16'h	2127;
28325	:douta	=	16'h	1947;
28326	:douta	=	16'h	1927;
28327	:douta	=	16'h	08a5;
28328	:douta	=	16'h	73d1;
28329	:douta	=	16'h	52ed;
28330	:douta	=	16'h	39e8;
28331	:douta	=	16'h	7bae;
28332	:douta	=	16'h	4a68;
28333	:douta	=	16'h	2966;
28334	:douta	=	16'h	6b6c;
28335	:douta	=	16'h	31e8;
28336	:douta	=	16'h	2986;
28337	:douta	=	16'h	2125;
28338	:douta	=	16'h	0042;
28339	:douta	=	16'h	0083;
28340	:douta	=	16'h	72ea;
28341	:douta	=	16'h	938b;
28342	:douta	=	16'h	a3aa;
28343	:douta	=	16'h	abeb;
28344	:douta	=	16'h	b44b;
28345	:douta	=	16'h	72a8;
28346	:douta	=	16'h	5249;
28347	:douta	=	16'h	21aa;
28348	:douta	=	16'h	1106;
28349	:douta	=	16'h	29c8;
28350	:douta	=	16'h	52cc;
28351	:douta	=	16'h	4acd;
28352	:douta	=	16'h	52ee;
28353	:douta	=	16'h	42ad;
28354	:douta	=	16'h	42cf;
28355	:douta	=	16'h	634f;
28356	:douta	=	16'h	4aad;
28357	:douta	=	16'h	42ce;
28358	:douta	=	16'h	4acf;
28359	:douta	=	16'h	322c;
28360	:douta	=	16'h	326c;
28361	:douta	=	16'h	3a4c;
28362	:douta	=	16'h	530f;
28363	:douta	=	16'h	4ace;
28364	:douta	=	16'h	4ace;
28365	:douta	=	16'h	3a6d;
28366	:douta	=	16'h	3a8d;
28367	:douta	=	16'h	31eb;
28368	:douta	=	16'h	63b1;
28369	:douta	=	16'h	63b1;
28370	:douta	=	16'h	3acf;
28371	:douta	=	16'h	3aaf;
28372	:douta	=	16'h	4b31;
28373	:douta	=	16'h	42d0;
28374	:douta	=	16'h	5350;
28375	:douta	=	16'h	4b30;
28376	:douta	=	16'h	430f;
28377	:douta	=	16'h	4b10;
28378	:douta	=	16'h	5a8b;
28379	:douta	=	16'h	51e7;
28380	:douta	=	16'h	4a08;
28381	:douta	=	16'h	51e8;
28382	:douta	=	16'h	5228;
28383	:douta	=	16'h	42cf;
28384	:douta	=	16'h	19ab;
28385	:douta	=	16'h	32d2;
28386	:douta	=	16'h	4c18;
28387	:douta	=	16'h	32f2;
28388	:douta	=	16'h	3b33;
28389	:douta	=	16'h	3313;
28390	:douta	=	16'h	7c32;
28391	:douta	=	16'h	730a;
28392	:douta	=	16'h	30c2;
28393	:douta	=	16'h	4184;
28394	:douta	=	16'h	4985;
28395	:douta	=	16'h	49c6;
28396	:douta	=	16'h	49a5;
28397	:douta	=	16'h	49c6;
28398	:douta	=	16'h	51e8;
28399	:douta	=	16'h	5a29;
28400	:douta	=	16'h	4a08;
28401	:douta	=	16'h	49c7;
28402	:douta	=	16'h	5229;
28403	:douta	=	16'h	41a7;
28404	:douta	=	16'h	41a7;
28405	:douta	=	16'h	41a7;
28406	:douta	=	16'h	41a6;
28407	:douta	=	16'h	41a7;
28408	:douta	=	16'h	49c7;
28409	:douta	=	16'h	49c7;
28410	:douta	=	16'h	41a7;
28411	:douta	=	16'h	41c7;
28412	:douta	=	16'h	3986;
28413	:douta	=	16'h	41a7;
28414	:douta	=	16'h	41a7;
28415	:douta	=	16'h	41a7;
28416	:douta	=	16'h	41a5;
28417	:douta	=	16'h	3944;
28418	:douta	=	16'h	6390;
28419	:douta	=	16'h	3103;
28420	:douta	=	16'h	3145;
28421	:douta	=	16'h	2924;
28422	:douta	=	16'h	2945;
28423	:douta	=	16'h	31a9;
28424	:douta	=	16'h	328e;
28425	:douta	=	16'h	29a9;
28426	:douta	=	16'h	2168;
28427	:douta	=	16'h	3a2c;
28428	:douta	=	16'h	4acf;
28429	:douta	=	16'h	6391;
28430	:douta	=	16'h	8c31;
28431	:douta	=	16'h	9cb4;
28432	:douta	=	16'h	8d39;
28433	:douta	=	16'h	8c95;
28434	:douta	=	16'h	a537;
28435	:douta	=	16'h	adb9;
28436	:douta	=	16'h	94f6;
28437	:douta	=	16'h	9d56;
28438	:douta	=	16'h	94f5;
28439	:douta	=	16'h	94d5;
28440	:douta	=	16'h	c5d7;
28441	:douta	=	16'h	d679;
28442	:douta	=	16'h	c619;
28443	:douta	=	16'h	8431;
28444	:douta	=	16'h	5b0e;
28445	:douta	=	16'h	7c12;
28446	:douta	=	16'h	ad97;
28447	:douta	=	16'h	de79;
28448	:douta	=	16'h	d69a;
28449	:douta	=	16'h	de14;
28450	:douta	=	16'h	de34;
28451	:douta	=	16'h	d5f3;
28452	:douta	=	16'h	c551;
28453	:douta	=	16'h	b512;
28454	:douta	=	16'h	9451;
28455	:douta	=	16'h	8c11;
28456	:douta	=	16'h	7bb0;
28457	:douta	=	16'h	7390;
28458	:douta	=	16'h	632f;
28459	:douta	=	16'h	28e3;
28460	:douta	=	16'h	b48d;
28461	:douta	=	16'h	b4ad;
28462	:douta	=	16'h	c54f;
28463	:douta	=	16'h	d5b0;
28464	:douta	=	16'h	e634;
28465	:douta	=	16'h	e654;
28466	:douta	=	16'h	e675;
28467	:douta	=	16'h	ee75;
28468	:douta	=	16'h	ddd2;
28469	:douta	=	16'h	e634;
28470	:douta	=	16'h	e654;
28471	:douta	=	16'h	e654;
28472	:douta	=	16'h	de13;
28473	:douta	=	16'h	d5f3;
28474	:douta	=	16'h	d5b2;
28475	:douta	=	16'h	c550;
28476	:douta	=	16'h	c531;
28477	:douta	=	16'h	b512;
28478	:douta	=	16'h	bd12;
28479	:douta	=	16'h	9c92;
28480	:douta	=	16'h	8452;
28481	:douta	=	16'h	8432;
28482	:douta	=	16'h	73b1;
28483	:douta	=	16'h	632f;
28484	:douta	=	16'h	632f;
28485	:douta	=	16'h	630e;
28486	:douta	=	16'h	5ace;
28487	:douta	=	16'h	4aae;
28488	:douta	=	16'h	2947;
28489	:douta	=	16'h	82a7;
28490	:douta	=	16'h	a389;
28491	:douta	=	16'h	e590;
28492	:douta	=	16'h	e633;
28493	:douta	=	16'h	ee34;
28494	:douta	=	16'h	eeb7;
28495	:douta	=	16'h	ee96;
28496	:douta	=	16'h	f6d7;
28497	:douta	=	16'h	eeb6;
28498	:douta	=	16'h	e675;
28499	:douta	=	16'h	eeb6;
28500	:douta	=	16'h	e634;
28501	:douta	=	16'h	e634;
28502	:douta	=	16'h	d5d3;
28503	:douta	=	16'h	cdb3;
28504	:douta	=	16'h	bd32;
28505	:douta	=	16'h	bd12;
28506	:douta	=	16'h	acb2;
28507	:douta	=	16'h	9452;
28508	:douta	=	16'h	9473;
28509	:douta	=	16'h	9c73;
28510	:douta	=	16'h	8c33;
28511	:douta	=	16'h	8432;
28512	:douta	=	16'h	7bb0;
28513	:douta	=	16'h	7bb0;
28514	:douta	=	16'h	7b8f;
28515	:douta	=	16'h	736e;
28516	:douta	=	16'h	732d;
28517	:douta	=	16'h	730d;
28518	:douta	=	16'h	72ec;
28519	:douta	=	16'h	732d;
28520	:douta	=	16'h	7b4d;
28521	:douta	=	16'h	6228;
28522	:douta	=	16'h	936a;
28523	:douta	=	16'h	b44b;
28524	:douta	=	16'h	a3e9;
28525	:douta	=	16'h	a3ca;
28526	:douta	=	16'h	b46b;
28527	:douta	=	16'h	cd0e;
28528	:douta	=	16'h	d590;
28529	:douta	=	16'h	d5d2;
28530	:douta	=	16'h	ddd2;
28531	:douta	=	16'h	cd92;
28532	:douta	=	16'h	cd32;
28533	:douta	=	16'h	c532;
28534	:douta	=	16'h	ac91;
28535	:douta	=	16'h	a492;
28536	:douta	=	16'h	9473;
28537	:douta	=	16'h	94b5;
28538	:douta	=	16'h	8cb5;
28539	:douta	=	16'h	7413;
28540	:douta	=	16'h	7413;
28541	:douta	=	16'h	7433;
28542	:douta	=	16'h	6bf3;
28543	:douta	=	16'h	7413;
28544	:douta	=	16'h	6c14;
28545	:douta	=	16'h	6c14;
28546	:douta	=	16'h	63d4;
28547	:douta	=	16'h	5bd4;
28548	:douta	=	16'h	4b52;
28549	:douta	=	16'h	3a8e;
28550	:douta	=	16'h	324d;
28551	:douta	=	16'h	29cb;
28552	:douta	=	16'h	320c;
28553	:douta	=	16'h	320c;
28554	:douta	=	16'h	2189;
28555	:douta	=	16'h	08c5;
28556	:douta	=	16'h	320b;
28557	:douta	=	16'h	29ea;
28558	:douta	=	16'h	21a9;
28559	:douta	=	16'h	1106;
28560	:douta	=	16'h	0884;
28561	:douta	=	16'h	10e5;
28562	:douta	=	16'h	10e5;
28563	:douta	=	16'h	10e5;
28564	:douta	=	16'h	10c5;
28565	:douta	=	16'h	10e5;
28566	:douta	=	16'h	10e5;
28567	:douta	=	16'h	10e5;
28568	:douta	=	16'h	10e5;
28569	:douta	=	16'h	1926;
28570	:douta	=	16'h	2147;
28571	:douta	=	16'h	1927;
28572	:douta	=	16'h	1947;
28573	:douta	=	16'h	1106;
28574	:douta	=	16'h	1926;
28575	:douta	=	16'h	1927;
28576	:douta	=	16'h	1947;
28577	:douta	=	16'h	1084;
28578	:douta	=	16'h	0000;
28579	:douta	=	16'h	0062;
28580	:douta	=	16'h	0062;
28581	:douta	=	16'h	0884;
28582	:douta	=	16'h	1906;
28583	:douta	=	16'h	10e5;
28584	:douta	=	16'h	7c74;
28585	:douta	=	16'h	7c75;
28586	:douta	=	16'h	84b6;
28587	:douta	=	16'h	6c14;
28588	:douta	=	16'h	6393;
28589	:douta	=	16'h	18e5;
28590	:douta	=	16'h	1906;
28591	:douta	=	16'h	1905;
28592	:douta	=	16'h	18e5;
28593	:douta	=	16'h	08a5;
28594	:douta	=	16'h	c50f;
28595	:douta	=	16'h	d50d;
28596	:douta	=	16'h	b42b;
28597	:douta	=	16'h	bc8c;
28598	:douta	=	16'h	b44b;
28599	:douta	=	16'h	4a4a;
28600	:douta	=	16'h	0086;
28601	:douta	=	16'h	8410;
28602	:douta	=	16'h	634d;
28603	:douta	=	16'h	2168;
28604	:douta	=	16'h	3209;
28605	:douta	=	16'h	426b;
28606	:douta	=	16'h	2188;
28607	:douta	=	16'h	4a8c;
28608	:douta	=	16'h	52ac;
28609	:douta	=	16'h	3a4b;
28610	:douta	=	16'h	29ca;
28611	:douta	=	16'h	320b;
28612	:douta	=	16'h	52ee;
28613	:douta	=	16'h	4ace;
28614	:douta	=	16'h	42ae;
28615	:douta	=	16'h	4b10;
28616	:douta	=	16'h	29aa;
28617	:douta	=	16'h	4ace;
28618	:douta	=	16'h	4ace;
28619	:douta	=	16'h	4b0f;
28620	:douta	=	16'h	634f;
28621	:douta	=	16'h	42ae;
28622	:douta	=	16'h	3a4c;
28623	:douta	=	16'h	530f;
28624	:douta	=	16'h	428d;
28625	:douta	=	16'h	3a6d;
28626	:douta	=	16'h	322d;
28627	:douta	=	16'h	5372;
28628	:douta	=	16'h	328e;
28629	:douta	=	16'h	5b71;
28630	:douta	=	16'h	4b51;
28631	:douta	=	16'h	42f0;
28632	:douta	=	16'h	4b0f;
28633	:douta	=	16'h	63d4;
28634	:douta	=	16'h	21a9;
28635	:douta	=	16'h	3a6c;
28636	:douta	=	16'h	41c7;
28637	:douta	=	16'h	5a49;
28638	:douta	=	16'h	4a08;
28639	:douta	=	16'h	49c7;
28640	:douta	=	16'h	5209;
28641	:douta	=	16'h	3187;
28642	:douta	=	16'h	328f;
28643	:douta	=	16'h	32f2;
28644	:douta	=	16'h	3a4b;
28645	:douta	=	16'h	3923;
28646	:douta	=	16'h	3922;
28647	:douta	=	16'h	4185;
28648	:douta	=	16'h	51c5;
28649	:douta	=	16'h	51c6;
28650	:douta	=	16'h	49a6;
28651	:douta	=	16'h	49a6;
28652	:douta	=	16'h	49c6;
28653	:douta	=	16'h	5228;
28654	:douta	=	16'h	3966;
28655	:douta	=	16'h	4186;
28656	:douta	=	16'h	49e7;
28657	:douta	=	16'h	49c7;
28658	:douta	=	16'h	49e8;
28659	:douta	=	16'h	49c7;
28660	:douta	=	16'h	49e8;
28661	:douta	=	16'h	41a7;
28662	:douta	=	16'h	49e7;
28663	:douta	=	16'h	39a6;
28664	:douta	=	16'h	41a7;
28665	:douta	=	16'h	49e8;
28666	:douta	=	16'h	49e7;
28667	:douta	=	16'h	49e8;
28668	:douta	=	16'h	49c7;
28669	:douta	=	16'h	4a08;
28670	:douta	=	16'h	4a08;
28671	:douta	=	16'h	49e7;
28672	:douta	=	16'h	41a5;
28673	:douta	=	16'h	3923;
28674	:douta	=	16'h	632e;
28675	:douta	=	16'h	3103;
28676	:douta	=	16'h	3125;
28677	:douta	=	16'h	2924;
28678	:douta	=	16'h	3146;
28679	:douta	=	16'h	2967;
28680	:douta	=	16'h	430f;
28681	:douta	=	16'h	29aa;
28682	:douta	=	16'h	21a9;
28683	:douta	=	16'h	1946;
28684	:douta	=	16'h	1926;
28685	:douta	=	16'h	2989;
28686	:douta	=	16'h	836d;
28687	:douta	=	16'h	ac71;
28688	:douta	=	16'h	9c30;
28689	:douta	=	16'h	ac4f;
28690	:douta	=	16'h	a46f;
28691	:douta	=	16'h	bcf1;
28692	:douta	=	16'h	a46f;
28693	:douta	=	16'h	d637;
28694	:douta	=	16'h	ad34;
28695	:douta	=	16'h	8c73;
28696	:douta	=	16'h	632e;
28697	:douta	=	16'h	9471;
28698	:douta	=	16'h	a514;
28699	:douta	=	16'h	b535;
28700	:douta	=	16'h	9492;
28701	:douta	=	16'h	94b4;
28702	:douta	=	16'h	a535;
28703	:douta	=	16'h	ef1a;
28704	:douta	=	16'h	e6fb;
28705	:douta	=	16'h	bd97;
28706	:douta	=	16'h	ee74;
28707	:douta	=	16'h	de13;
28708	:douta	=	16'h	c552;
28709	:douta	=	16'h	acf1;
28710	:douta	=	16'h	9410;
28711	:douta	=	16'h	7b90;
28712	:douta	=	16'h	7b90;
28713	:douta	=	16'h	6b2f;
28714	:douta	=	16'h	39e9;
28715	:douta	=	16'h	936a;
28716	:douta	=	16'h	ac8d;
28717	:douta	=	16'h	c50f;
28718	:douta	=	16'h	d591;
28719	:douta	=	16'h	ddd2;
28720	:douta	=	16'h	e634;
28721	:douta	=	16'h	ee96;
28722	:douta	=	16'h	e654;
28723	:douta	=	16'h	ee96;
28724	:douta	=	16'h	e634;
28725	:douta	=	16'h	e613;
28726	:douta	=	16'h	ddd2;
28727	:douta	=	16'h	ddf3;
28728	:douta	=	16'h	de13;
28729	:douta	=	16'h	d5d2;
28730	:douta	=	16'h	c531;
28731	:douta	=	16'h	bcf0;
28732	:douta	=	16'h	b4d1;
28733	:douta	=	16'h	9c91;
28734	:douta	=	16'h	9c91;
28735	:douta	=	16'h	9c93;
28736	:douta	=	16'h	8433;
28737	:douta	=	16'h	8452;
28738	:douta	=	16'h	7c12;
28739	:douta	=	16'h	73b0;
28740	:douta	=	16'h	630d;
28741	:douta	=	16'h	630f;
28742	:douta	=	16'h	6b71;
28743	:douta	=	16'h	3145;
28744	:douta	=	16'h	40e2;
28745	:douta	=	16'h	b40b;
28746	:douta	=	16'h	c4ae;
28747	:douta	=	16'h	ee53;
28748	:douta	=	16'h	eeb6;
28749	:douta	=	16'h	ee95;
28750	:douta	=	16'h	eeb6;
28751	:douta	=	16'h	ee95;
28752	:douta	=	16'h	ee96;
28753	:douta	=	16'h	ee96;
28754	:douta	=	16'h	e655;
28755	:douta	=	16'h	ee75;
28756	:douta	=	16'h	ddf3;
28757	:douta	=	16'h	d5d3;
28758	:douta	=	16'h	d5b3;
28759	:douta	=	16'h	cd73;
28760	:douta	=	16'h	bd32;
28761	:douta	=	16'h	b512;
28762	:douta	=	16'h	a4b2;
28763	:douta	=	16'h	8c52;
28764	:douta	=	16'h	8c32;
28765	:douta	=	16'h	9473;
28766	:douta	=	16'h	8c53;
28767	:douta	=	16'h	8411;
28768	:douta	=	16'h	7b6f;
28769	:douta	=	16'h	7b4e;
28770	:douta	=	16'h	7b6e;
28771	:douta	=	16'h	736d;
28772	:douta	=	16'h	732c;
28773	:douta	=	16'h	730c;
28774	:douta	=	16'h	732d;
28775	:douta	=	16'h	72eb;
28776	:douta	=	16'h	6227;
28777	:douta	=	16'h	72c8;
28778	:douta	=	16'h	9b6a;
28779	:douta	=	16'h	b42a;
28780	:douta	=	16'h	ddd0;
28781	:douta	=	16'h	e5f2;
28782	:douta	=	16'h	d570;
28783	:douta	=	16'h	ddb1;
28784	:douta	=	16'h	ddd1;
28785	:douta	=	16'h	ddf2;
28786	:douta	=	16'h	ddf3;
28787	:douta	=	16'h	d5b2;
28788	:douta	=	16'h	c532;
28789	:douta	=	16'h	b4f1;
28790	:douta	=	16'h	acd2;
28791	:douta	=	16'h	a4b2;
28792	:douta	=	16'h	9473;
28793	:douta	=	16'h	9494;
28794	:douta	=	16'h	94b5;
28795	:douta	=	16'h	8454;
28796	:douta	=	16'h	7c34;
28797	:douta	=	16'h	7413;
28798	:douta	=	16'h	6bf2;
28799	:douta	=	16'h	6bf3;
28800	:douta	=	16'h	6bf3;
28801	:douta	=	16'h	63d3;
28802	:douta	=	16'h	63d3;
28803	:douta	=	16'h	5b93;
28804	:douta	=	16'h	4b31;
28805	:douta	=	16'h	3aaf;
28806	:douta	=	16'h	3a6e;
28807	:douta	=	16'h	2a0c;
28808	:douta	=	16'h	29eb;
28809	:douta	=	16'h	29ca;
28810	:douta	=	16'h	218a;
28811	:douta	=	16'h	29aa;
28812	:douta	=	16'h	1927;
28813	:douta	=	16'h	2167;
28814	:douta	=	16'h	29a9;
28815	:douta	=	16'h	320c;
28816	:douta	=	16'h	322c;
28817	:douta	=	16'h	1927;
28818	:douta	=	16'h	10c4;
28819	:douta	=	16'h	10e5;
28820	:douta	=	16'h	10e5;
28821	:douta	=	16'h	10e5;
28822	:douta	=	16'h	18e5;
28823	:douta	=	16'h	10c5;
28824	:douta	=	16'h	10e5;
28825	:douta	=	16'h	1927;
28826	:douta	=	16'h	1967;
28827	:douta	=	16'h	2147;
28828	:douta	=	16'h	2147;
28829	:douta	=	16'h	1906;
28830	:douta	=	16'h	1927;
28831	:douta	=	16'h	1927;
28832	:douta	=	16'h	1946;
28833	:douta	=	16'h	2147;
28834	:douta	=	16'h	1926;
28835	:douta	=	16'h	10e5;
28836	:douta	=	16'h	0883;
28837	:douta	=	16'h	0021;
28838	:douta	=	16'h	0042;
28839	:douta	=	16'h	0041;
28840	:douta	=	16'h	10a4;
28841	:douta	=	16'h	2146;
28842	:douta	=	16'h	4acc;
28843	:douta	=	16'h	6370;
28844	:douta	=	16'h	7c14;
28845	:douta	=	16'h	0884;
28846	:douta	=	16'h	2147;
28847	:douta	=	16'h	1906;
28848	:douta	=	16'h	18e5;
28849	:douta	=	16'h	29c9;
28850	:douta	=	16'h	73b0;
28851	:douta	=	16'h	734d;
28852	:douta	=	16'h	834b;
28853	:douta	=	16'h	49e5;
28854	:douta	=	16'h	5228;
28855	:douta	=	16'h	29eb;
28856	:douta	=	16'h	422c;
28857	:douta	=	16'h	4aab;
28858	:douta	=	16'h	634e;
28859	:douta	=	16'h	422b;
28860	:douta	=	16'h	52ed;
28861	:douta	=	16'h	73b0;
28862	:douta	=	16'h	08a6;
28863	:douta	=	16'h	1968;
28864	:douta	=	16'h	52ee;
28865	:douta	=	16'h	4a8b;
28866	:douta	=	16'h	6b8f;
28867	:douta	=	16'h	426c;
28868	:douta	=	16'h	320c;
28869	:douta	=	16'h	324c;
28870	:douta	=	16'h	5b2f;
28871	:douta	=	16'h	4aae;
28872	:douta	=	16'h	530f;
28873	:douta	=	16'h	5b70;
28874	:douta	=	16'h	42af;
28875	:douta	=	16'h	320b;
28876	:douta	=	16'h	320b;
28877	:douta	=	16'h	322b;
28878	:douta	=	16'h	6b90;
28879	:douta	=	16'h	63b1;
28880	:douta	=	16'h	21aa;
28881	:douta	=	16'h	3a2d;
28882	:douta	=	16'h	530f;
28883	:douta	=	16'h	42ef;
28884	:douta	=	16'h	5b92;
28885	:douta	=	16'h	4311;
28886	:douta	=	16'h	3aaf;
28887	:douta	=	16'h	5352;
28888	:douta	=	16'h	29ea;
28889	:douta	=	16'h	31ca;
28890	:douta	=	16'h	21aa;
28891	:douta	=	16'h	31ea;
28892	:douta	=	16'h	840f;
28893	:douta	=	16'h	6aab;
28894	:douta	=	16'h	5229;
28895	:douta	=	16'h	49c7;
28896	:douta	=	16'h	49c6;
28897	:douta	=	16'h	3ab0;
28898	:douta	=	16'h	4396;
28899	:douta	=	16'h	3166;
28900	:douta	=	16'h	38e1;
28901	:douta	=	16'h	4164;
28902	:douta	=	16'h	49c6;
28903	:douta	=	16'h	51e7;
28904	:douta	=	16'h	49c6;
28905	:douta	=	16'h	49a6;
28906	:douta	=	16'h	51e7;
28907	:douta	=	16'h	51e7;
28908	:douta	=	16'h	49c7;
28909	:douta	=	16'h	49e8;
28910	:douta	=	16'h	41c7;
28911	:douta	=	16'h	4186;
28912	:douta	=	16'h	49e8;
28913	:douta	=	16'h	49c7;
28914	:douta	=	16'h	41a7;
28915	:douta	=	16'h	49e8;
28916	:douta	=	16'h	49e7;
28917	:douta	=	16'h	41a7;
28918	:douta	=	16'h	49e7;
28919	:douta	=	16'h	41a7;
28920	:douta	=	16'h	41c7;
28921	:douta	=	16'h	49c7;
28922	:douta	=	16'h	49c7;
28923	:douta	=	16'h	41a7;
28924	:douta	=	16'h	41a7;
28925	:douta	=	16'h	41c7;
28926	:douta	=	16'h	41c7;
28927	:douta	=	16'h	49e7;
28928	:douta	=	16'h	41a5;
28929	:douta	=	16'h	3944;
28930	:douta	=	16'h	4a09;
28931	:douta	=	16'h	3965;
28932	:douta	=	16'h	3945;
28933	:douta	=	16'h	3125;
28934	:douta	=	16'h	3125;
28935	:douta	=	16'h	20e5;
28936	:douta	=	16'h	4b50;
28937	:douta	=	16'h	29ca;
28938	:douta	=	16'h	322b;
28939	:douta	=	16'h	2189;
28940	:douta	=	16'h	2168;
28941	:douta	=	16'h	29a9;
28942	:douta	=	16'h	6aea;
28943	:douta	=	16'h	b490;
28944	:douta	=	16'h	ac2e;
28945	:douta	=	16'h	ac2e;
28946	:douta	=	16'h	a42e;
28947	:douta	=	16'h	9bed;
28948	:douta	=	16'h	a42d;
28949	:douta	=	16'h	c4af;
28950	:douta	=	16'h	9c2e;
28951	:douta	=	16'h	630d;
28952	:douta	=	16'h	634e;
28953	:douta	=	16'h	7bd0;
28954	:douta	=	16'h	6bd0;
28955	:douta	=	16'h	6baf;
28956	:douta	=	16'h	638f;
28957	:douta	=	16'h	6b8f;
28958	:douta	=	16'h	73f0;
28959	:douta	=	16'h	634e;
28960	:douta	=	16'h	7bf0;
28961	:douta	=	16'h	8c52;
28962	:douta	=	16'h	7c31;
28963	:douta	=	16'h	9450;
28964	:douta	=	16'h	ddd3;
28965	:douta	=	16'h	acb1;
28966	:douta	=	16'h	8bcf;
28967	:douta	=	16'h	736f;
28968	:douta	=	16'h	62ef;
28969	:douta	=	16'h	7288;
28970	:douta	=	16'h	ac4b;
28971	:douta	=	16'h	c52f;
28972	:douta	=	16'h	cd6f;
28973	:douta	=	16'h	ddd2;
28974	:douta	=	16'h	e654;
28975	:douta	=	16'h	ee75;
28976	:douta	=	16'h	e675;
28977	:douta	=	16'h	ee75;
28978	:douta	=	16'h	e675;
28979	:douta	=	16'h	e654;
28980	:douta	=	16'h	ee75;
28981	:douta	=	16'h	ddd2;
28982	:douta	=	16'h	d5b2;
28983	:douta	=	16'h	d591;
28984	:douta	=	16'h	cd72;
28985	:douta	=	16'h	cd92;
28986	:douta	=	16'h	c572;
28987	:douta	=	16'h	a4b2;
28988	:douta	=	16'h	a4b2;
28989	:douta	=	16'h	9472;
28990	:douta	=	16'h	8c32;
28991	:douta	=	16'h	7bf1;
28992	:douta	=	16'h	7bd1;
28993	:douta	=	16'h	7bd1;
28994	:douta	=	16'h	734f;
28995	:douta	=	16'h	6b2e;
28996	:douta	=	16'h	6b4f;
28997	:douta	=	16'h	31a7;
28998	:douta	=	16'h	30e2;
28999	:douta	=	16'h	9b88;
29000	:douta	=	16'h	a3ea;
29001	:douta	=	16'h	d56e;
29002	:douta	=	16'h	f6b5;
29003	:douta	=	16'h	cdb2;
29004	:douta	=	16'h	c4cf;
29005	:douta	=	16'h	f6b6;
29006	:douta	=	16'h	ee76;
29007	:douta	=	16'h	ee75;
29008	:douta	=	16'h	ee75;
29009	:douta	=	16'h	e654;
29010	:douta	=	16'h	de14;
29011	:douta	=	16'h	cd72;
29012	:douta	=	16'h	d5d3;
29013	:douta	=	16'h	cd73;
29014	:douta	=	16'h	b512;
29015	:douta	=	16'h	b4f3;
29016	:douta	=	16'h	a4d3;
29017	:douta	=	16'h	a493;
29018	:douta	=	16'h	9c93;
29019	:douta	=	16'h	9452;
29020	:douta	=	16'h	8c52;
29021	:douta	=	16'h	7bd0;
29022	:douta	=	16'h	83d0;
29023	:douta	=	16'h	8c11;
29024	:douta	=	16'h	7b6e;
29025	:douta	=	16'h	736d;
29026	:douta	=	16'h	732c;
29027	:douta	=	16'h	732d;
29028	:douta	=	16'h	834e;
29029	:douta	=	16'h	72ea;
29030	:douta	=	16'h	6a69;
29031	:douta	=	16'h	932a;
29032	:douta	=	16'h	abea;
29033	:douta	=	16'h	d54e;
29034	:douta	=	16'h	e653;
29035	:douta	=	16'h	eeb6;
29036	:douta	=	16'h	ee75;
29037	:douta	=	16'h	ee75;
29038	:douta	=	16'h	ee75;
29039	:douta	=	16'h	e674;
29040	:douta	=	16'h	e654;
29041	:douta	=	16'h	ddd3;
29042	:douta	=	16'h	cd71;
29043	:douta	=	16'h	bd12;
29044	:douta	=	16'h	acb2;
29045	:douta	=	16'h	a492;
29046	:douta	=	16'h	9452;
29047	:douta	=	16'h	9432;
29048	:douta	=	16'h	7bf1;
29049	:douta	=	16'h	8433;
29050	:douta	=	16'h	8433;
29051	:douta	=	16'h	8474;
29052	:douta	=	16'h	8454;
29053	:douta	=	16'h	73f2;
29054	:douta	=	16'h	6b91;
29055	:douta	=	16'h	6371;
29056	:douta	=	16'h	5b51;
29057	:douta	=	16'h	5331;
29058	:douta	=	16'h	5331;
29059	:douta	=	16'h	5351;
29060	:douta	=	16'h	5351;
29061	:douta	=	16'h	428f;
29062	:douta	=	16'h	322d;
29063	:douta	=	16'h	324d;
29064	:douta	=	16'h	4af0;
29065	:douta	=	16'h	42f1;
29066	:douta	=	16'h	322c;
29067	:douta	=	16'h	21ca;
29068	:douta	=	16'h	5310;
29069	:douta	=	16'h	3a2c;
29070	:douta	=	16'h	29ea;
29071	:douta	=	16'h	2168;
29072	:douta	=	16'h	10e6;
29073	:douta	=	16'h	1084;
29074	:douta	=	16'h	29aa;
29075	:douta	=	16'h	320c;
29076	:douta	=	16'h	21ca;
29077	:douta	=	16'h	1906;
29078	:douta	=	16'h	2147;
29079	:douta	=	16'h	1926;
29080	:douta	=	16'h	1927;
29081	:douta	=	16'h	2168;
29082	:douta	=	16'h	1927;
29083	:douta	=	16'h	1927;
29084	:douta	=	16'h	1926;
29085	:douta	=	16'h	1927;
29086	:douta	=	16'h	1926;
29087	:douta	=	16'h	1927;
29088	:douta	=	16'h	1927;
29089	:douta	=	16'h	1926;
29090	:douta	=	16'h	1106;
29091	:douta	=	16'h	1906;
29092	:douta	=	16'h	1105;
29093	:douta	=	16'h	1926;
29094	:douta	=	16'h	2127;
29095	:douta	=	16'h	2127;
29096	:douta	=	16'h	2126;
29097	:douta	=	16'h	1905;
29098	:douta	=	16'h	18e5;
29099	:douta	=	16'h	0021;
29100	:douta	=	16'h	0000;
29101	:douta	=	16'h	0021;
29102	:douta	=	16'h	0001;
29103	:douta	=	16'h	0021;
29104	:douta	=	16'h	0842;
29105	:douta	=	16'h	10c4;
29106	:douta	=	16'h	6391;
29107	:douta	=	16'h	6bf4;
29108	:douta	=	16'h	8d1a;
29109	:douta	=	16'h	4b10;
29110	:douta	=	16'h	10e5;
29111	:douta	=	16'h	1106;
29112	:douta	=	16'h	08a4;
29113	:douta	=	16'h	3a2a;
29114	:douta	=	16'h	426b;
29115	:douta	=	16'h	52ad;
29116	:douta	=	16'h	636f;
29117	:douta	=	16'h	52ac;
29118	:douta	=	16'h	636e;
29119	:douta	=	16'h	5b0e;
29120	:douta	=	16'h	424a;
29121	:douta	=	16'h	6b8f;
29122	:douta	=	16'h	52cc;
29123	:douta	=	16'h	3a2c;
29124	:douta	=	16'h	52ee;
29125	:douta	=	16'h	42ae;
29126	:douta	=	16'h	3a6c;
29127	:douta	=	16'h	5b50;
29128	:douta	=	16'h	8453;
29129	:douta	=	16'h	42ce;
29130	:douta	=	16'h	3a2b;
29131	:douta	=	16'h	42ad;
29132	:douta	=	16'h	29eb;
29133	:douta	=	16'h	6bd1;
29134	:douta	=	16'h	63b1;
29135	:douta	=	16'h	21ca;
29136	:douta	=	16'h	4acf;
29137	:douta	=	16'h	5350;
29138	:douta	=	16'h	320b;
29139	:douta	=	16'h	5b2f;
29140	:douta	=	16'h	5350;
29141	:douta	=	16'h	42ad;
29142	:douta	=	16'h	29aa;
29143	:douta	=	16'h	320a;
29144	:douta	=	16'h	3a6d;
29145	:douta	=	16'h	4a4b;
29146	:douta	=	16'h	93ed;
29147	:douta	=	16'h	6ac9;
29148	:douta	=	16'h	49a7;
29149	:douta	=	16'h	5207;
29150	:douta	=	16'h	524b;
29151	:douta	=	16'h	2a8f;
29152	:douta	=	16'h	32d1;
29153	:douta	=	16'h	4985;
29154	:douta	=	16'h	5142;
29155	:douta	=	16'h	51a5;
29156	:douta	=	16'h	5a06;
29157	:douta	=	16'h	5a07;
29158	:douta	=	16'h	4185;
29159	:douta	=	16'h	49c6;
29160	:douta	=	16'h	49e7;
29161	:douta	=	16'h	41a6;
29162	:douta	=	16'h	4166;
29163	:douta	=	16'h	4186;
29164	:douta	=	16'h	41a7;
29165	:douta	=	16'h	49e8;
29166	:douta	=	16'h	49e8;
29167	:douta	=	16'h	49e8;
29168	:douta	=	16'h	4a08;
29169	:douta	=	16'h	49e8;
29170	:douta	=	16'h	49e8;
29171	:douta	=	16'h	49e7;
29172	:douta	=	16'h	49e7;
29173	:douta	=	16'h	41a7;
29174	:douta	=	16'h	41a7;
29175	:douta	=	16'h	41c7;
29176	:douta	=	16'h	41a6;
29177	:douta	=	16'h	41a7;
29178	:douta	=	16'h	41c7;
29179	:douta	=	16'h	41c7;
29180	:douta	=	16'h	49c7;
29181	:douta	=	16'h	49c7;
29182	:douta	=	16'h	41a7;
29183	:douta	=	16'h	49e7;
29184	:douta	=	16'h	4185;
29185	:douta	=	16'h	3964;
29186	:douta	=	16'h	3966;
29187	:douta	=	16'h	4228;
29188	:douta	=	16'h	3145;
29189	:douta	=	16'h	3124;
29190	:douta	=	16'h	3145;
29191	:douta	=	16'h	20e4;
29192	:douta	=	16'h	4b50;
29193	:douta	=	16'h	29a9;
29194	:douta	=	16'h	29a9;
29195	:douta	=	16'h	29a9;
29196	:douta	=	16'h	2167;
29197	:douta	=	16'h	31ca;
29198	:douta	=	16'h	5a6a;
29199	:douta	=	16'h	ac2e;
29200	:douta	=	16'h	a40e;
29201	:douta	=	16'h	ac4e;
29202	:douta	=	16'h	a40e;
29203	:douta	=	16'h	a3ee;
29204	:douta	=	16'h	ac4e;
29205	:douta	=	16'h	bcce;
29206	:douta	=	16'h	940e;
29207	:douta	=	16'h	630d;
29208	:douta	=	16'h	6b6f;
29209	:douta	=	16'h	73d0;
29210	:douta	=	16'h	73d0;
29211	:douta	=	16'h	73f0;
29212	:douta	=	16'h	73d1;
29213	:douta	=	16'h	638f;
29214	:douta	=	16'h	73d1;
29215	:douta	=	16'h	6bb1;
29216	:douta	=	16'h	6370;
29217	:douta	=	16'h	6bf1;
29218	:douta	=	16'h	6390;
29219	:douta	=	16'h	3aab;
29220	:douta	=	16'h	bcf1;
29221	:douta	=	16'h	cd73;
29222	:douta	=	16'h	736e;
29223	:douta	=	16'h	62ad;
29224	:douta	=	16'h	41a8;
29225	:douta	=	16'h	c4cd;
29226	:douta	=	16'h	c50d;
29227	:douta	=	16'h	d590;
29228	:douta	=	16'h	d5d2;
29229	:douta	=	16'h	e634;
29230	:douta	=	16'h	e694;
29231	:douta	=	16'h	ee96;
29232	:douta	=	16'h	ee75;
29233	:douta	=	16'h	e613;
29234	:douta	=	16'h	ee75;
29235	:douta	=	16'h	e654;
29236	:douta	=	16'h	e654;
29237	:douta	=	16'h	ddf3;
29238	:douta	=	16'h	d591;
29239	:douta	=	16'h	cd91;
29240	:douta	=	16'h	c531;
29241	:douta	=	16'h	bd31;
29242	:douta	=	16'h	cd93;
29243	:douta	=	16'h	a4d3;
29244	:douta	=	16'h	9c93;
29245	:douta	=	16'h	9453;
29246	:douta	=	16'h	8c32;
29247	:douta	=	16'h	7bd1;
29248	:douta	=	16'h	734e;
29249	:douta	=	16'h	734e;
29250	:douta	=	16'h	732e;
29251	:douta	=	16'h	6b4e;
29252	:douta	=	16'h	5acc;
29253	:douta	=	16'h	4143;
29254	:douta	=	16'h	82c6;
29255	:douta	=	16'h	ac0b;
29256	:douta	=	16'h	c4ac;
29257	:douta	=	16'h	ddd0;
29258	:douta	=	16'h	ff18;
29259	:douta	=	16'h	e674;
29260	:douta	=	16'h	7b2d;
29261	:douta	=	16'h	d52f;
29262	:douta	=	16'h	eeb6;
29263	:douta	=	16'h	e653;
29264	:douta	=	16'h	e654;
29265	:douta	=	16'h	de13;
29266	:douta	=	16'h	ddf3;
29267	:douta	=	16'h	c552;
29268	:douta	=	16'h	c533;
29269	:douta	=	16'h	bd13;
29270	:douta	=	16'h	a4d3;
29271	:douta	=	16'h	acd3;
29272	:douta	=	16'h	a4b3;
29273	:douta	=	16'h	9c72;
29274	:douta	=	16'h	9452;
29275	:douta	=	16'h	8c32;
29276	:douta	=	16'h	8c11;
29277	:douta	=	16'h	7bb0;
29278	:douta	=	16'h	736e;
29279	:douta	=	16'h	7b8f;
29280	:douta	=	16'h	7b8f;
29281	:douta	=	16'h	7b8e;
29282	:douta	=	16'h	7b6e;
29283	:douta	=	16'h	7b8e;
29284	:douta	=	16'h	6268;
29285	:douta	=	16'h	938a;
29286	:douta	=	16'h	bc6d;
29287	:douta	=	16'h	c50e;
29288	:douta	=	16'h	ddb0;
29289	:douta	=	16'h	ee95;
29290	:douta	=	16'h	ee96;
29291	:douta	=	16'h	e695;
29292	:douta	=	16'h	ee96;
29293	:douta	=	16'h	eeb5;
29294	:douta	=	16'h	e655;
29295	:douta	=	16'h	de13;
29296	:douta	=	16'h	d5f2;
29297	:douta	=	16'h	cd52;
29298	:douta	=	16'h	bcb1;
29299	:douta	=	16'h	a472;
29300	:douta	=	16'h	9c72;
29301	:douta	=	16'h	9c92;
29302	:douta	=	16'h	9431;
29303	:douta	=	16'h	7bf1;
29304	:douta	=	16'h	7bd1;
29305	:douta	=	16'h	7c12;
29306	:douta	=	16'h	7bf2;
29307	:douta	=	16'h	7c12;
29308	:douta	=	16'h	7c13;
29309	:douta	=	16'h	73d2;
29310	:douta	=	16'h	6bb2;
29311	:douta	=	16'h	73d2;
29312	:douta	=	16'h	5b50;
29313	:douta	=	16'h	5b51;
29314	:douta	=	16'h	6392;
29315	:douta	=	16'h	63f4;
29316	:douta	=	16'h	6435;
29317	:douta	=	16'h	5372;
29318	:douta	=	16'h	4af0;
29319	:douta	=	16'h	4af0;
29320	:douta	=	16'h	5374;
29321	:douta	=	16'h	3aaf;
29322	:douta	=	16'h	42cf;
29323	:douta	=	16'h	2189;
29324	:douta	=	16'h	5310;
29325	:douta	=	16'h	4b10;
29326	:douta	=	16'h	3a8e;
29327	:douta	=	16'h	324e;
29328	:douta	=	16'h	328e;
29329	:douta	=	16'h	2168;
29330	:douta	=	16'h	0882;
29331	:douta	=	16'h	18e5;
29332	:douta	=	16'h	32ae;
29333	:douta	=	16'h	3a8f;
29334	:douta	=	16'h	10e6;
29335	:douta	=	16'h	1948;
29336	:douta	=	16'h	1947;
29337	:douta	=	16'h	2147;
29338	:douta	=	16'h	1927;
29339	:douta	=	16'h	1906;
29340	:douta	=	16'h	1927;
29341	:douta	=	16'h	1947;
29342	:douta	=	16'h	1927;
29343	:douta	=	16'h	1947;
29344	:douta	=	16'h	1946;
29345	:douta	=	16'h	1906;
29346	:douta	=	16'h	1926;
29347	:douta	=	16'h	10c5;
29348	:douta	=	16'h	10e5;
29349	:douta	=	16'h	1926;
29350	:douta	=	16'h	1926;
29351	:douta	=	16'h	1926;
29352	:douta	=	16'h	1926;
29353	:douta	=	16'h	1927;
29354	:douta	=	16'h	1926;
29355	:douta	=	16'h	2127;
29356	:douta	=	16'h	2147;
29357	:douta	=	16'h	18e5;
29358	:douta	=	16'h	18e5;
29359	:douta	=	16'h	0883;
29360	:douta	=	16'h	0863;
29361	:douta	=	16'h	0001;
29362	:douta	=	16'h	0000;
29363	:douta	=	16'h	10a2;
29364	:douta	=	16'h	426d;
29365	:douta	=	16'h	3a2b;
29366	:douta	=	16'h	10e5;
29367	:douta	=	16'h	1927;
29368	:douta	=	16'h	1906;
29369	:douta	=	16'h	0022;
29370	:douta	=	16'h	52ad;
29371	:douta	=	16'h	634e;
29372	:douta	=	16'h	424b;
29373	:douta	=	16'h	52ed;
29374	:douta	=	16'h	73d0;
29375	:douta	=	16'h	5b2e;
29376	:douta	=	16'h	3a0a;
29377	:douta	=	16'h	3a4b;
29378	:douta	=	16'h	4aad;
29379	:douta	=	16'h	08e5;
29380	:douta	=	16'h	426b;
29381	:douta	=	16'h	3a8d;
29382	:douta	=	16'h	6b90;
29383	:douta	=	16'h	532e;
29384	:douta	=	16'h	5b50;
29385	:douta	=	16'h	322c;
29386	:douta	=	16'h	6390;
29387	:douta	=	16'h	3a4c;
29388	:douta	=	16'h	636f;
29389	:douta	=	16'h	532f;
29390	:douta	=	16'h	5b2f;
29391	:douta	=	16'h	320b;
29392	:douta	=	16'h	5b50;
29393	:douta	=	16'h	4b30;
29394	:douta	=	16'h	4acd;
29395	:douta	=	16'h	29e9;
29396	:douta	=	16'h	31a8;
29397	:douta	=	16'h	428c;
29398	:douta	=	16'h	29aa;
29399	:douta	=	16'h	31e9;
29400	:douta	=	16'h	4a6a;
29401	:douta	=	16'h	62a9;
29402	:douta	=	16'h	49a7;
29403	:douta	=	16'h	5207;
29404	:douta	=	16'h	5208;
29405	:douta	=	16'h	49c7;
29406	:douta	=	16'h	53f5;
29407	:douta	=	16'h	21a9;
29408	:douta	=	16'h	5207;
29409	:douta	=	16'h	59e4;
29410	:douta	=	16'h	5a25;
29411	:douta	=	16'h	6227;
29412	:douta	=	16'h	49a5;
29413	:douta	=	16'h	4165;
29414	:douta	=	16'h	6228;
29415	:douta	=	16'h	5207;
29416	:douta	=	16'h	4186;
29417	:douta	=	16'h	41c7;
29418	:douta	=	16'h	4187;
29419	:douta	=	16'h	41a7;
29420	:douta	=	16'h	3966;
29421	:douta	=	16'h	49e8;
29422	:douta	=	16'h	49c7;
29423	:douta	=	16'h	49c7;
29424	:douta	=	16'h	49c7;
29425	:douta	=	16'h	49e8;
29426	:douta	=	16'h	49e8;
29427	:douta	=	16'h	49c7;
29428	:douta	=	16'h	49e7;
29429	:douta	=	16'h	41c7;
29430	:douta	=	16'h	41c7;
29431	:douta	=	16'h	41c7;
29432	:douta	=	16'h	41c7;
29433	:douta	=	16'h	49e8;
29434	:douta	=	16'h	41a7;
29435	:douta	=	16'h	41c7;
29436	:douta	=	16'h	49e8;
29437	:douta	=	16'h	49e7;
29438	:douta	=	16'h	41c7;
29439	:douta	=	16'h	41c7;
29440	:douta	=	16'h	3924;
29441	:douta	=	16'h	4165;
29442	:douta	=	16'h	30e3;
29443	:douta	=	16'h	5b2e;
29444	:douta	=	16'h	3145;
29445	:douta	=	16'h	3124;
29446	:douta	=	16'h	3125;
29447	:douta	=	16'h	2904;
29448	:douta	=	16'h	4a6b;
29449	:douta	=	16'h	2a2b;
29450	:douta	=	16'h	2168;
29451	:douta	=	16'h	29c9;
29452	:douta	=	16'h	2188;
29453	:douta	=	16'h	2188;
29454	:douta	=	16'h	522a;
29455	:douta	=	16'h	a3ed;
29456	:douta	=	16'h	a42e;
29457	:douta	=	16'h	ac2e;
29458	:douta	=	16'h	a42e;
29459	:douta	=	16'h	9bed;
29460	:douta	=	16'h	ac4e;
29461	:douta	=	16'h	ac6e;
29462	:douta	=	16'h	83ae;
29463	:douta	=	16'h	52cd;
29464	:douta	=	16'h	632e;
29465	:douta	=	16'h	6b6f;
29466	:douta	=	16'h	73cf;
29467	:douta	=	16'h	6baf;
29468	:douta	=	16'h	636e;
29469	:douta	=	16'h	6b8f;
29470	:douta	=	16'h	6baf;
29471	:douta	=	16'h	6bb0;
29472	:douta	=	16'h	6bd0;
29473	:douta	=	16'h	7411;
29474	:douta	=	16'h	6bd0;
29475	:douta	=	16'h	636f;
29476	:douta	=	16'h	63af;
29477	:douta	=	16'h	530d;
29478	:douta	=	16'h	7bef;
29479	:douta	=	16'h	bc8d;
29480	:douta	=	16'h	dd8f;
29481	:douta	=	16'h	cd6f;
29482	:douta	=	16'h	ddd2;
29483	:douta	=	16'h	de53;
29484	:douta	=	16'h	e674;
29485	:douta	=	16'h	e655;
29486	:douta	=	16'h	eeb6;
29487	:douta	=	16'h	eeb6;
29488	:douta	=	16'h	e634;
29489	:douta	=	16'h	e675;
29490	:douta	=	16'h	e654;
29491	:douta	=	16'h	e674;
29492	:douta	=	16'h	e654;
29493	:douta	=	16'h	d5b2;
29494	:douta	=	16'h	c552;
29495	:douta	=	16'h	bd11;
29496	:douta	=	16'h	a493;
29497	:douta	=	16'h	9c72;
29498	:douta	=	16'h	a4d2;
29499	:douta	=	16'h	9c92;
29500	:douta	=	16'h	9472;
29501	:douta	=	16'h	8412;
29502	:douta	=	16'h	7bf1;
29503	:douta	=	16'h	7b70;
29504	:douta	=	16'h	736f;
29505	:douta	=	16'h	734e;
29506	:douta	=	16'h	736f;
29507	:douta	=	16'h	5a6a;
29508	:douta	=	16'h	6245;
29509	:douta	=	16'h	ac2c;
29510	:douta	=	16'h	b44a;
29511	:douta	=	16'h	e5d0;
29512	:douta	=	16'h	ee75;
29513	:douta	=	16'h	f6b6;
29514	:douta	=	16'h	eeb6;
29515	:douta	=	16'h	f6f7;
29516	:douta	=	16'h	93ee;
29517	:douta	=	16'h	62ce;
29518	:douta	=	16'h	c4ef;
29519	:douta	=	16'h	e613;
29520	:douta	=	16'h	ddd2;
29521	:douta	=	16'h	c552;
29522	:douta	=	16'h	b4f2;
29523	:douta	=	16'h	acb2;
29524	:douta	=	16'h	a4b3;
29525	:douta	=	16'h	a4b3;
29526	:douta	=	16'h	9c72;
29527	:douta	=	16'h	9452;
29528	:douta	=	16'h	9452;
29529	:douta	=	16'h	9452;
29530	:douta	=	16'h	8c10;
29531	:douta	=	16'h	83d0;
29532	:douta	=	16'h	7b8e;
29533	:douta	=	16'h	734d;
29534	:douta	=	16'h	732d;
29535	:douta	=	16'h	732d;
29536	:douta	=	16'h	6b0c;
29537	:douta	=	16'h	6b0d;
29538	:douta	=	16'h	4165;
29539	:douta	=	16'h	51a5;
29540	:douta	=	16'h	834a;
29541	:douta	=	16'h	ac0a;
29542	:douta	=	16'h	bc8c;
29543	:douta	=	16'h	d58f;
29544	:douta	=	16'h	de12;
29545	:douta	=	16'h	e613;
29546	:douta	=	16'h	e655;
29547	:douta	=	16'h	e675;
29548	:douta	=	16'h	e613;
29549	:douta	=	16'h	ddd2;
29550	:douta	=	16'h	ddf3;
29551	:douta	=	16'h	ddd2;
29552	:douta	=	16'h	d5b3;
29553	:douta	=	16'h	c531;
29554	:douta	=	16'h	bd12;
29555	:douta	=	16'h	b4d2;
29556	:douta	=	16'h	9c72;
29557	:douta	=	16'h	9452;
29558	:douta	=	16'h	9c72;
29559	:douta	=	16'h	9452;
29560	:douta	=	16'h	8412;
29561	:douta	=	16'h	7bf2;
29562	:douta	=	16'h	7bf2;
29563	:douta	=	16'h	6b4f;
29564	:douta	=	16'h	6b70;
29565	:douta	=	16'h	6b70;
29566	:douta	=	16'h	6b91;
29567	:douta	=	16'h	6b91;
29568	:douta	=	16'h	73d2;
29569	:douta	=	16'h	6bb1;
29570	:douta	=	16'h	6371;
29571	:douta	=	16'h	5b10;
29572	:douta	=	16'h	5b10;
29573	:douta	=	16'h	52ad;
29574	:douta	=	16'h	4ace;
29575	:douta	=	16'h	5aee;
29576	:douta	=	16'h	bcef;
29577	:douta	=	16'h	acf3;
29578	:douta	=	16'h	5331;
29579	:douta	=	16'h	3a4d;
29580	:douta	=	16'h	3a4d;
29581	:douta	=	16'h	6bd3;
29582	:douta	=	16'h	5351;
29583	:douta	=	16'h	3aae;
29584	:douta	=	16'h	42af;
29585	:douta	=	16'h	4b10;
29586	:douta	=	16'h	322d;
29587	:douta	=	16'h	29cb;
29588	:douta	=	16'h	1106;
29589	:douta	=	16'h	0863;
29590	:douta	=	16'h	29ca;
29591	:douta	=	16'h	322d;
29592	:douta	=	16'h	2989;
29593	:douta	=	16'h	1947;
29594	:douta	=	16'h	1926;
29595	:douta	=	16'h	1907;
29596	:douta	=	16'h	1926;
29597	:douta	=	16'h	1947;
29598	:douta	=	16'h	1946;
29599	:douta	=	16'h	1927;
29600	:douta	=	16'h	1906;
29601	:douta	=	16'h	1106;
29602	:douta	=	16'h	1105;
29603	:douta	=	16'h	10e5;
29604	:douta	=	16'h	10e6;
29605	:douta	=	16'h	1906;
29606	:douta	=	16'h	1906;
29607	:douta	=	16'h	1105;
29608	:douta	=	16'h	10e6;
29609	:douta	=	16'h	1926;
29610	:douta	=	16'h	10e5;
29611	:douta	=	16'h	10e5;
29612	:douta	=	16'h	18e5;
29613	:douta	=	16'h	1905;
29614	:douta	=	16'h	1905;
29615	:douta	=	16'h	1926;
29616	:douta	=	16'h	1926;
29617	:douta	=	16'h	2187;
29618	:douta	=	16'h	2168;
29619	:douta	=	16'h	2988;
29620	:douta	=	16'h	2147;
29621	:douta	=	16'h	10c5;
29622	:douta	=	16'h	0862;
29623	:douta	=	16'h	0000;
29624	:douta	=	16'h	0862;
29625	:douta	=	16'h	0863;
29626	:douta	=	16'h	4aad;
29627	:douta	=	16'h	5373;
29628	:douta	=	16'h	4b0f;
29629	:douta	=	16'h	422a;
29630	:douta	=	16'h	5b2f;
29631	:douta	=	16'h	6b90;
29632	:douta	=	16'h	8410;
29633	:douta	=	16'h	426b;
29634	:douta	=	16'h	31ea;
29635	:douta	=	16'h	5b0e;
29636	:douta	=	16'h	6b70;
29637	:douta	=	16'h	632e;
29638	:douta	=	16'h	634f;
29639	:douta	=	16'h	5b70;
29640	:douta	=	16'h	322b;
29641	:douta	=	16'h	5b50;
29642	:douta	=	16'h	3a2b;
29643	:douta	=	16'h	5b50;
29644	:douta	=	16'h	6370;
29645	:douta	=	16'h	428d;
29646	:douta	=	16'h	428d;
29647	:douta	=	16'h	5330;
29648	:douta	=	16'h	322b;
29649	:douta	=	16'h	530e;
29650	:douta	=	16'h	1906;
29651	:douta	=	16'h	29a8;
29652	:douta	=	16'h	4229;
29653	:douta	=	16'h	a48e;
29654	:douta	=	16'h	a48d;
29655	:douta	=	16'h	6268;
29656	:douta	=	16'h	5a48;
29657	:douta	=	16'h	6247;
29658	:douta	=	16'h	52ac;
29659	:douta	=	16'h	4aaf;
29660	:douta	=	16'h	2a4e;
29661	:douta	=	16'h	4b94;
29662	:douta	=	16'h	5248;
29663	:douta	=	16'h	6a66;
29664	:douta	=	16'h	6246;
29665	:douta	=	16'h	6a68;
29666	:douta	=	16'h	51e6;
29667	:douta	=	16'h	51e6;
29668	:douta	=	16'h	5a28;
29669	:douta	=	16'h	5a29;
29670	:douta	=	16'h	41a7;
29671	:douta	=	16'h	49c8;
29672	:douta	=	16'h	49c8;
29673	:douta	=	16'h	41a7;
29674	:douta	=	16'h	49c8;
29675	:douta	=	16'h	49e8;
29676	:douta	=	16'h	41a7;
29677	:douta	=	16'h	49c7;
29678	:douta	=	16'h	49c7;
29679	:douta	=	16'h	41a7;
29680	:douta	=	16'h	41a7;
29681	:douta	=	16'h	41c7;
29682	:douta	=	16'h	49c7;
29683	:douta	=	16'h	49c7;
29684	:douta	=	16'h	49c8;
29685	:douta	=	16'h	49e7;
29686	:douta	=	16'h	49e8;
29687	:douta	=	16'h	49c7;
29688	:douta	=	16'h	49e8;
29689	:douta	=	16'h	49e8;
29690	:douta	=	16'h	49e8;
29691	:douta	=	16'h	49e8;
29692	:douta	=	16'h	41a6;
29693	:douta	=	16'h	41c7;
29694	:douta	=	16'h	41a7;
29695	:douta	=	16'h	41c7;
29696	:douta	=	16'h	3105;
29697	:douta	=	16'h	4185;
29698	:douta	=	16'h	3903;
29699	:douta	=	16'h	5b4f;
29700	:douta	=	16'h	3124;
29701	:douta	=	16'h	3125;
29702	:douta	=	16'h	3125;
29703	:douta	=	16'h	2924;
29704	:douta	=	16'h	4a2a;
29705	:douta	=	16'h	29ca;
29706	:douta	=	16'h	2189;
29707	:douta	=	16'h	29c9;
29708	:douta	=	16'h	2988;
29709	:douta	=	16'h	2188;
29710	:douta	=	16'h	3188;
29711	:douta	=	16'h	936c;
29712	:douta	=	16'h	ac6e;
29713	:douta	=	16'h	ac4e;
29714	:douta	=	16'h	a3ed;
29715	:douta	=	16'h	9bee;
29716	:douta	=	16'h	b46e;
29717	:douta	=	16'h	a44e;
29718	:douta	=	16'h	838e;
29719	:douta	=	16'h	52ac;
29720	:douta	=	16'h	634e;
29721	:douta	=	16'h	6b6f;
29722	:douta	=	16'h	73d0;
29723	:douta	=	16'h	6baf;
29724	:douta	=	16'h	634e;
29725	:douta	=	16'h	636e;
29726	:douta	=	16'h	636e;
29727	:douta	=	16'h	73d0;
29728	:douta	=	16'h	6bd0;
29729	:douta	=	16'h	6bd0;
29730	:douta	=	16'h	6bf0;
29731	:douta	=	16'h	6b8f;
29732	:douta	=	16'h	6bae;
29733	:douta	=	16'h	63af;
29734	:douta	=	16'h	5b8e;
29735	:douta	=	16'h	ee33;
29736	:douta	=	16'h	eeb5;
29737	:douta	=	16'h	d5b1;
29738	:douta	=	16'h	e633;
29739	:douta	=	16'h	e654;
29740	:douta	=	16'h	e674;
29741	:douta	=	16'h	e675;
29742	:douta	=	16'h	ee96;
29743	:douta	=	16'h	eeb6;
29744	:douta	=	16'h	e634;
29745	:douta	=	16'h	ee54;
29746	:douta	=	16'h	e654;
29747	:douta	=	16'h	de13;
29748	:douta	=	16'h	e614;
29749	:douta	=	16'h	d5b2;
29750	:douta	=	16'h	c532;
29751	:douta	=	16'h	b4d2;
29752	:douta	=	16'h	9c92;
29753	:douta	=	16'h	9472;
29754	:douta	=	16'h	9c93;
29755	:douta	=	16'h	8c52;
29756	:douta	=	16'h	8c52;
29757	:douta	=	16'h	8412;
29758	:douta	=	16'h	7bf1;
29759	:douta	=	16'h	738f;
29760	:douta	=	16'h	732e;
29761	:douta	=	16'h	6b4e;
29762	:douta	=	16'h	5249;
29763	:douta	=	16'h	41a5;
29764	:douta	=	16'h	a3ca;
29765	:douta	=	16'h	bc8c;
29766	:douta	=	16'h	cced;
29767	:douta	=	16'h	ee74;
29768	:douta	=	16'h	eeb6;
29769	:douta	=	16'h	eeb7;
29770	:douta	=	16'h	ee96;
29771	:douta	=	16'h	eeb6;
29772	:douta	=	16'h	cd92;
29773	:douta	=	16'h	836e;
29774	:douta	=	16'h	7b4d;
29775	:douta	=	16'h	c531;
29776	:douta	=	16'h	d592;
29777	:douta	=	16'h	bd12;
29778	:douta	=	16'h	b4f2;
29779	:douta	=	16'h	b4d3;
29780	:douta	=	16'h	a493;
29781	:douta	=	16'h	9473;
29782	:douta	=	16'h	8c52;
29783	:douta	=	16'h	8c11;
29784	:douta	=	16'h	83f1;
29785	:douta	=	16'h	8bf1;
29786	:douta	=	16'h	8410;
29787	:douta	=	16'h	7b8f;
29788	:douta	=	16'h	736d;
29789	:douta	=	16'h	732d;
29790	:douta	=	16'h	7b6d;
29791	:douta	=	16'h	732d;
29792	:douta	=	16'h	6b2c;
29793	:douta	=	16'h	49c7;
29794	:douta	=	16'h	6a87;
29795	:douta	=	16'h	8b29;
29796	:douta	=	16'h	bcad;
29797	:douta	=	16'h	ddb0;
29798	:douta	=	16'h	e5f3;
29799	:douta	=	16'h	e613;
29800	:douta	=	16'h	e633;
29801	:douta	=	16'h	e633;
29802	:douta	=	16'h	e612;
29803	:douta	=	16'h	e633;
29804	:douta	=	16'h	e654;
29805	:douta	=	16'h	ddd2;
29806	:douta	=	16'h	cd51;
29807	:douta	=	16'h	c510;
29808	:douta	=	16'h	c531;
29809	:douta	=	16'h	bd11;
29810	:douta	=	16'h	bcd2;
29811	:douta	=	16'h	ac92;
29812	:douta	=	16'h	9452;
29813	:douta	=	16'h	8411;
29814	:douta	=	16'h	83f1;
29815	:douta	=	16'h	8412;
29816	:douta	=	16'h	7bd1;
29817	:douta	=	16'h	7bb1;
29818	:douta	=	16'h	6b4f;
29819	:douta	=	16'h	6b4f;
29820	:douta	=	16'h	6b91;
29821	:douta	=	16'h	73b2;
29822	:douta	=	16'h	6bb2;
29823	:douta	=	16'h	73b1;
29824	:douta	=	16'h	6bd2;
29825	:douta	=	16'h	73b1;
29826	:douta	=	16'h	6391;
29827	:douta	=	16'h	6370;
29828	:douta	=	16'h	5b0f;
29829	:douta	=	16'h	424d;
29830	:douta	=	16'h	4a2d;
29831	:douta	=	16'h	d591;
29832	:douta	=	16'h	a4f4;
29833	:douta	=	16'h	73f3;
29834	:douta	=	16'h	6351;
29835	:douta	=	16'h	42ce;
29836	:douta	=	16'h	322c;
29837	:douta	=	16'h	6bd3;
29838	:douta	=	16'h	5b92;
29839	:douta	=	16'h	3a8e;
29840	:douta	=	16'h	3aae;
29841	:douta	=	16'h	4b10;
29842	:douta	=	16'h	42af;
29843	:douta	=	16'h	42af;
29844	:douta	=	16'h	2a0c;
29845	:douta	=	16'h	21aa;
29846	:douta	=	16'h	0884;
29847	:douta	=	16'h	29aa;
29848	:douta	=	16'h	3a6f;
29849	:douta	=	16'h	1927;
29850	:douta	=	16'h	18e6;
29851	:douta	=	16'h	1947;
29852	:douta	=	16'h	2148;
29853	:douta	=	16'h	1907;
29854	:douta	=	16'h	1906;
29855	:douta	=	16'h	1106;
29856	:douta	=	16'h	1906;
29857	:douta	=	16'h	1926;
29858	:douta	=	16'h	1926;
29859	:douta	=	16'h	10e5;
29860	:douta	=	16'h	1906;
29861	:douta	=	16'h	1906;
29862	:douta	=	16'h	1906;
29863	:douta	=	16'h	1905;
29864	:douta	=	16'h	10e5;
29865	:douta	=	16'h	1105;
29866	:douta	=	16'h	10e5;
29867	:douta	=	16'h	10c5;
29868	:douta	=	16'h	1905;
29869	:douta	=	16'h	1926;
29870	:douta	=	16'h	1905;
29871	:douta	=	16'h	1906;
29872	:douta	=	16'h	1906;
29873	:douta	=	16'h	10e5;
29874	:douta	=	16'h	1906;
29875	:douta	=	16'h	10e6;
29876	:douta	=	16'h	2168;
29877	:douta	=	16'h	2988;
29878	:douta	=	16'h	2168;
29879	:douta	=	16'h	10e4;
29880	:douta	=	16'h	0062;
29881	:douta	=	16'h	0000;
29882	:douta	=	16'h	2987;
29883	:douta	=	16'h	7c97;
29884	:douta	=	16'h	6c76;
29885	:douta	=	16'h	29eb;
29886	:douta	=	16'h	2126;
29887	:douta	=	16'h	4acd;
29888	:douta	=	16'h	7bf1;
29889	:douta	=	16'h	4a8c;
29890	:douta	=	16'h	4aad;
29891	:douta	=	16'h	6b6f;
29892	:douta	=	16'h	4acc;
29893	:douta	=	16'h	6bb0;
29894	:douta	=	16'h	634f;
29895	:douta	=	16'h	3a2c;
29896	:douta	=	16'h	94b3;
29897	:douta	=	16'h	636f;
29898	:douta	=	16'h	29ea;
29899	:douta	=	16'h	21aa;
29900	:douta	=	16'h	6390;
29901	:douta	=	16'h	1128;
29902	:douta	=	16'h	428c;
29903	:douta	=	16'h	5b71;
29904	:douta	=	16'h	2146;
29905	:douta	=	16'h	1965;
29906	:douta	=	16'h	3a4a;
29907	:douta	=	16'h	29c9;
29908	:douta	=	16'h	bd11;
29909	:douta	=	16'h	8b6b;
29910	:douta	=	16'h	59e7;
29911	:douta	=	16'h	6a88;
29912	:douta	=	16'h	6a67;
29913	:douta	=	16'h	4a09;
29914	:douta	=	16'h	4b11;
29915	:douta	=	16'h	4312;
29916	:douta	=	16'h	63f6;
29917	:douta	=	16'h	4b53;
29918	:douta	=	16'h	82c6;
29919	:douta	=	16'h	6247;
29920	:douta	=	16'h	6246;
29921	:douta	=	16'h	6247;
29922	:douta	=	16'h	51e6;
29923	:douta	=	16'h	5a48;
29924	:douta	=	16'h	51e7;
29925	:douta	=	16'h	49c7;
29926	:douta	=	16'h	41a7;
29927	:douta	=	16'h	41a7;
29928	:douta	=	16'h	49e8;
29929	:douta	=	16'h	4a08;
29930	:douta	=	16'h	49c8;
29931	:douta	=	16'h	49e8;
29932	:douta	=	16'h	49e8;
29933	:douta	=	16'h	49c7;
29934	:douta	=	16'h	49c7;
29935	:douta	=	16'h	41c7;
29936	:douta	=	16'h	4186;
29937	:douta	=	16'h	41c7;
29938	:douta	=	16'h	49e8;
29939	:douta	=	16'h	49c7;
29940	:douta	=	16'h	49c7;
29941	:douta	=	16'h	49e8;
29942	:douta	=	16'h	49e8;
29943	:douta	=	16'h	5249;
29944	:douta	=	16'h	49e8;
29945	:douta	=	16'h	49c7;
29946	:douta	=	16'h	49e7;
29947	:douta	=	16'h	41a7;
29948	:douta	=	16'h	41a6;
29949	:douta	=	16'h	41a7;
29950	:douta	=	16'h	41a6;
29951	:douta	=	16'h	41a7;
29952	:douta	=	16'h	3124;
29953	:douta	=	16'h	4165;
29954	:douta	=	16'h	4165;
29955	:douta	=	16'h	5b4f;
29956	:douta	=	16'h	30e3;
29957	:douta	=	16'h	3145;
29958	:douta	=	16'h	3124;
29959	:douta	=	16'h	3145;
29960	:douta	=	16'h	49e8;
29961	:douta	=	16'h	2168;
29962	:douta	=	16'h	2189;
29963	:douta	=	16'h	29a9;
29964	:douta	=	16'h	2188;
29965	:douta	=	16'h	2188;
29966	:douta	=	16'h	2989;
29967	:douta	=	16'h	6aab;
29968	:douta	=	16'h	a42e;
29969	:douta	=	16'h	ac2e;
29970	:douta	=	16'h	9bed;
29971	:douta	=	16'h	a40e;
29972	:douta	=	16'h	ac6e;
29973	:douta	=	16'h	9c0e;
29974	:douta	=	16'h	734d;
29975	:douta	=	16'h	5aee;
29976	:douta	=	16'h	636f;
29977	:douta	=	16'h	6b8f;
29978	:douta	=	16'h	634e;
29979	:douta	=	16'h	6b6e;
29980	:douta	=	16'h	6b6e;
29981	:douta	=	16'h	6bd0;
29982	:douta	=	16'h	73d1;
29983	:douta	=	16'h	6bb0;
29984	:douta	=	16'h	73f0;
29985	:douta	=	16'h	6bb0;
29986	:douta	=	16'h	63cf;
29987	:douta	=	16'h	638f;
29988	:douta	=	16'h	6bcf;
29989	:douta	=	16'h	6baf;
29990	:douta	=	16'h	73f0;
29991	:douta	=	16'h	636e;
29992	:douta	=	16'h	bcf0;
29993	:douta	=	16'h	e654;
29994	:douta	=	16'h	e654;
29995	:douta	=	16'h	e674;
29996	:douta	=	16'h	e655;
29997	:douta	=	16'h	e675;
29998	:douta	=	16'h	ee96;
29999	:douta	=	16'h	e696;
30000	:douta	=	16'h	e654;
30001	:douta	=	16'h	d5d2;
30002	:douta	=	16'h	d5b2;
30003	:douta	=	16'h	d5b2;
30004	:douta	=	16'h	cd92;
30005	:douta	=	16'h	bd11;
30006	:douta	=	16'h	a471;
30007	:douta	=	16'h	9c71;
30008	:douta	=	16'h	9471;
30009	:douta	=	16'h	9452;
30010	:douta	=	16'h	8433;
30011	:douta	=	16'h	7bd0;
30012	:douta	=	16'h	7390;
30013	:douta	=	16'h	736f;
30014	:douta	=	16'h	7b90;
30015	:douta	=	16'h	7b90;
30016	:douta	=	16'h	62ec;
30017	:douta	=	16'h	49e6;
30018	:douta	=	16'h	8b6a;
30019	:douta	=	16'h	b44b;
30020	:douta	=	16'h	bcee;
30021	:douta	=	16'h	ddf2;
30022	:douta	=	16'h	e655;
30023	:douta	=	16'h	eeb7;
30024	:douta	=	16'h	eeb6;
30025	:douta	=	16'h	ee95;
30026	:douta	=	16'h	ee96;
30027	:douta	=	16'h	e674;
30028	:douta	=	16'h	ddd2;
30029	:douta	=	16'h	ddf4;
30030	:douta	=	16'h	ac6f;
30031	:douta	=	16'h	8bce;
30032	:douta	=	16'h	734d;
30033	:douta	=	16'h	7b6e;
30034	:douta	=	16'h	9410;
30035	:douta	=	16'h	a493;
30036	:douta	=	16'h	9cb3;
30037	:douta	=	16'h	9c94;
30038	:douta	=	16'h	9452;
30039	:douta	=	16'h	8c32;
30040	:douta	=	16'h	8c31;
30041	:douta	=	16'h	8c11;
30042	:douta	=	16'h	7bae;
30043	:douta	=	16'h	7b8e;
30044	:douta	=	16'h	7bae;
30045	:douta	=	16'h	7b8f;
30046	:douta	=	16'h	7b6f;
30047	:douta	=	16'h	49c7;
30048	:douta	=	16'h	7ac7;
30049	:douta	=	16'h	bc6d;
30050	:douta	=	16'h	bc4b;
30051	:douta	=	16'h	dd90;
30052	:douta	=	16'h	ddf3;
30053	:douta	=	16'h	ee95;
30054	:douta	=	16'h	ee75;
30055	:douta	=	16'h	ee96;
30056	:douta	=	16'h	ee96;
30057	:douta	=	16'h	eeb6;
30058	:douta	=	16'h	ee95;
30059	:douta	=	16'h	e654;
30060	:douta	=	16'h	ee95;
30061	:douta	=	16'h	ee74;
30062	:douta	=	16'h	e612;
30063	:douta	=	16'h	ddb2;
30064	:douta	=	16'h	d592;
30065	:douta	=	16'h	bd11;
30066	:douta	=	16'h	acb1;
30067	:douta	=	16'h	9c93;
30068	:douta	=	16'h	8412;
30069	:douta	=	16'h	83f1;
30070	:douta	=	16'h	83f1;
30071	:douta	=	16'h	7bb0;
30072	:douta	=	16'h	7b6f;
30073	:douta	=	16'h	736f;
30074	:douta	=	16'h	6b4f;
30075	:douta	=	16'h	630d;
30076	:douta	=	16'h	62cd;
30077	:douta	=	16'h	62cd;
30078	:douta	=	16'h	6b2e;
30079	:douta	=	16'h	736f;
30080	:douta	=	16'h	6b2e;
30081	:douta	=	16'h	6b70;
30082	:douta	=	16'h	5b0e;
30083	:douta	=	16'h	62cd;
30084	:douta	=	16'h	9bad;
30085	:douta	=	16'h	ee53;
30086	:douta	=	16'h	e633;
30087	:douta	=	16'h	b4f1;
30088	:douta	=	16'h	b4d2;
30089	:douta	=	16'h	acd2;
30090	:douta	=	16'h	73f2;
30091	:douta	=	16'h	6392;
30092	:douta	=	16'h	2a0c;
30093	:douta	=	16'h	6392;
30094	:douta	=	16'h	6bf3;
30095	:douta	=	16'h	5b72;
30096	:douta	=	16'h	4af0;
30097	:douta	=	16'h	42d0;
30098	:douta	=	16'h	4acf;
30099	:douta	=	16'h	42ae;
30100	:douta	=	16'h	42af;
30101	:douta	=	16'h	4b10;
30102	:douta	=	16'h	3a4d;
30103	:douta	=	16'h	2189;
30104	:douta	=	16'h	1128;
30105	:douta	=	16'h	322d;
30106	:douta	=	16'h	42af;
30107	:douta	=	16'h	320c;
30108	:douta	=	16'h	2168;
30109	:douta	=	16'h	1967;
30110	:douta	=	16'h	10e4;
30111	:douta	=	16'h	10c5;
30112	:douta	=	16'h	10e6;
30113	:douta	=	16'h	10e6;
30114	:douta	=	16'h	1926;
30115	:douta	=	16'h	10e6;
30116	:douta	=	16'h	18e5;
30117	:douta	=	16'h	1926;
30118	:douta	=	16'h	10c5;
30119	:douta	=	16'h	1105;
30120	:douta	=	16'h	10e5;
30121	:douta	=	16'h	18e5;
30122	:douta	=	16'h	10e5;
30123	:douta	=	16'h	10e5;
30124	:douta	=	16'h	1906;
30125	:douta	=	16'h	1905;
30126	:douta	=	16'h	2146;
30127	:douta	=	16'h	18e5;
30128	:douta	=	16'h	10c4;
30129	:douta	=	16'h	10e5;
30130	:douta	=	16'h	18e5;
30131	:douta	=	16'h	1905;
30132	:douta	=	16'h	18e5;
30133	:douta	=	16'h	10e4;
30134	:douta	=	16'h	10e4;
30135	:douta	=	16'h	1905;
30136	:douta	=	16'h	1906;
30137	:douta	=	16'h	2167;
30138	:douta	=	16'h	2188;
30139	:douta	=	16'h	0000;
30140	:douta	=	16'h	2126;
30141	:douta	=	16'h	3a0a;
30142	:douta	=	16'h	1926;
30143	:douta	=	16'h	1947;
30144	:douta	=	16'h	10e5;
30145	:douta	=	16'h	3a2b;
30146	:douta	=	16'h	5b4f;
30147	:douta	=	16'h	6b90;
30148	:douta	=	16'h	5b2e;
30149	:douta	=	16'h	632e;
30150	:douta	=	16'h	9cd3;
30151	:douta	=	16'h	8c31;
30152	:douta	=	16'h	4acd;
30153	:douta	=	16'h	4ace;
30154	:douta	=	16'h	6bb0;
30155	:douta	=	16'h	5b30;
30156	:douta	=	16'h	21ca;
30157	:douta	=	16'h	5b0e;
30158	:douta	=	16'h	7c32;
30159	:douta	=	16'h	1925;
30160	:douta	=	16'h	5acc;
30161	:douta	=	16'h	a513;
30162	:douta	=	16'h	b48e;
30163	:douta	=	16'h	93ab;
30164	:douta	=	16'h	6227;
30165	:douta	=	16'h	6a67;
30166	:douta	=	16'h	5a29;
30167	:douta	=	16'h	3a6d;
30168	:douta	=	16'h	19aa;
30169	:douta	=	16'h	42ce;
30170	:douta	=	16'h	3ab0;
30171	:douta	=	16'h	6c14;
30172	:douta	=	16'h	32b0;
30173	:douta	=	16'h	528d;
30174	:douta	=	16'h	72c9;
30175	:douta	=	16'h	6a47;
30176	:douta	=	16'h	6267;
30177	:douta	=	16'h	5a48;
30178	:douta	=	16'h	5207;
30179	:douta	=	16'h	5a29;
30180	:douta	=	16'h	5a49;
30181	:douta	=	16'h	5228;
30182	:douta	=	16'h	49e8;
30183	:douta	=	16'h	4a08;
30184	:douta	=	16'h	4a08;
30185	:douta	=	16'h	49e8;
30186	:douta	=	16'h	4a28;
30187	:douta	=	16'h	4a08;
30188	:douta	=	16'h	49c7;
30189	:douta	=	16'h	41a7;
30190	:douta	=	16'h	41a7;
30191	:douta	=	16'h	3987;
30192	:douta	=	16'h	49c7;
30193	:douta	=	16'h	49c7;
30194	:douta	=	16'h	41a7;
30195	:douta	=	16'h	49e8;
30196	:douta	=	16'h	49c7;
30197	:douta	=	16'h	41a7;
30198	:douta	=	16'h	41c7;
30199	:douta	=	16'h	49e8;
30200	:douta	=	16'h	5228;
30201	:douta	=	16'h	5228;
30202	:douta	=	16'h	49c7;
30203	:douta	=	16'h	49c7;
30204	:douta	=	16'h	41a7;
30205	:douta	=	16'h	41a7;
30206	:douta	=	16'h	41a7;
30207	:douta	=	16'h	41a7;
30208	:douta	=	16'h	41c5;
30209	:douta	=	16'h	4165;
30210	:douta	=	16'h	4165;
30211	:douta	=	16'h	5b0e;
30212	:douta	=	16'h	30e2;
30213	:douta	=	16'h	3124;
30214	:douta	=	16'h	3145;
30215	:douta	=	16'h	3945;
30216	:douta	=	16'h	41c7;
30217	:douta	=	16'h	2189;
30218	:douta	=	16'h	2168;
30219	:douta	=	16'h	2188;
30220	:douta	=	16'h	29a9;
30221	:douta	=	16'h	31ea;
30222	:douta	=	16'h	2147;
30223	:douta	=	16'h	6aab;
30224	:douta	=	16'h	ac2e;
30225	:douta	=	16'h	ac2e;
30226	:douta	=	16'h	93cd;
30227	:douta	=	16'h	9bed;
30228	:douta	=	16'h	b46f;
30229	:douta	=	16'h	93cd;
30230	:douta	=	16'h	736d;
30231	:douta	=	16'h	4a8c;
30232	:douta	=	16'h	6bb0;
30233	:douta	=	16'h	6b8f;
30234	:douta	=	16'h	634e;
30235	:douta	=	16'h	6b6f;
30236	:douta	=	16'h	634e;
30237	:douta	=	16'h	6bb0;
30238	:douta	=	16'h	6bd0;
30239	:douta	=	16'h	6bd0;
30240	:douta	=	16'h	6bb0;
30241	:douta	=	16'h	73f1;
30242	:douta	=	16'h	6bd0;
30243	:douta	=	16'h	638e;
30244	:douta	=	16'h	6bcf;
30245	:douta	=	16'h	6baf;
30246	:douta	=	16'h	6bd0;
30247	:douta	=	16'h	63b0;
30248	:douta	=	16'h	5b6e;
30249	:douta	=	16'h	ff16;
30250	:douta	=	16'h	e6b5;
30251	:douta	=	16'h	e675;
30252	:douta	=	16'h	e655;
30253	:douta	=	16'h	e675;
30254	:douta	=	16'h	e675;
30255	:douta	=	16'h	ee96;
30256	:douta	=	16'h	de34;
30257	:douta	=	16'h	d5b2;
30258	:douta	=	16'h	cd92;
30259	:douta	=	16'h	c552;
30260	:douta	=	16'h	c552;
30261	:douta	=	16'h	acd1;
30262	:douta	=	16'h	9451;
30263	:douta	=	16'h	9431;
30264	:douta	=	16'h	9472;
30265	:douta	=	16'h	8c32;
30266	:douta	=	16'h	7bf2;
30267	:douta	=	16'h	738f;
30268	:douta	=	16'h	734f;
30269	:douta	=	16'h	6b2e;
30270	:douta	=	16'h	6b2f;
30271	:douta	=	16'h	7bb0;
30272	:douta	=	16'h	4985;
30273	:douta	=	16'h	7287;
30274	:douta	=	16'h	ac2a;
30275	:douta	=	16'h	c4ad;
30276	:douta	=	16'h	d5b1;
30277	:douta	=	16'h	e675;
30278	:douta	=	16'h	eeb6;
30279	:douta	=	16'h	f6b6;
30280	:douta	=	16'h	ee95;
30281	:douta	=	16'h	ee95;
30282	:douta	=	16'h	ee95;
30283	:douta	=	16'h	e635;
30284	:douta	=	16'h	d592;
30285	:douta	=	16'h	cd72;
30286	:douta	=	16'h	bd33;
30287	:douta	=	16'h	a491;
30288	:douta	=	16'h	83af;
30289	:douta	=	16'h	630d;
30290	:douta	=	16'h	62ed;
30291	:douta	=	16'h	7370;
30292	:douta	=	16'h	9453;
30293	:douta	=	16'h	9473;
30294	:douta	=	16'h	9452;
30295	:douta	=	16'h	8411;
30296	:douta	=	16'h	83f0;
30297	:douta	=	16'h	83f0;
30298	:douta	=	16'h	83cf;
30299	:douta	=	16'h	83d0;
30300	:douta	=	16'h	83af;
30301	:douta	=	16'h	7b8f;
30302	:douta	=	16'h	62cb;
30303	:douta	=	16'h	5a26;
30304	:douta	=	16'h	bc4b;
30305	:douta	=	16'h	d52e;
30306	:douta	=	16'h	ddf2;
30307	:douta	=	16'h	f6d6;
30308	:douta	=	16'h	ddf2;
30309	:douta	=	16'h	ee95;
30310	:douta	=	16'h	e634;
30311	:douta	=	16'h	ee95;
30312	:douta	=	16'h	e654;
30313	:douta	=	16'h	e653;
30314	:douta	=	16'h	e5d3;
30315	:douta	=	16'h	d591;
30316	:douta	=	16'h	cd52;
30317	:douta	=	16'h	cd73;
30318	:douta	=	16'h	c4f1;
30319	:douta	=	16'h	b4d1;
30320	:douta	=	16'h	acb1;
30321	:douta	=	16'h	a4b2;
30322	:douta	=	16'h	a493;
30323	:douta	=	16'h	9432;
30324	:douta	=	16'h	7bb0;
30325	:douta	=	16'h	7bb0;
30326	:douta	=	16'h	7b6f;
30327	:douta	=	16'h	734e;
30328	:douta	=	16'h	734e;
30329	:douta	=	16'h	732e;
30330	:douta	=	16'h	6b0e;
30331	:douta	=	16'h	732e;
30332	:douta	=	16'h	732e;
30333	:douta	=	16'h	62ed;
30334	:douta	=	16'h	6b0e;
30335	:douta	=	16'h	734e;
30336	:douta	=	16'h	5acd;
30337	:douta	=	16'h	528c;
30338	:douta	=	16'h	732c;
30339	:douta	=	16'h	ccad;
30340	:douta	=	16'h	d54f;
30341	:douta	=	16'h	de34;
30342	:douta	=	16'h	ddf3;
30343	:douta	=	16'h	bd12;
30344	:douta	=	16'h	9472;
30345	:douta	=	16'h	8c93;
30346	:douta	=	16'h	6371;
30347	:douta	=	16'h	5b11;
30348	:douta	=	16'h	428e;
30349	:douta	=	16'h	5b71;
30350	:douta	=	16'h	63b3;
30351	:douta	=	16'h	5b72;
30352	:douta	=	16'h	5331;
30353	:douta	=	16'h	4af0;
30354	:douta	=	16'h	42af;
30355	:douta	=	16'h	42af;
30356	:douta	=	16'h	4af0;
30357	:douta	=	16'h	42af;
30358	:douta	=	16'h	3a8e;
30359	:douta	=	16'h	29aa;
30360	:douta	=	16'h	322d;
30361	:douta	=	16'h	324e;
30362	:douta	=	16'h	21aa;
30363	:douta	=	16'h	3a6d;
30364	:douta	=	16'h	21a8;
30365	:douta	=	16'h	29c9;
30366	:douta	=	16'h	21c9;
30367	:douta	=	16'h	29ca;
30368	:douta	=	16'h	2168;
30369	:douta	=	16'h	10e5;
30370	:douta	=	16'h	10c4;
30371	:douta	=	16'h	10e5;
30372	:douta	=	16'h	1906;
30373	:douta	=	16'h	1906;
30374	:douta	=	16'h	10e5;
30375	:douta	=	16'h	10e5;
30376	:douta	=	16'h	10e5;
30377	:douta	=	16'h	10e5;
30378	:douta	=	16'h	10e5;
30379	:douta	=	16'h	10c5;
30380	:douta	=	16'h	1905;
30381	:douta	=	16'h	10e5;
30382	:douta	=	16'h	1926;
30383	:douta	=	16'h	18e5;
30384	:douta	=	16'h	10e5;
30385	:douta	=	16'h	10c4;
30386	:douta	=	16'h	1905;
30387	:douta	=	16'h	1905;
30388	:douta	=	16'h	18e5;
30389	:douta	=	16'h	10e5;
30390	:douta	=	16'h	10c5;
30391	:douta	=	16'h	10e5;
30392	:douta	=	16'h	10e5;
30393	:douta	=	16'h	1105;
30394	:douta	=	16'h	1906;
30395	:douta	=	16'h	29a9;
30396	:douta	=	16'h	0001;
30397	:douta	=	16'h	0000;
30398	:douta	=	16'h	2147;
30399	:douta	=	16'h	2188;
30400	:douta	=	16'h	1948;
30401	:douta	=	16'h	1926;
30402	:douta	=	16'h	324c;
30403	:douta	=	16'h	73d1;
30404	:douta	=	16'h	4aad;
30405	:douta	=	16'h	52ed;
30406	:douta	=	16'h	5b0d;
30407	:douta	=	16'h	428c;
30408	:douta	=	16'h	6b8e;
30409	:douta	=	16'h	6b90;
30410	:douta	=	16'h	94b4;
30411	:douta	=	16'h	4aed;
30412	:douta	=	16'h	530f;
30413	:douta	=	16'h	3a6b;
30414	:douta	=	16'h	1906;
30415	:douta	=	16'h	8c31;
30416	:douta	=	16'h	b4ef;
30417	:douta	=	16'h	b4cf;
30418	:douta	=	16'h	61e6;
30419	:douta	=	16'h	6247;
30420	:douta	=	16'h	6a66;
30421	:douta	=	16'h	39e9;
30422	:douta	=	16'h	1149;
30423	:douta	=	16'h	21cb;
30424	:douta	=	16'h	29eb;
30425	:douta	=	16'h	3a8e;
30426	:douta	=	16'h	63d4;
30427	:douta	=	16'h	4b31;
30428	:douta	=	16'h	3ad1;
30429	:douta	=	16'h	4209;
30430	:douta	=	16'h	6a67;
30431	:douta	=	16'h	6a69;
30432	:douta	=	16'h	6a88;
30433	:douta	=	16'h	5a28;
30434	:douta	=	16'h	5208;
30435	:douta	=	16'h	5208;
30436	:douta	=	16'h	5229;
30437	:douta	=	16'h	49e8;
30438	:douta	=	16'h	49e8;
30439	:douta	=	16'h	49e8;
30440	:douta	=	16'h	49e8;
30441	:douta	=	16'h	5229;
30442	:douta	=	16'h	49e8;
30443	:douta	=	16'h	41a7;
30444	:douta	=	16'h	41a7;
30445	:douta	=	16'h	41c7;
30446	:douta	=	16'h	41a7;
30447	:douta	=	16'h	41a7;
30448	:douta	=	16'h	41c7;
30449	:douta	=	16'h	49c7;
30450	:douta	=	16'h	49c7;
30451	:douta	=	16'h	49e8;
30452	:douta	=	16'h	49e8;
30453	:douta	=	16'h	49c7;
30454	:douta	=	16'h	49e8;
30455	:douta	=	16'h	41a7;
30456	:douta	=	16'h	49e7;
30457	:douta	=	16'h	41a7;
30458	:douta	=	16'h	41a7;
30459	:douta	=	16'h	3986;
30460	:douta	=	16'h	49e7;
30461	:douta	=	16'h	49c7;
30462	:douta	=	16'h	41c7;
30463	:douta	=	16'h	41a7;
30464	:douta	=	16'h	8b88;
30465	:douta	=	16'h	4165;
30466	:douta	=	16'h	4165;
30467	:douta	=	16'h	4a09;
30468	:douta	=	16'h	3124;
30469	:douta	=	16'h	3124;
30470	:douta	=	16'h	3145;
30471	:douta	=	16'h	3124;
30472	:douta	=	16'h	3145;
30473	:douta	=	16'h	29c9;
30474	:douta	=	16'h	2168;
30475	:douta	=	16'h	29a9;
30476	:douta	=	16'h	29c9;
30477	:douta	=	16'h	2188;
30478	:douta	=	16'h	39e9;
30479	:douta	=	16'h	7b4c;
30480	:douta	=	16'h	8b8d;
30481	:douta	=	16'h	93cd;
30482	:douta	=	16'h	8bad;
30483	:douta	=	16'h	ac4e;
30484	:douta	=	16'h	ac4e;
30485	:douta	=	16'h	9c0e;
30486	:douta	=	16'h	6b2d;
30487	:douta	=	16'h	5aed;
30488	:douta	=	16'h	634e;
30489	:douta	=	16'h	634e;
30490	:douta	=	16'h	6b8f;
30491	:douta	=	16'h	636e;
30492	:douta	=	16'h	6bb0;
30493	:douta	=	16'h	6bd0;
30494	:douta	=	16'h	6bd0;
30495	:douta	=	16'h	73d0;
30496	:douta	=	16'h	6bb0;
30497	:douta	=	16'h	638f;
30498	:douta	=	16'h	6baf;
30499	:douta	=	16'h	636f;
30500	:douta	=	16'h	638f;
30501	:douta	=	16'h	6baf;
30502	:douta	=	16'h	6bcf;
30503	:douta	=	16'h	6baf;
30504	:douta	=	16'h	6bd0;
30505	:douta	=	16'h	5b4e;
30506	:douta	=	16'h	c511;
30507	:douta	=	16'h	f6f6;
30508	:douta	=	16'h	ee96;
30509	:douta	=	16'h	ee96;
30510	:douta	=	16'h	ee96;
30511	:douta	=	16'h	de34;
30512	:douta	=	16'h	ddf3;
30513	:douta	=	16'h	cd92;
30514	:douta	=	16'h	c552;
30515	:douta	=	16'h	b4d1;
30516	:douta	=	16'h	ac91;
30517	:douta	=	16'h	a471;
30518	:douta	=	16'h	9451;
30519	:douta	=	16'h	9431;
30520	:douta	=	16'h	7bf1;
30521	:douta	=	16'h	7bf1;
30522	:douta	=	16'h	736f;
30523	:douta	=	16'h	6b4f;
30524	:douta	=	16'h	734f;
30525	:douta	=	16'h	736f;
30526	:douta	=	16'h	62cd;
30527	:douta	=	16'h	51e5;
30528	:douta	=	16'h	a42b;
30529	:douta	=	16'h	bccc;
30530	:douta	=	16'h	c50f;
30531	:douta	=	16'h	d591;
30532	:douta	=	16'h	e695;
30533	:douta	=	16'h	eeb7;
30534	:douta	=	16'h	f6b6;
30535	:douta	=	16'h	ee95;
30536	:douta	=	16'h	ee75;
30537	:douta	=	16'h	e675;
30538	:douta	=	16'h	e613;
30539	:douta	=	16'h	d5d3;
30540	:douta	=	16'h	cd73;
30541	:douta	=	16'h	c552;
30542	:douta	=	16'h	b4b2;
30543	:douta	=	16'h	9c93;
30544	:douta	=	16'h	9494;
30545	:douta	=	16'h	9494;
30546	:douta	=	16'h	9474;
30547	:douta	=	16'h	8c54;
30548	:douta	=	16'h	7390;
30549	:douta	=	16'h	6b91;
30550	:douta	=	16'h	73d1;
30551	:douta	=	16'h	7bf2;
30552	:douta	=	16'h	7391;
30553	:douta	=	16'h	6b70;
30554	:douta	=	16'h	7390;
30555	:douta	=	16'h	5aef;
30556	:douta	=	16'h	520a;
30557	:douta	=	16'h	6a48;
30558	:douta	=	16'h	936a;
30559	:douta	=	16'h	cd0e;
30560	:douta	=	16'h	e633;
30561	:douta	=	16'h	ee95;
30562	:douta	=	16'h	e612;
30563	:douta	=	16'h	d570;
30564	:douta	=	16'h	ee75;
30565	:douta	=	16'h	e654;
30566	:douta	=	16'h	e634;
30567	:douta	=	16'h	ddf3;
30568	:douta	=	16'h	e634;
30569	:douta	=	16'h	ddd2;
30570	:douta	=	16'h	d591;
30571	:douta	=	16'h	cd50;
30572	:douta	=	16'h	acb1;
30573	:douta	=	16'h	ac91;
30574	:douta	=	16'h	9431;
30575	:douta	=	16'h	9411;
30576	:douta	=	16'h	9411;
30577	:douta	=	16'h	8c11;
30578	:douta	=	16'h	83b0;
30579	:douta	=	16'h	838f;
30580	:douta	=	16'h	732c;
30581	:douta	=	16'h	734e;
30582	:douta	=	16'h	732d;
30583	:douta	=	16'h	730d;
30584	:douta	=	16'h	7b6e;
30585	:douta	=	16'h	7b4e;
30586	:douta	=	16'h	734e;
30587	:douta	=	16'h	62cd;
30588	:douta	=	16'h	5acc;
30589	:douta	=	16'h	5acb;
30590	:douta	=	16'h	836d;
30591	:douta	=	16'h	734d;
30592	:douta	=	16'h	a3ec;
30593	:douta	=	16'h	e5f2;
30594	:douta	=	16'h	f6b7;
30595	:douta	=	16'h	eeb7;
30596	:douta	=	16'h	e675;
30597	:douta	=	16'h	e655;
30598	:douta	=	16'h	cd93;
30599	:douta	=	16'h	a4b2;
30600	:douta	=	16'h	a4b3;
30601	:douta	=	16'h	9cb4;
30602	:douta	=	16'h	6b91;
30603	:douta	=	16'h	5b50;
30604	:douta	=	16'h	5310;
30605	:douta	=	16'h	6392;
30606	:douta	=	16'h	6392;
30607	:douta	=	16'h	5b72;
30608	:douta	=	16'h	5331;
30609	:douta	=	16'h	4b10;
30610	:douta	=	16'h	42af;
30611	:douta	=	16'h	4acf;
30612	:douta	=	16'h	4acf;
30613	:douta	=	16'h	426d;
30614	:douta	=	16'h	320c;
30615	:douta	=	16'h	42af;
30616	:douta	=	16'h	42cf;
30617	:douta	=	16'h	326f;
30618	:douta	=	16'h	3a2d;
30619	:douta	=	16'h	21aa;
30620	:douta	=	16'h	3a6d;
30621	:douta	=	16'h	2169;
30622	:douta	=	16'h	2189;
30623	:douta	=	16'h	10a5;
30624	:douta	=	16'h	10e5;
30625	:douta	=	16'h	1927;
30626	:douta	=	16'h	2189;
30627	:douta	=	16'h	29ca;
30628	:douta	=	16'h	21a9;
30629	:douta	=	16'h	1906;
30630	:douta	=	16'h	08c4;
30631	:douta	=	16'h	10e5;
30632	:douta	=	16'h	1905;
30633	:douta	=	16'h	10e5;
30634	:douta	=	16'h	10c5;
30635	:douta	=	16'h	18e5;
30636	:douta	=	16'h	10e5;
30637	:douta	=	16'h	10e5;
30638	:douta	=	16'h	18e5;
30639	:douta	=	16'h	1905;
30640	:douta	=	16'h	10e5;
30641	:douta	=	16'h	10c4;
30642	:douta	=	16'h	1906;
30643	:douta	=	16'h	1906;
30644	:douta	=	16'h	1905;
30645	:douta	=	16'h	18e5;
30646	:douta	=	16'h	10c5;
30647	:douta	=	16'h	1905;
30648	:douta	=	16'h	1905;
30649	:douta	=	16'h	18e5;
30650	:douta	=	16'h	1905;
30651	:douta	=	16'h	18e5;
30652	:douta	=	16'h	18e5;
30653	:douta	=	16'h	1926;
30654	:douta	=	16'h	1927;
30655	:douta	=	16'h	0884;
30656	:douta	=	16'h	08a3;
30657	:douta	=	16'h	29ca;
30658	:douta	=	16'h	7477;
30659	:douta	=	16'h	3a8d;
30660	:douta	=	16'h	530f;
30661	:douta	=	16'h	8452;
30662	:douta	=	16'h	6b90;
30663	:douta	=	16'h	5b0e;
30664	:douta	=	16'h	94d3;
30665	:douta	=	16'h	73d0;
30666	:douta	=	16'h	2166;
30667	:douta	=	16'h	4a4a;
30668	:douta	=	16'h	322a;
30669	:douta	=	16'h	b511;
30670	:douta	=	16'h	c530;
30671	:douta	=	16'h	7aa8;
30672	:douta	=	16'h	7aa6;
30673	:douta	=	16'h	7aa7;
30674	:douta	=	16'h	5229;
30675	:douta	=	16'h	29a9;
30676	:douta	=	16'h	2a4c;
30677	:douta	=	16'h	4acf;
30678	:douta	=	16'h	3a4c;
30679	:douta	=	16'h	5b51;
30680	:douta	=	16'h	3aae;
30681	:douta	=	16'h	5b50;
30682	:douta	=	16'h	3a6e;
30683	:douta	=	16'h	322d;
30684	:douta	=	16'h	222e;
30685	:douta	=	16'h	4a6c;
30686	:douta	=	16'h	72a9;
30687	:douta	=	16'h	6a68;
30688	:douta	=	16'h	6249;
30689	:douta	=	16'h	49e8;
30690	:douta	=	16'h	5228;
30691	:douta	=	16'h	5a49;
30692	:douta	=	16'h	5208;
30693	:douta	=	16'h	49e8;
30694	:douta	=	16'h	5229;
30695	:douta	=	16'h	5249;
30696	:douta	=	16'h	49e8;
30697	:douta	=	16'h	49c7;
30698	:douta	=	16'h	49e8;
30699	:douta	=	16'h	49c7;
30700	:douta	=	16'h	41a7;
30701	:douta	=	16'h	41c7;
30702	:douta	=	16'h	41a7;
30703	:douta	=	16'h	41a7;
30704	:douta	=	16'h	41a7;
30705	:douta	=	16'h	3966;
30706	:douta	=	16'h	39a6;
30707	:douta	=	16'h	49e8;
30708	:douta	=	16'h	49e8;
30709	:douta	=	16'h	41a7;
30710	:douta	=	16'h	41a7;
30711	:douta	=	16'h	49e7;
30712	:douta	=	16'h	41c7;
30713	:douta	=	16'h	3986;
30714	:douta	=	16'h	41a7;
30715	:douta	=	16'h	41a7;
30716	:douta	=	16'h	41a7;
30717	:douta	=	16'h	49c7;
30718	:douta	=	16'h	49e7;
30719	:douta	=	16'h	41a7;
30720	:douta	=	16'h	ac69;
30721	:douta	=	16'h	4185;
30722	:douta	=	16'h	4165;
30723	:douta	=	16'h	4186;
30724	:douta	=	16'h	39a6;
30725	:douta	=	16'h	3104;
30726	:douta	=	16'h	3125;
30727	:douta	=	16'h	3145;
30728	:douta	=	16'h	2925;
30729	:douta	=	16'h	320b;
30730	:douta	=	16'h	2188;
30731	:douta	=	16'h	2969;
30732	:douta	=	16'h	2168;
30733	:douta	=	16'h	2168;
30734	:douta	=	16'h	526b;
30735	:douta	=	16'h	7b2c;
30736	:douta	=	16'h	732c;
30737	:douta	=	16'h	7b2c;
30738	:douta	=	16'h	834c;
30739	:douta	=	16'h	a40d;
30740	:douta	=	16'h	9bed;
30741	:douta	=	16'h	7b6d;
30742	:douta	=	16'h	52cc;
30743	:douta	=	16'h	52cd;
30744	:douta	=	16'h	636f;
30745	:douta	=	16'h	636f;
30746	:douta	=	16'h	636e;
30747	:douta	=	16'h	634e;
30748	:douta	=	16'h	73d0;
30749	:douta	=	16'h	7411;
30750	:douta	=	16'h	7411;
30751	:douta	=	16'h	73f1;
30752	:douta	=	16'h	7c11;
30753	:douta	=	16'h	6bd0;
30754	:douta	=	16'h	63af;
30755	:douta	=	16'h	5b4e;
30756	:douta	=	16'h	5b4e;
30757	:douta	=	16'h	638e;
30758	:douta	=	16'h	6baf;
30759	:douta	=	16'h	6bcf;
30760	:douta	=	16'h	6bd0;
30761	:douta	=	16'h	63d0;
30762	:douta	=	16'h	5b4e;
30763	:douta	=	16'h	feb5;
30764	:douta	=	16'h	ee96;
30765	:douta	=	16'h	e696;
30766	:douta	=	16'h	e675;
30767	:douta	=	16'h	e655;
30768	:douta	=	16'h	d5b2;
30769	:douta	=	16'h	cd93;
30770	:douta	=	16'h	c531;
30771	:douta	=	16'h	a490;
30772	:douta	=	16'h	a471;
30773	:douta	=	16'h	9c51;
30774	:douta	=	16'h	9c72;
30775	:douta	=	16'h	9432;
30776	:douta	=	16'h	73b0;
30777	:douta	=	16'h	738f;
30778	:douta	=	16'h	738f;
30779	:douta	=	16'h	6b4f;
30780	:douta	=	16'h	734e;
30781	:douta	=	16'h	5aad;
30782	:douta	=	16'h	4187;
30783	:douta	=	16'h	a3ea;
30784	:douta	=	16'h	bcad;
30785	:douta	=	16'h	cd4f;
30786	:douta	=	16'h	ddf3;
30787	:douta	=	16'h	e654;
30788	:douta	=	16'h	f6d7;
30789	:douta	=	16'h	eeb6;
30790	:douta	=	16'h	eeb7;
30791	:douta	=	16'h	ee95;
30792	:douta	=	16'h	ee75;
30793	:douta	=	16'h	e654;
30794	:douta	=	16'h	d5d2;
30795	:douta	=	16'h	d591;
30796	:douta	=	16'h	bcf2;
30797	:douta	=	16'h	acb2;
30798	:douta	=	16'h	acd3;
30799	:douta	=	16'h	9494;
30800	:douta	=	16'h	8c54;
30801	:douta	=	16'h	8c54;
30802	:douta	=	16'h	8c54;
30803	:douta	=	16'h	8c53;
30804	:douta	=	16'h	8c73;
30805	:douta	=	16'h	7bf2;
30806	:douta	=	16'h	6b90;
30807	:douta	=	16'h	6370;
30808	:douta	=	16'h	6330;
30809	:douta	=	16'h	5b0e;
30810	:douta	=	16'h	6b2e;
30811	:douta	=	16'h	49e7;
30812	:douta	=	16'h	59e6;
30813	:douta	=	16'h	9b69;
30814	:douta	=	16'h	b42b;
30815	:douta	=	16'h	bcee;
30816	:douta	=	16'h	ff17;
30817	:douta	=	16'h	f6d7;
30818	:douta	=	16'h	eeb6;
30819	:douta	=	16'h	e654;
30820	:douta	=	16'h	ac0c;
30821	:douta	=	16'h	ee95;
30822	:douta	=	16'h	e673;
30823	:douta	=	16'h	cd30;
30824	:douta	=	16'h	ddd1;
30825	:douta	=	16'h	bcd1;
30826	:douta	=	16'h	ac70;
30827	:douta	=	16'h	b4d1;
30828	:douta	=	16'h	a472;
30829	:douta	=	16'h	a491;
30830	:douta	=	16'h	9c31;
30831	:douta	=	16'h	8c10;
30832	:douta	=	16'h	8bf1;
30833	:douta	=	16'h	8bf0;
30834	:douta	=	16'h	8c11;
30835	:douta	=	16'h	7b8f;
30836	:douta	=	16'h	7b6e;
30837	:douta	=	16'h	732d;
30838	:douta	=	16'h	730c;
30839	:douta	=	16'h	6aeb;
30840	:douta	=	16'h	734d;
30841	:douta	=	16'h	734d;
30842	:douta	=	16'h	732d;
30843	:douta	=	16'h	41ea;
30844	:douta	=	16'h	298a;
30845	:douta	=	16'h	a42f;
30846	:douta	=	16'h	c50f;
30847	:douta	=	16'h	cd71;
30848	:douta	=	16'h	b48e;
30849	:douta	=	16'h	cd72;
30850	:douta	=	16'h	e696;
30851	:douta	=	16'h	de35;
30852	:douta	=	16'h	d5f4;
30853	:douta	=	16'h	c574;
30854	:douta	=	16'h	acb3;
30855	:douta	=	16'h	9c94;
30856	:douta	=	16'h	9493;
30857	:douta	=	16'h	8c73;
30858	:douta	=	16'h	6371;
30859	:douta	=	16'h	530f;
30860	:douta	=	16'h	5330;
30861	:douta	=	16'h	5b71;
30862	:douta	=	16'h	6392;
30863	:douta	=	16'h	5351;
30864	:douta	=	16'h	5330;
30865	:douta	=	16'h	5310;
30866	:douta	=	16'h	42ae;
30867	:douta	=	16'h	428e;
30868	:douta	=	16'h	42af;
30869	:douta	=	16'h	3a4d;
30870	:douta	=	16'h	42ae;
30871	:douta	=	16'h	4ad0;
30872	:douta	=	16'h	4b10;
30873	:douta	=	16'h	31ca;
30874	:douta	=	16'h	734d;
30875	:douta	=	16'h	218a;
30876	:douta	=	16'h	4b10;
30877	:douta	=	16'h	29ca;
30878	:douta	=	16'h	324d;
30879	:douta	=	16'h	2988;
30880	:douta	=	16'h	2147;
30881	:douta	=	16'h	10e5;
30882	:douta	=	16'h	1084;
30883	:douta	=	16'h	10e5;
30884	:douta	=	16'h	2147;
30885	:douta	=	16'h	29ca;
30886	:douta	=	16'h	2167;
30887	:douta	=	16'h	1926;
30888	:douta	=	16'h	10e5;
30889	:douta	=	16'h	10e5;
30890	:douta	=	16'h	10e5;
30891	:douta	=	16'h	18e5;
30892	:douta	=	16'h	18e5;
30893	:douta	=	16'h	10e5;
30894	:douta	=	16'h	1905;
30895	:douta	=	16'h	10c4;
30896	:douta	=	16'h	10e5;
30897	:douta	=	16'h	10a4;
30898	:douta	=	16'h	1905;
30899	:douta	=	16'h	18e5;
30900	:douta	=	16'h	10e5;
30901	:douta	=	16'h	10e5;
30902	:douta	=	16'h	10e5;
30903	:douta	=	16'h	1926;
30904	:douta	=	16'h	1905;
30905	:douta	=	16'h	1926;
30906	:douta	=	16'h	1905;
30907	:douta	=	16'h	1905;
30908	:douta	=	16'h	1905;
30909	:douta	=	16'h	10e5;
30910	:douta	=	16'h	1926;
30911	:douta	=	16'h	2147;
30912	:douta	=	16'h	0021;
30913	:douta	=	16'h	0863;
30914	:douta	=	16'h	530f;
30915	:douta	=	16'h	6c14;
30916	:douta	=	16'h	6391;
30917	:douta	=	16'h	6370;
30918	:douta	=	16'h	7411;
30919	:douta	=	16'h	636f;
30920	:douta	=	16'h	6b8e;
30921	:douta	=	16'h	52cb;
30922	:douta	=	16'h	4aab;
30923	:douta	=	16'h	a4d2;
30924	:douta	=	16'h	c5b3;
30925	:douta	=	16'h	ac2b;
30926	:douta	=	16'h	7ac7;
30927	:douta	=	16'h	7aa7;
30928	:douta	=	16'h	6227;
30929	:douta	=	16'h	628b;
30930	:douta	=	16'h	2a0c;
30931	:douta	=	16'h	2a2c;
30932	:douta	=	16'h	3aae;
30933	:douta	=	16'h	42ad;
30934	:douta	=	16'h	4aee;
30935	:douta	=	16'h	4acf;
30936	:douta	=	16'h	42ad;
30937	:douta	=	16'h	6371;
30938	:douta	=	16'h	3a4c;
30939	:douta	=	16'h	31eb;
30940	:douta	=	16'h	4b52;
30941	:douta	=	16'h	5b2f;
30942	:douta	=	16'h	6a88;
30943	:douta	=	16'h	6a69;
30944	:douta	=	16'h	5228;
30945	:douta	=	16'h	5228;
30946	:douta	=	16'h	5228;
30947	:douta	=	16'h	5228;
30948	:douta	=	16'h	49e7;
30949	:douta	=	16'h	49e8;
30950	:douta	=	16'h	5249;
30951	:douta	=	16'h	5249;
30952	:douta	=	16'h	5209;
30953	:douta	=	16'h	49c7;
30954	:douta	=	16'h	49c7;
30955	:douta	=	16'h	41c7;
30956	:douta	=	16'h	4186;
30957	:douta	=	16'h	41a7;
30958	:douta	=	16'h	41c7;
30959	:douta	=	16'h	41c7;
30960	:douta	=	16'h	41c7;
30961	:douta	=	16'h	3986;
30962	:douta	=	16'h	3987;
30963	:douta	=	16'h	49c7;
30964	:douta	=	16'h	49c8;
30965	:douta	=	16'h	49e8;
30966	:douta	=	16'h	49e7;
30967	:douta	=	16'h	49c7;
30968	:douta	=	16'h	49e7;
30969	:douta	=	16'h	41a7;
30970	:douta	=	16'h	3986;
30971	:douta	=	16'h	41a7;
30972	:douta	=	16'h	49e7;
30973	:douta	=	16'h	49c7;
30974	:douta	=	16'h	49e7;
30975	:douta	=	16'h	49e7;
30976	:douta	=	16'h	e58b;
30977	:douta	=	16'h	28e5;
30978	:douta	=	16'h	4165;
30979	:douta	=	16'h	30e2;
30980	:douta	=	16'h	528b;
30981	:douta	=	16'h	28c2;
30982	:douta	=	16'h	3124;
30983	:douta	=	16'h	3145;
30984	:douta	=	16'h	2904;
30985	:douta	=	16'h	31ea;
30986	:douta	=	16'h	2168;
30987	:douta	=	16'h	2988;
30988	:douta	=	16'h	21a8;
30989	:douta	=	16'h	1947;
30990	:douta	=	16'h	5aab;
30991	:douta	=	16'h	62ac;
30992	:douta	=	16'h	6acc;
30993	:douta	=	16'h	6aec;
30994	:douta	=	16'h	7b4d;
30995	:douta	=	16'h	730c;
30996	:douta	=	16'h	836d;
30997	:douta	=	16'h	528b;
30998	:douta	=	16'h	4a8c;
30999	:douta	=	16'h	52cc;
31000	:douta	=	16'h	5b0e;
31001	:douta	=	16'h	634f;
31002	:douta	=	16'h	73d0;
31003	:douta	=	16'h	6bb0;
31004	:douta	=	16'h	73d0;
31005	:douta	=	16'h	6b8f;
31006	:douta	=	16'h	6bb0;
31007	:douta	=	16'h	6bb0;
31008	:douta	=	16'h	6bd0;
31009	:douta	=	16'h	73f0;
31010	:douta	=	16'h	7411;
31011	:douta	=	16'h	6baf;
31012	:douta	=	16'h	638f;
31013	:douta	=	16'h	6baf;
31014	:douta	=	16'h	638f;
31015	:douta	=	16'h	6bcf;
31016	:douta	=	16'h	6bd0;
31017	:douta	=	16'h	6baf;
31018	:douta	=	16'h	73f0;
31019	:douta	=	16'h	534e;
31020	:douta	=	16'h	d572;
31021	:douta	=	16'h	feb5;
31022	:douta	=	16'h	de35;
31023	:douta	=	16'h	e634;
31024	:douta	=	16'h	ddf4;
31025	:douta	=	16'h	b511;
31026	:douta	=	16'h	ac91;
31027	:douta	=	16'h	acb2;
31028	:douta	=	16'h	a470;
31029	:douta	=	16'h	a492;
31030	:douta	=	16'h	9432;
31031	:douta	=	16'h	83d1;
31032	:douta	=	16'h	736f;
31033	:douta	=	16'h	7370;
31034	:douta	=	16'h	734e;
31035	:douta	=	16'h	7370;
31036	:douta	=	16'h	528c;
31037	:douta	=	16'h	8328;
31038	:douta	=	16'h	bcaa;
31039	:douta	=	16'h	cd2f;
31040	:douta	=	16'h	e633;
31041	:douta	=	16'h	e675;
31042	:douta	=	16'h	eeb7;
31043	:douta	=	16'h	eeb7;
31044	:douta	=	16'h	eeb7;
31045	:douta	=	16'h	eeb7;
31046	:douta	=	16'h	eeb6;
31047	:douta	=	16'h	e675;
31048	:douta	=	16'h	de13;
31049	:douta	=	16'h	d5f3;
31050	:douta	=	16'h	c532;
31051	:douta	=	16'h	b4d2;
31052	:douta	=	16'h	9473;
31053	:douta	=	16'h	8c94;
31054	:douta	=	16'h	8c74;
31055	:douta	=	16'h	8c74;
31056	:douta	=	16'h	8c95;
31057	:douta	=	16'h	8454;
31058	:douta	=	16'h	8413;
31059	:douta	=	16'h	83f1;
31060	:douta	=	16'h	7b90;
31061	:douta	=	16'h	6b4e;
31062	:douta	=	16'h	734f;
31063	:douta	=	16'h	6b0e;
31064	:douta	=	16'h	5acd;
31065	:douta	=	16'h	4a6b;
31066	:douta	=	16'h	4164;
31067	:douta	=	16'h	9369;
31068	:douta	=	16'h	b42c;
31069	:douta	=	16'h	ee74;
31070	:douta	=	16'h	e654;
31071	:douta	=	16'h	f6f7;
31072	:douta	=	16'h	a40b;
31073	:douta	=	16'h	d550;
31074	:douta	=	16'h	ee95;
31075	:douta	=	16'h	ee95;
31076	:douta	=	16'h	ee95;
31077	:douta	=	16'h	832b;
31078	:douta	=	16'h	b4ae;
31079	:douta	=	16'h	bcf0;
31080	:douta	=	16'h	bcd0;
31081	:douta	=	16'h	ac90;
31082	:douta	=	16'h	9431;
31083	:douta	=	16'h	9411;
31084	:douta	=	16'h	93f0;
31085	:douta	=	16'h	8bcf;
31086	:douta	=	16'h	8bf0;
31087	:douta	=	16'h	83d0;
31088	:douta	=	16'h	7b8f;
31089	:douta	=	16'h	7b6e;
31090	:douta	=	16'h	734d;
31091	:douta	=	16'h	7b6e;
31092	:douta	=	16'h	7b6d;
31093	:douta	=	16'h	7b2d;
31094	:douta	=	16'h	62cb;
31095	:douta	=	16'h	62cc;
31096	:douta	=	16'h	62ab;
31097	:douta	=	16'h	730c;
31098	:douta	=	16'h	9c0e;
31099	:douta	=	16'h	e613;
31100	:douta	=	16'h	f675;
31101	:douta	=	16'h	e656;
31102	:douta	=	16'h	eeb7;
31103	:douta	=	16'h	eeb7;
31104	:douta	=	16'h	e696;
31105	:douta	=	16'h	e656;
31106	:douta	=	16'h	de15;
31107	:douta	=	16'h	d5d5;
31108	:douta	=	16'h	cdb4;
31109	:douta	=	16'h	b554;
31110	:douta	=	16'h	b514;
31111	:douta	=	16'h	9cd4;
31112	:douta	=	16'h	9cb4;
31113	:douta	=	16'h	94b4;
31114	:douta	=	16'h	73d2;
31115	:douta	=	16'h	6371;
31116	:douta	=	16'h	5b30;
31117	:douta	=	16'h	6371;
31118	:douta	=	16'h	5b51;
31119	:douta	=	16'h	530f;
31120	:douta	=	16'h	4acf;
31121	:douta	=	16'h	4aaf;
31122	:douta	=	16'h	4aef;
31123	:douta	=	16'h	4acf;
31124	:douta	=	16'h	5330;
31125	:douta	=	16'h	5b51;
31126	:douta	=	16'h	52f0;
31127	:douta	=	16'h	326f;
31128	:douta	=	16'h	31ec;
31129	:douta	=	16'h	bd54;
31130	:douta	=	16'h	6c15;
31131	:douta	=	16'h	2a2c;
31132	:douta	=	16'h	5331;
31133	:douta	=	16'h	42af;
31134	:douta	=	16'h	3a8e;
31135	:douta	=	16'h	42af;
31136	:douta	=	16'h	322c;
31137	:douta	=	16'h	21ca;
31138	:douta	=	16'h	21a9;
31139	:douta	=	16'h	2168;
31140	:douta	=	16'h	2147;
31141	:douta	=	16'h	10e5;
31142	:douta	=	16'h	1905;
31143	:douta	=	16'h	1906;
31144	:douta	=	16'h	29ea;
31145	:douta	=	16'h	21a9;
31146	:douta	=	16'h	21a9;
31147	:douta	=	16'h	2147;
31148	:douta	=	16'h	10e5;
31149	:douta	=	16'h	10e5;
31150	:douta	=	16'h	0884;
31151	:douta	=	16'h	10e5;
31152	:douta	=	16'h	10c4;
31153	:douta	=	16'h	10c5;
31154	:douta	=	16'h	10e5;
31155	:douta	=	16'h	10e5;
31156	:douta	=	16'h	10e5;
31157	:douta	=	16'h	10c5;
31158	:douta	=	16'h	10e5;
31159	:douta	=	16'h	10e5;
31160	:douta	=	16'h	10e5;
31161	:douta	=	16'h	10e5;
31162	:douta	=	16'h	10e5;
31163	:douta	=	16'h	1905;
31164	:douta	=	16'h	10e5;
31165	:douta	=	16'h	10c5;
31166	:douta	=	16'h	10c4;
31167	:douta	=	16'h	10c5;
31168	:douta	=	16'h	1925;
31169	:douta	=	16'h	10e5;
31170	:douta	=	16'h	0063;
31171	:douta	=	16'h	0000;
31172	:douta	=	16'h	2187;
31173	:douta	=	16'h	10a4;
31174	:douta	=	16'h	1927;
31175	:douta	=	16'h	2988;
31176	:douta	=	16'h	93ef;
31177	:douta	=	16'h	ad10;
31178	:douta	=	16'h	c50f;
31179	:douta	=	16'h	7a67;
31180	:douta	=	16'h	82c7;
31181	:douta	=	16'h	8b08;
31182	:douta	=	16'h	6289;
31183	:douta	=	16'h	21cb;
31184	:douta	=	16'h	42ae;
31185	:douta	=	16'h	3a2d;
31186	:douta	=	16'h	3a6d;
31187	:douta	=	16'h	322c;
31188	:douta	=	16'h	530f;
31189	:douta	=	16'h	4b0f;
31190	:douta	=	16'h	2a0b;
31191	:douta	=	16'h	6bb2;
31192	:douta	=	16'h	530f;
31193	:douta	=	16'h	4b10;
31194	:douta	=	16'h	42cf;
31195	:douta	=	16'h	42f0;
31196	:douta	=	16'h	4b11;
31197	:douta	=	16'h	3aaf;
31198	:douta	=	16'h	7287;
31199	:douta	=	16'h	6289;
31200	:douta	=	16'h	5a48;
31201	:douta	=	16'h	5249;
31202	:douta	=	16'h	5228;
31203	:douta	=	16'h	5208;
31204	:douta	=	16'h	5208;
31205	:douta	=	16'h	5228;
31206	:douta	=	16'h	49e8;
31207	:douta	=	16'h	49e8;
31208	:douta	=	16'h	49c7;
31209	:douta	=	16'h	49c7;
31210	:douta	=	16'h	41c7;
31211	:douta	=	16'h	41a7;
31212	:douta	=	16'h	49e8;
31213	:douta	=	16'h	41c7;
31214	:douta	=	16'h	41c7;
31215	:douta	=	16'h	49c7;
31216	:douta	=	16'h	49c7;
31217	:douta	=	16'h	49e7;
31218	:douta	=	16'h	3986;
31219	:douta	=	16'h	3966;
31220	:douta	=	16'h	41a7;
31221	:douta	=	16'h	41a6;
31222	:douta	=	16'h	3986;
31223	:douta	=	16'h	41a7;
31224	:douta	=	16'h	41a6;
31225	:douta	=	16'h	41c7;
31226	:douta	=	16'h	49c7;
31227	:douta	=	16'h	49c7;
31228	:douta	=	16'h	41c7;
31229	:douta	=	16'h	49c7;
31230	:douta	=	16'h	41a7;
31231	:douta	=	16'h	41a7;
31232	:douta	=	16'h	f5cb;
31233	:douta	=	16'h	20c4;
31234	:douta	=	16'h	4185;
31235	:douta	=	16'h	38e3;
31236	:douta	=	16'h	52ed;
31237	:douta	=	16'h	30e3;
31238	:douta	=	16'h	3124;
31239	:douta	=	16'h	3124;
31240	:douta	=	16'h	2904;
31241	:douta	=	16'h	320b;
31242	:douta	=	16'h	2168;
31243	:douta	=	16'h	2188;
31244	:douta	=	16'h	2188;
31245	:douta	=	16'h	2168;
31246	:douta	=	16'h	5aac;
31247	:douta	=	16'h	5a8b;
31248	:douta	=	16'h	62cc;
31249	:douta	=	16'h	62cc;
31250	:douta	=	16'h	72ec;
31251	:douta	=	16'h	6aec;
31252	:douta	=	16'h	730d;
31253	:douta	=	16'h	4a8c;
31254	:douta	=	16'h	4a8b;
31255	:douta	=	16'h	4aad;
31256	:douta	=	16'h	52ee;
31257	:douta	=	16'h	5b0d;
31258	:douta	=	16'h	636f;
31259	:douta	=	16'h	6b8f;
31260	:douta	=	16'h	6bb0;
31261	:douta	=	16'h	6bd0;
31262	:douta	=	16'h	6bb0;
31263	:douta	=	16'h	6bd0;
31264	:douta	=	16'h	7411;
31265	:douta	=	16'h	7411;
31266	:douta	=	16'h	73f1;
31267	:douta	=	16'h	6bcf;
31268	:douta	=	16'h	638f;
31269	:douta	=	16'h	638f;
31270	:douta	=	16'h	6baf;
31271	:douta	=	16'h	638f;
31272	:douta	=	16'h	6bcf;
31273	:douta	=	16'h	638f;
31274	:douta	=	16'h	6bf0;
31275	:douta	=	16'h	6bd0;
31276	:douta	=	16'h	5b0d;
31277	:douta	=	16'h	b4d2;
31278	:douta	=	16'h	e634;
31279	:douta	=	16'h	d5d3;
31280	:douta	=	16'h	d5b2;
31281	:douta	=	16'h	a470;
31282	:douta	=	16'h	a450;
31283	:douta	=	16'h	a4b1;
31284	:douta	=	16'h	b4d2;
31285	:douta	=	16'h	83f0;
31286	:douta	=	16'h	6b2f;
31287	:douta	=	16'h	6b2e;
31288	:douta	=	16'h	7370;
31289	:douta	=	16'h	734f;
31290	:douta	=	16'h	734f;
31291	:douta	=	16'h	420a;
31292	:douta	=	16'h	4187;
31293	:douta	=	16'h	cd2d;
31294	:douta	=	16'h	cd2e;
31295	:douta	=	16'h	d5b0;
31296	:douta	=	16'h	eeb6;
31297	:douta	=	16'h	eeb6;
31298	:douta	=	16'h	eed7;
31299	:douta	=	16'h	eeb6;
31300	:douta	=	16'h	eeb6;
31301	:douta	=	16'h	ee97;
31302	:douta	=	16'h	ee96;
31303	:douta	=	16'h	e634;
31304	:douta	=	16'h	d5f3;
31305	:douta	=	16'h	cd93;
31306	:douta	=	16'h	bcf2;
31307	:douta	=	16'h	acb3;
31308	:douta	=	16'h	9cb4;
31309	:douta	=	16'h	94b5;
31310	:douta	=	16'h	8455;
31311	:douta	=	16'h	8455;
31312	:douta	=	16'h	8454;
31313	:douta	=	16'h	7c12;
31314	:douta	=	16'h	7bd1;
31315	:douta	=	16'h	7bd1;
31316	:douta	=	16'h	7b90;
31317	:douta	=	16'h	6b4f;
31318	:douta	=	16'h	62ed;
31319	:douta	=	16'h	632e;
31320	:douta	=	16'h	528b;
31321	:douta	=	16'h	3145;
31322	:douta	=	16'h	72a8;
31323	:douta	=	16'h	c4ac;
31324	:douta	=	16'h	cd0e;
31325	:douta	=	16'h	d5b1;
31326	:douta	=	16'h	eed7;
31327	:douta	=	16'h	ee95;
31328	:douta	=	16'h	d591;
31329	:douta	=	16'h	d591;
31330	:douta	=	16'h	e654;
31331	:douta	=	16'h	ee95;
31332	:douta	=	16'h	ee94;
31333	:douta	=	16'h	a42e;
31334	:douta	=	16'h	93cd;
31335	:douta	=	16'h	ac70;
31336	:douta	=	16'h	ac90;
31337	:douta	=	16'h	ac90;
31338	:douta	=	16'h	8c10;
31339	:douta	=	16'h	8bf0;
31340	:douta	=	16'h	838e;
31341	:douta	=	16'h	83cf;
31342	:douta	=	16'h	838e;
31343	:douta	=	16'h	7b4d;
31344	:douta	=	16'h	730c;
31345	:douta	=	16'h	730c;
31346	:douta	=	16'h	730c;
31347	:douta	=	16'h	732c;
31348	:douta	=	16'h	838e;
31349	:douta	=	16'h	8bce;
31350	:douta	=	16'h	7b4d;
31351	:douta	=	16'h	6acb;
31352	:douta	=	16'h	628b;
31353	:douta	=	16'h	cd52;
31354	:douta	=	16'h	ee75;
31355	:douta	=	16'h	d5d4;
31356	:douta	=	16'h	de15;
31357	:douta	=	16'h	e697;
31358	:douta	=	16'h	eeb8;
31359	:douta	=	16'h	ee97;
31360	:douta	=	16'h	d5f5;
31361	:douta	=	16'h	cdb4;
31362	:douta	=	16'h	bd54;
31363	:douta	=	16'h	ad14;
31364	:douta	=	16'h	ad15;
31365	:douta	=	16'h	a4d5;
31366	:douta	=	16'h	a4b4;
31367	:douta	=	16'h	9c94;
31368	:douta	=	16'h	9494;
31369	:douta	=	16'h	8c73;
31370	:douta	=	16'h	7bf2;
31371	:douta	=	16'h	73b1;
31372	:douta	=	16'h	6350;
31373	:douta	=	16'h	5b50;
31374	:douta	=	16'h	5b30;
31375	:douta	=	16'h	530f;
31376	:douta	=	16'h	4acf;
31377	:douta	=	16'h	5310;
31378	:douta	=	16'h	532f;
31379	:douta	=	16'h	5330;
31380	:douta	=	16'h	5b50;
31381	:douta	=	16'h	5330;
31382	:douta	=	16'h	4af0;
31383	:douta	=	16'h	630e;
31384	:douta	=	16'h	c4f0;
31385	:douta	=	16'h	7434;
31386	:douta	=	16'h	5bb2;
31387	:douta	=	16'h	3a6e;
31388	:douta	=	16'h	63b2;
31389	:douta	=	16'h	4acf;
31390	:douta	=	16'h	42af;
31391	:douta	=	16'h	4af0;
31392	:douta	=	16'h	328e;
31393	:douta	=	16'h	324d;
31394	:douta	=	16'h	322c;
31395	:douta	=	16'h	2189;
31396	:douta	=	16'h	21aa;
31397	:douta	=	16'h	1926;
31398	:douta	=	16'h	1927;
31399	:douta	=	16'h	1927;
31400	:douta	=	16'h	1947;
31401	:douta	=	16'h	1906;
31402	:douta	=	16'h	3aaf;
31403	:douta	=	16'h	2a2c;
31404	:douta	=	16'h	2148;
31405	:douta	=	16'h	2127;
31406	:douta	=	16'h	2167;
31407	:douta	=	16'h	29a9;
31408	:douta	=	16'h	29a9;
31409	:douta	=	16'h	1926;
31410	:douta	=	16'h	18e5;
31411	:douta	=	16'h	10e4;
31412	:douta	=	16'h	10c4;
31413	:douta	=	16'h	10e4;
31414	:douta	=	16'h	1947;
31415	:douta	=	16'h	1926;
31416	:douta	=	16'h	10c5;
31417	:douta	=	16'h	1906;
31418	:douta	=	16'h	18e5;
31419	:douta	=	16'h	18e5;
31420	:douta	=	16'h	10e5;
31421	:douta	=	16'h	10c5;
31422	:douta	=	16'h	10c4;
31423	:douta	=	16'h	10a4;
31424	:douta	=	16'h	1905;
31425	:douta	=	16'h	10c5;
31426	:douta	=	16'h	10e5;
31427	:douta	=	16'h	0042;
31428	:douta	=	16'h	0000;
31429	:douta	=	16'h	2167;
31430	:douta	=	16'h	2146;
31431	:douta	=	16'h	10c6;
31432	:douta	=	16'h	cd92;
31433	:douta	=	16'h	d54f;
31434	:douta	=	16'h	8267;
31435	:douta	=	16'h	9327;
31436	:douta	=	16'h	82e9;
31437	:douta	=	16'h	422a;
31438	:douta	=	16'h	324d;
31439	:douta	=	16'h	6391;
31440	:douta	=	16'h	29cb;
31441	:douta	=	16'h	29cb;
31442	:douta	=	16'h	4aad;
31443	:douta	=	16'h	29eb;
31444	:douta	=	16'h	5b50;
31445	:douta	=	16'h	530f;
31446	:douta	=	16'h	4b0f;
31447	:douta	=	16'h	5330;
31448	:douta	=	16'h	5b71;
31449	:douta	=	16'h	324d;
31450	:douta	=	16'h	328f;
31451	:douta	=	16'h	4b10;
31452	:douta	=	16'h	6bf4;
31453	:douta	=	16'h	32af;
31454	:douta	=	16'h	6acc;
31455	:douta	=	16'h	6268;
31456	:douta	=	16'h	6289;
31457	:douta	=	16'h	5249;
31458	:douta	=	16'h	5229;
31459	:douta	=	16'h	5228;
31460	:douta	=	16'h	5249;
31461	:douta	=	16'h	5249;
31462	:douta	=	16'h	49e8;
31463	:douta	=	16'h	41a7;
31464	:douta	=	16'h	41a7;
31465	:douta	=	16'h	41a7;
31466	:douta	=	16'h	41a7;
31467	:douta	=	16'h	41a7;
31468	:douta	=	16'h	41c7;
31469	:douta	=	16'h	49c7;
31470	:douta	=	16'h	41c7;
31471	:douta	=	16'h	41c7;
31472	:douta	=	16'h	41a7;
31473	:douta	=	16'h	41c7;
31474	:douta	=	16'h	41a6;
31475	:douta	=	16'h	41a7;
31476	:douta	=	16'h	41c7;
31477	:douta	=	16'h	41a7;
31478	:douta	=	16'h	39a6;
31479	:douta	=	16'h	41a6;
31480	:douta	=	16'h	41c7;
31481	:douta	=	16'h	41a7;
31482	:douta	=	16'h	41c7;
31483	:douta	=	16'h	41a7;
31484	:douta	=	16'h	49c7;
31485	:douta	=	16'h	49e8;
31486	:douta	=	16'h	49c8;
31487	:douta	=	16'h	41a7;
31488	:douta	=	16'h	ed8b;
31489	:douta	=	16'h	41a5;
31490	:douta	=	16'h	3124;
31491	:douta	=	16'h	3944;
31492	:douta	=	16'h	634f;
31493	:douta	=	16'h	41c7;
31494	:douta	=	16'h	3144;
31495	:douta	=	16'h	3124;
31496	:douta	=	16'h	3124;
31497	:douta	=	16'h	424b;
31498	:douta	=	16'h	29ca;
31499	:douta	=	16'h	29a8;
31500	:douta	=	16'h	29a9;
31501	:douta	=	16'h	2989;
31502	:douta	=	16'h	52ac;
31503	:douta	=	16'h	4a4a;
31504	:douta	=	16'h	5a8b;
31505	:douta	=	16'h	5a8b;
31506	:douta	=	16'h	526a;
31507	:douta	=	16'h	5aac;
31508	:douta	=	16'h	5acd;
31509	:douta	=	16'h	52cc;
31510	:douta	=	16'h	426b;
31511	:douta	=	16'h	52cd;
31512	:douta	=	16'h	530e;
31513	:douta	=	16'h	5b2e;
31514	:douta	=	16'h	634e;
31515	:douta	=	16'h	636f;
31516	:douta	=	16'h	6bd0;
31517	:douta	=	16'h	73f1;
31518	:douta	=	16'h	73f1;
31519	:douta	=	16'h	6bd0;
31520	:douta	=	16'h	73f0;
31521	:douta	=	16'h	6bf1;
31522	:douta	=	16'h	73f1;
31523	:douta	=	16'h	6bcf;
31524	:douta	=	16'h	6bd0;
31525	:douta	=	16'h	638f;
31526	:douta	=	16'h	6baf;
31527	:douta	=	16'h	638f;
31528	:douta	=	16'h	6baf;
31529	:douta	=	16'h	6bef;
31530	:douta	=	16'h	6bcf;
31531	:douta	=	16'h	6bd0;
31532	:douta	=	16'h	634e;
31533	:douta	=	16'h	5b6e;
31534	:douta	=	16'h	736e;
31535	:douta	=	16'h	c531;
31536	:douta	=	16'h	cd52;
31537	:douta	=	16'h	a490;
31538	:douta	=	16'h	ac90;
31539	:douta	=	16'h	8bcf;
31540	:douta	=	16'h	8bf0;
31541	:douta	=	16'h	9431;
31542	:douta	=	16'h	7bd0;
31543	:douta	=	16'h	7b6f;
31544	:douta	=	16'h	734e;
31545	:douta	=	16'h	732e;
31546	:douta	=	16'h	3a2b;
31547	:douta	=	16'h	9b6a;
31548	:douta	=	16'h	bc4b;
31549	:douta	=	16'h	ee76;
31550	:douta	=	16'h	d5d2;
31551	:douta	=	16'h	ee96;
31552	:douta	=	16'h	eeb6;
31553	:douta	=	16'h	f6d7;
31554	:douta	=	16'h	eeb7;
31555	:douta	=	16'h	eeb7;
31556	:douta	=	16'h	e676;
31557	:douta	=	16'h	e675;
31558	:douta	=	16'h	e634;
31559	:douta	=	16'h	d5b3;
31560	:douta	=	16'h	bd32;
31561	:douta	=	16'h	a4b3;
31562	:douta	=	16'h	9c93;
31563	:douta	=	16'h	9474;
31564	:douta	=	16'h	8c53;
31565	:douta	=	16'h	8453;
31566	:douta	=	16'h	8454;
31567	:douta	=	16'h	7bd1;
31568	:douta	=	16'h	7390;
31569	:douta	=	16'h	6b4f;
31570	:douta	=	16'h	6b4e;
31571	:douta	=	16'h	6b2e;
31572	:douta	=	16'h	6b0e;
31573	:douta	=	16'h	630d;
31574	:douta	=	16'h	62cd;
31575	:douta	=	16'h	49a7;
31576	:douta	=	16'h	7287;
31577	:douta	=	16'h	ac2c;
31578	:douta	=	16'h	8b28;
31579	:douta	=	16'h	ee75;
31580	:douta	=	16'h	ee75;
31581	:douta	=	16'h	ddf3;
31582	:douta	=	16'h	bcac;
31583	:douta	=	16'h	f6d7;
31584	:douta	=	16'h	a470;
31585	:douta	=	16'h	730b;
31586	:douta	=	16'h	ee54;
31587	:douta	=	16'h	e674;
31588	:douta	=	16'h	cd71;
31589	:douta	=	16'h	acd1;
31590	:douta	=	16'h	a490;
31591	:douta	=	16'h	a471;
31592	:douta	=	16'h	9431;
31593	:douta	=	16'h	7bd0;
31594	:douta	=	16'h	83cf;
31595	:douta	=	16'h	7baf;
31596	:douta	=	16'h	734e;
31597	:douta	=	16'h	6b2d;
31598	:douta	=	16'h	730d;
31599	:douta	=	16'h	7b6e;
31600	:douta	=	16'h	838e;
31601	:douta	=	16'h	732d;
31602	:douta	=	16'h	62aa;
31603	:douta	=	16'h	5249;
31604	:douta	=	16'h	41e8;
31605	:douta	=	16'h	39a8;
31606	:douta	=	16'h	832b;
31607	:douta	=	16'h	bc8f;
31608	:douta	=	16'h	c531;
31609	:douta	=	16'h	ac6d;
31610	:douta	=	16'h	ac6d;
31611	:douta	=	16'h	d5d4;
31612	:douta	=	16'h	c573;
31613	:douta	=	16'h	cd94;
31614	:douta	=	16'h	d5d4;
31615	:douta	=	16'h	cdd5;
31616	:douta	=	16'h	cdb5;
31617	:douta	=	16'h	c575;
31618	:douta	=	16'h	bd55;
31619	:douta	=	16'h	b535;
31620	:douta	=	16'h	ad15;
31621	:douta	=	16'h	9cb5;
31622	:douta	=	16'h	9cd5;
31623	:douta	=	16'h	9494;
31624	:douta	=	16'h	8c93;
31625	:douta	=	16'h	9494;
31626	:douta	=	16'h	8433;
31627	:douta	=	16'h	73d1;
31628	:douta	=	16'h	73b1;
31629	:douta	=	16'h	6350;
31630	:douta	=	16'h	6350;
31631	:douta	=	16'h	5b30;
31632	:douta	=	16'h	5b0f;
31633	:douta	=	16'h	4aae;
31634	:douta	=	16'h	52ee;
31635	:douta	=	16'h	4ace;
31636	:douta	=	16'h	4ace;
31637	:douta	=	16'h	632f;
31638	:douta	=	16'h	cd11;
31639	:douta	=	16'h	ddd3;
31640	:douta	=	16'h	ee35;
31641	:douta	=	16'h	7c74;
31642	:douta	=	16'h	6bf3;
31643	:douta	=	16'h	5350;
31644	:douta	=	16'h	6bd3;
31645	:douta	=	16'h	5b72;
31646	:douta	=	16'h	5310;
31647	:douta	=	16'h	4af0;
31648	:douta	=	16'h	3a8e;
31649	:douta	=	16'h	322c;
31650	:douta	=	16'h	322c;
31651	:douta	=	16'h	29ca;
31652	:douta	=	16'h	29ca;
31653	:douta	=	16'h	2189;
31654	:douta	=	16'h	1947;
31655	:douta	=	16'h	1927;
31656	:douta	=	16'h	29ca;
31657	:douta	=	16'h	21aa;
31658	:douta	=	16'h	29cb;
31659	:douta	=	16'h	42d0;
31660	:douta	=	16'h	29cb;
31661	:douta	=	16'h	1968;
31662	:douta	=	16'h	10e5;
31663	:douta	=	16'h	2147;
31664	:douta	=	16'h	1927;
31665	:douta	=	16'h	2128;
31666	:douta	=	16'h	2168;
31667	:douta	=	16'h	2169;
31668	:douta	=	16'h	29aa;
31669	:douta	=	16'h	29eb;
31670	:douta	=	16'h	29eb;
31671	:douta	=	16'h	29aa;
31672	:douta	=	16'h	1906;
31673	:douta	=	16'h	0863;
31674	:douta	=	16'h	10c3;
31675	:douta	=	16'h	10e5;
31676	:douta	=	16'h	10e5;
31677	:douta	=	16'h	10c5;
31678	:douta	=	16'h	10e5;
31679	:douta	=	16'h	10e5;
31680	:douta	=	16'h	1905;
31681	:douta	=	16'h	10c5;
31682	:douta	=	16'h	0884;
31683	:douta	=	16'h	10c4;
31684	:douta	=	16'h	1905;
31685	:douta	=	16'h	2126;
31686	:douta	=	16'h	08a3;
31687	:douta	=	16'h	10e5;
31688	:douta	=	16'h	08c6;
31689	:douta	=	16'h	10e6;
31690	:douta	=	16'h	7b2b;
31691	:douta	=	16'h	3a4d;
31692	:douta	=	16'h	320c;
31693	:douta	=	16'h	532f;
31694	:douta	=	16'h	7413;
31695	:douta	=	16'h	428e;
31696	:douta	=	16'h	320c;
31697	:douta	=	16'h	3a4d;
31698	:douta	=	16'h	4aad;
31699	:douta	=	16'h	7c13;
31700	:douta	=	16'h	5b71;
31701	:douta	=	16'h	5b50;
31702	:douta	=	16'h	5b71;
31703	:douta	=	16'h	5330;
31704	:douta	=	16'h	42af;
31705	:douta	=	16'h	42d0;
31706	:douta	=	16'h	4b0f;
31707	:douta	=	16'h	73f4;
31708	:douta	=	16'h	3a8e;
31709	:douta	=	16'h	3aaf;
31710	:douta	=	16'h	4b31;
31711	:douta	=	16'h	ad34;
31712	:douta	=	16'h	6248;
31713	:douta	=	16'h	6269;
31714	:douta	=	16'h	5229;
31715	:douta	=	16'h	5249;
31716	:douta	=	16'h	5208;
31717	:douta	=	16'h	49e8;
31718	:douta	=	16'h	49c8;
31719	:douta	=	16'h	49c7;
31720	:douta	=	16'h	41a7;
31721	:douta	=	16'h	41a7;
31722	:douta	=	16'h	41a7;
31723	:douta	=	16'h	49c7;
31724	:douta	=	16'h	49e8;
31725	:douta	=	16'h	41a7;
31726	:douta	=	16'h	3986;
31727	:douta	=	16'h	39a6;
31728	:douta	=	16'h	49c7;
31729	:douta	=	16'h	41a7;
31730	:douta	=	16'h	41a7;
31731	:douta	=	16'h	4186;
31732	:douta	=	16'h	4186;
31733	:douta	=	16'h	39a6;
31734	:douta	=	16'h	41a6;
31735	:douta	=	16'h	3986;
31736	:douta	=	16'h	39a6;
31737	:douta	=	16'h	41a6;
31738	:douta	=	16'h	41a7;
31739	:douta	=	16'h	41a7;
31740	:douta	=	16'h	49e7;
31741	:douta	=	16'h	49c8;
31742	:douta	=	16'h	4187;
31743	:douta	=	16'h	49e8;
31744	:douta	=	16'h	e52a;
31745	:douta	=	16'h	6ac7;
31746	:douta	=	16'h	28e3;
31747	:douta	=	16'h	3965;
31748	:douta	=	16'h	632f;
31749	:douta	=	16'h	528b;
31750	:douta	=	16'h	3145;
31751	:douta	=	16'h	3124;
31752	:douta	=	16'h	3124;
31753	:douta	=	16'h	422a;
31754	:douta	=	16'h	3a6c;
31755	:douta	=	16'h	2168;
31756	:douta	=	16'h	2168;
31757	:douta	=	16'h	31ca;
31758	:douta	=	16'h	528b;
31759	:douta	=	16'h	422a;
31760	:douta	=	16'h	4a0a;
31761	:douta	=	16'h	526b;
31762	:douta	=	16'h	4209;
31763	:douta	=	16'h	528b;
31764	:douta	=	16'h	52cc;
31765	:douta	=	16'h	528c;
31766	:douta	=	16'h	426b;
31767	:douta	=	16'h	52ce;
31768	:douta	=	16'h	5b0e;
31769	:douta	=	16'h	634f;
31770	:douta	=	16'h	634f;
31771	:douta	=	16'h	6390;
31772	:douta	=	16'h	6b90;
31773	:douta	=	16'h	6bb0;
31774	:douta	=	16'h	6bd0;
31775	:douta	=	16'h	73f1;
31776	:douta	=	16'h	73f1;
31777	:douta	=	16'h	6bf1;
31778	:douta	=	16'h	7411;
31779	:douta	=	16'h	6bd0;
31780	:douta	=	16'h	6baf;
31781	:douta	=	16'h	638f;
31782	:douta	=	16'h	6bcf;
31783	:douta	=	16'h	638f;
31784	:douta	=	16'h	63af;
31785	:douta	=	16'h	6bd0;
31786	:douta	=	16'h	6bcf;
31787	:douta	=	16'h	636e;
31788	:douta	=	16'h	5b0d;
31789	:douta	=	16'h	4aab;
31790	:douta	=	16'h	3a6b;
31791	:douta	=	16'h	426b;
31792	:douta	=	16'h	ddb2;
31793	:douta	=	16'h	ac90;
31794	:douta	=	16'h	ac90;
31795	:douta	=	16'h	93ef;
31796	:douta	=	16'h	7b6e;
31797	:douta	=	16'h	6b0d;
31798	:douta	=	16'h	734e;
31799	:douta	=	16'h	6b0d;
31800	:douta	=	16'h	5aab;
31801	:douta	=	16'h	6b0d;
31802	:douta	=	16'h	3987;
31803	:douta	=	16'h	cd0e;
31804	:douta	=	16'h	c50c;
31805	:douta	=	16'h	ee96;
31806	:douta	=	16'h	de13;
31807	:douta	=	16'h	eeb6;
31808	:douta	=	16'h	eed7;
31809	:douta	=	16'h	eeb7;
31810	:douta	=	16'h	eeb7;
31811	:douta	=	16'h	ee96;
31812	:douta	=	16'h	e655;
31813	:douta	=	16'h	de15;
31814	:douta	=	16'h	d5d3;
31815	:douta	=	16'h	c552;
31816	:douta	=	16'h	b513;
31817	:douta	=	16'h	a4b4;
31818	:douta	=	16'h	8c74;
31819	:douta	=	16'h	8454;
31820	:douta	=	16'h	8413;
31821	:douta	=	16'h	8453;
31822	:douta	=	16'h	8412;
31823	:douta	=	16'h	73b0;
31824	:douta	=	16'h	6b6f;
31825	:douta	=	16'h	6b4e;
31826	:douta	=	16'h	6b4e;
31827	:douta	=	16'h	6b0d;
31828	:douta	=	16'h	62cd;
31829	:douta	=	16'h	630d;
31830	:douta	=	16'h	49a6;
31831	:douta	=	16'h	59c6;
31832	:douta	=	16'h	9348;
31833	:douta	=	16'h	d52e;
31834	:douta	=	16'h	d570;
31835	:douta	=	16'h	ee75;
31836	:douta	=	16'h	ee96;
31837	:douta	=	16'h	f6f8;
31838	:douta	=	16'h	e633;
31839	:douta	=	16'h	ee75;
31840	:douta	=	16'h	ee73;
31841	:douta	=	16'h	acaf;
31842	:douta	=	16'h	8b6b;
31843	:douta	=	16'h	ac6e;
31844	:douta	=	16'h	c511;
31845	:douta	=	16'h	a4b1;
31846	:douta	=	16'h	a491;
31847	:douta	=	16'h	9431;
31848	:douta	=	16'h	9411;
31849	:douta	=	16'h	83f1;
31850	:douta	=	16'h	7b90;
31851	:douta	=	16'h	734e;
31852	:douta	=	16'h	732d;
31853	:douta	=	16'h	6b0d;
31854	:douta	=	16'h	6acc;
31855	:douta	=	16'h	6aec;
31856	:douta	=	16'h	732c;
31857	:douta	=	16'h	834d;
31858	:douta	=	16'h	7b4d;
31859	:douta	=	16'h	62cc;
31860	:douta	=	16'h	62aa;
31861	:douta	=	16'h	8b4c;
31862	:douta	=	16'h	d52e;
31863	:douta	=	16'h	ddd1;
31864	:douta	=	16'h	f6b6;
31865	:douta	=	16'h	eeb7;
31866	:douta	=	16'h	d5f4;
31867	:douta	=	16'h	ddf4;
31868	:douta	=	16'h	e655;
31869	:douta	=	16'h	bd12;
31870	:douta	=	16'h	cd93;
31871	:douta	=	16'h	c594;
31872	:douta	=	16'h	acd3;
31873	:douta	=	16'h	acf4;
31874	:douta	=	16'h	b535;
31875	:douta	=	16'h	ad15;
31876	:douta	=	16'h	a4f5;
31877	:douta	=	16'h	a4d5;
31878	:douta	=	16'h	9cd4;
31879	:douta	=	16'h	94b4;
31880	:douta	=	16'h	8c73;
31881	:douta	=	16'h	8432;
31882	:douta	=	16'h	7bf1;
31883	:douta	=	16'h	7bf2;
31884	:douta	=	16'h	7390;
31885	:douta	=	16'h	634f;
31886	:douta	=	16'h	634f;
31887	:douta	=	16'h	5b0e;
31888	:douta	=	16'h	5aee;
31889	:douta	=	16'h	5b0f;
31890	:douta	=	16'h	4aae;
31891	:douta	=	16'h	4a8d;
31892	:douta	=	16'h	93ee;
31893	:douta	=	16'h	d552;
31894	:douta	=	16'h	e655;
31895	:douta	=	16'h	cdb5;
31896	:douta	=	16'h	a4b3;
31897	:douta	=	16'h	7433;
31898	:douta	=	16'h	6371;
31899	:douta	=	16'h	4acf;
31900	:douta	=	16'h	5b50;
31901	:douta	=	16'h	5310;
31902	:douta	=	16'h	4ad0;
31903	:douta	=	16'h	4aef;
31904	:douta	=	16'h	428e;
31905	:douta	=	16'h	3a6d;
31906	:douta	=	16'h	3a4d;
31907	:douta	=	16'h	29aa;
31908	:douta	=	16'h	29aa;
31909	:douta	=	16'h	29aa;
31910	:douta	=	16'h	2168;
31911	:douta	=	16'h	29a9;
31912	:douta	=	16'h	1127;
31913	:douta	=	16'h	4aae;
31914	:douta	=	16'h	21aa;
31915	:douta	=	16'h	5311;
31916	:douta	=	16'h	21aa;
31917	:douta	=	16'h	2a2c;
31918	:douta	=	16'h	1967;
31919	:douta	=	16'h	29cb;
31920	:douta	=	16'h	3a4e;
31921	:douta	=	16'h	29aa;
31922	:douta	=	16'h	1989;
31923	:douta	=	16'h	21a9;
31924	:douta	=	16'h	2189;
31925	:douta	=	16'h	21ec;
31926	:douta	=	16'h	2a0b;
31927	:douta	=	16'h	218a;
31928	:douta	=	16'h	29cb;
31929	:douta	=	16'h	2168;
31930	:douta	=	16'h	29a9;
31931	:douta	=	16'h	1906;
31932	:douta	=	16'h	10e4;
31933	:douta	=	16'h	10e5;
31934	:douta	=	16'h	10e5;
31935	:douta	=	16'h	10e5;
31936	:douta	=	16'h	1905;
31937	:douta	=	16'h	10e5;
31938	:douta	=	16'h	1084;
31939	:douta	=	16'h	08a4;
31940	:douta	=	16'h	10e5;
31941	:douta	=	16'h	1926;
31942	:douta	=	16'h	1105;
31943	:douta	=	16'h	10c4;
31944	:douta	=	16'h	1906;
31945	:douta	=	16'h	10e5;
31946	:douta	=	16'h	428e;
31947	:douta	=	16'h	29eb;
31948	:douta	=	16'h	428d;
31949	:douta	=	16'h	6b91;
31950	:douta	=	16'h	5b30;
31951	:douta	=	16'h	52ef;
31952	:douta	=	16'h	5b50;
31953	:douta	=	16'h	3a4d;
31954	:douta	=	16'h	6bd2;
31955	:douta	=	16'h	6b71;
31956	:douta	=	16'h	5b30;
31957	:douta	=	16'h	7c55;
31958	:douta	=	16'h	6371;
31959	:douta	=	16'h	4b10;
31960	:douta	=	16'h	5b93;
31961	:douta	=	16'h	5b73;
31962	:douta	=	16'h	5b92;
31963	:douta	=	16'h	5351;
31964	:douta	=	16'h	5351;
31965	:douta	=	16'h	3ad0;
31966	:douta	=	16'h	6c14;
31967	:douta	=	16'h	c67b;
31968	:douta	=	16'h	b5b7;
31969	:douta	=	16'h	6229;
31970	:douta	=	16'h	5a28;
31971	:douta	=	16'h	49e8;
31972	:douta	=	16'h	5228;
31973	:douta	=	16'h	49e8;
31974	:douta	=	16'h	49c8;
31975	:douta	=	16'h	41a7;
31976	:douta	=	16'h	41a7;
31977	:douta	=	16'h	41c7;
31978	:douta	=	16'h	41c7;
31979	:douta	=	16'h	41a7;
31980	:douta	=	16'h	41c7;
31981	:douta	=	16'h	49e7;
31982	:douta	=	16'h	41a7;
31983	:douta	=	16'h	41a7;
31984	:douta	=	16'h	41a7;
31985	:douta	=	16'h	41a7;
31986	:douta	=	16'h	41a7;
31987	:douta	=	16'h	41a6;
31988	:douta	=	16'h	41a7;
31989	:douta	=	16'h	41a6;
31990	:douta	=	16'h	3986;
31991	:douta	=	16'h	41a7;
31992	:douta	=	16'h	3986;
31993	:douta	=	16'h	41c7;
31994	:douta	=	16'h	39a6;
31995	:douta	=	16'h	41a7;
31996	:douta	=	16'h	49c8;
31997	:douta	=	16'h	41a7;
31998	:douta	=	16'h	41a7;
31999	:douta	=	16'h	41a7;
32000	:douta	=	16'h	dd0b;
32001	:douta	=	16'h	b468;
32002	:douta	=	16'h	3145;
32003	:douta	=	16'h	4165;
32004	:douta	=	16'h	4a49;
32005	:douta	=	16'h	5b2e;
32006	:douta	=	16'h	3124;
32007	:douta	=	16'h	3945;
32008	:douta	=	16'h	3124;
32009	:douta	=	16'h	3167;
32010	:douta	=	16'h	29c9;
32011	:douta	=	16'h	29a8;
32012	:douta	=	16'h	2168;
32013	:douta	=	16'h	3a2b;
32014	:douta	=	16'h	422a;
32015	:douta	=	16'h	422a;
32016	:douta	=	16'h	422a;
32017	:douta	=	16'h	4a2b;
32018	:douta	=	16'h	31a7;
32019	:douta	=	16'h	4a8c;
32020	:douta	=	16'h	52ad;
32021	:douta	=	16'h	426c;
32022	:douta	=	16'h	426c;
32023	:douta	=	16'h	52cd;
32024	:douta	=	16'h	4acd;
32025	:douta	=	16'h	5b0e;
32026	:douta	=	16'h	636f;
32027	:douta	=	16'h	638f;
32028	:douta	=	16'h	73d1;
32029	:douta	=	16'h	6bb0;
32030	:douta	=	16'h	6bd0;
32031	:douta	=	16'h	6bb0;
32032	:douta	=	16'h	6bd0;
32033	:douta	=	16'h	6bd1;
32034	:douta	=	16'h	73f1;
32035	:douta	=	16'h	638f;
32036	:douta	=	16'h	638f;
32037	:douta	=	16'h	63af;
32038	:douta	=	16'h	5b6e;
32039	:douta	=	16'h	6baf;
32040	:douta	=	16'h	73d0;
32041	:douta	=	16'h	6bf0;
32042	:douta	=	16'h	6bcf;
32043	:douta	=	16'h	6bd0;
32044	:douta	=	16'h	638f;
32045	:douta	=	16'h	6baf;
32046	:douta	=	16'h	638e;
32047	:douta	=	16'h	5b4e;
32048	:douta	=	16'h	328b;
32049	:douta	=	16'h	9430;
32050	:douta	=	16'h	b4d1;
32051	:douta	=	16'h	940f;
32052	:douta	=	16'h	732d;
32053	:douta	=	16'h	7b6e;
32054	:douta	=	16'h	6b2d;
32055	:douta	=	16'h	6b0e;
32056	:douta	=	16'h	5acd;
32057	:douta	=	16'h	3168;
32058	:douta	=	16'h	edd0;
32059	:douta	=	16'h	de12;
32060	:douta	=	16'h	ee54;
32061	:douta	=	16'h	e676;
32062	:douta	=	16'h	e654;
32063	:douta	=	16'h	eeb6;
32064	:douta	=	16'h	eeb7;
32065	:douta	=	16'h	f6f8;
32066	:douta	=	16'h	e676;
32067	:douta	=	16'h	e675;
32068	:douta	=	16'h	d5d3;
32069	:douta	=	16'h	cdb4;
32070	:douta	=	16'h	cd93;
32071	:douta	=	16'h	c573;
32072	:douta	=	16'h	b513;
32073	:douta	=	16'h	9494;
32074	:douta	=	16'h	94b5;
32075	:douta	=	16'h	8c74;
32076	:douta	=	16'h	8c54;
32077	:douta	=	16'h	8413;
32078	:douta	=	16'h	7bf2;
32079	:douta	=	16'h	6b70;
32080	:douta	=	16'h	7390;
32081	:douta	=	16'h	632e;
32082	:douta	=	16'h	630d;
32083	:douta	=	16'h	6aed;
32084	:douta	=	16'h	49e8;
32085	:douta	=	16'h	3945;
32086	:douta	=	16'h	934a;
32087	:douta	=	16'h	abe9;
32088	:douta	=	16'h	d58f;
32089	:douta	=	16'h	ddf2;
32090	:douta	=	16'h	ac2d;
32091	:douta	=	16'h	ee73;
32092	:douta	=	16'h	ee95;
32093	:douta	=	16'h	e654;
32094	:douta	=	16'h	ee95;
32095	:douta	=	16'h	b4af;
32096	:douta	=	16'h	cd31;
32097	:douta	=	16'h	b4b1;
32098	:douta	=	16'h	bd12;
32099	:douta	=	16'h	ac91;
32100	:douta	=	16'h	83cf;
32101	:douta	=	16'h	62cc;
32102	:douta	=	16'h	734f;
32103	:douta	=	16'h	8bf0;
32104	:douta	=	16'h	8c10;
32105	:douta	=	16'h	83d0;
32106	:douta	=	16'h	8bf0;
32107	:douta	=	16'h	83f0;
32108	:douta	=	16'h	7b8f;
32109	:douta	=	16'h	734d;
32110	:douta	=	16'h	62ec;
32111	:douta	=	16'h	6aec;
32112	:douta	=	16'h	62ab;
32113	:douta	=	16'h	526a;
32114	:douta	=	16'h	524a;
32115	:douta	=	16'h	b44d;
32116	:douta	=	16'h	dd91;
32117	:douta	=	16'h	e634;
32118	:douta	=	16'h	e675;
32119	:douta	=	16'h	f6f8;
32120	:douta	=	16'h	e655;
32121	:douta	=	16'h	e675;
32122	:douta	=	16'h	e655;
32123	:douta	=	16'h	de15;
32124	:douta	=	16'h	de15;
32125	:douta	=	16'h	d5b4;
32126	:douta	=	16'h	cdb4;
32127	:douta	=	16'h	ddf4;
32128	:douta	=	16'h	cdb4;
32129	:douta	=	16'h	bd34;
32130	:douta	=	16'h	9cb2;
32131	:douta	=	16'h	8c32;
32132	:douta	=	16'h	8c32;
32133	:douta	=	16'h	83f1;
32134	:douta	=	16'h	8c32;
32135	:douta	=	16'h	8411;
32136	:douta	=	16'h	8412;
32137	:douta	=	16'h	8412;
32138	:douta	=	16'h	736f;
32139	:douta	=	16'h	7370;
32140	:douta	=	16'h	738f;
32141	:douta	=	16'h	6b4f;
32142	:douta	=	16'h	7b90;
32143	:douta	=	16'h	7370;
32144	:douta	=	16'h	630e;
32145	:douta	=	16'h	836f;
32146	:douta	=	16'h	b48f;
32147	:douta	=	16'h	ddb2;
32148	:douta	=	16'h	d5d4;
32149	:douta	=	16'h	d5d4;
32150	:douta	=	16'h	bd54;
32151	:douta	=	16'h	8c95;
32152	:douta	=	16'h	8474;
32153	:douta	=	16'h	6bb1;
32154	:douta	=	16'h	6330;
32155	:douta	=	16'h	4ace;
32156	:douta	=	16'h	5b50;
32157	:douta	=	16'h	52ef;
32158	:douta	=	16'h	4aae;
32159	:douta	=	16'h	4ace;
32160	:douta	=	16'h	428d;
32161	:douta	=	16'h	322c;
32162	:douta	=	16'h	322c;
32163	:douta	=	16'h	39eb;
32164	:douta	=	16'h	31eb;
32165	:douta	=	16'h	31ca;
32166	:douta	=	16'h	1127;
32167	:douta	=	16'h	1127;
32168	:douta	=	16'h	bd34;
32169	:douta	=	16'h	8453;
32170	:douta	=	16'h	31ec;
32171	:douta	=	16'h	6bf3;
32172	:douta	=	16'h	322d;
32173	:douta	=	16'h	3a6d;
32174	:douta	=	16'h	322d;
32175	:douta	=	16'h	21eb;
32176	:douta	=	16'h	3aae;
32177	:douta	=	16'h	322c;
32178	:douta	=	16'h	21ca;
32179	:douta	=	16'h	29eb;
32180	:douta	=	16'h	324c;
32181	:douta	=	16'h	324d;
32182	:douta	=	16'h	5b30;
32183	:douta	=	16'h	1969;
32184	:douta	=	16'h	21aa;
32185	:douta	=	16'h	1927;
32186	:douta	=	16'h	1106;
32187	:douta	=	16'h	1947;
32188	:douta	=	16'h	1926;
32189	:douta	=	16'h	2168;
32190	:douta	=	16'h	1926;
32191	:douta	=	16'h	10e5;
32192	:douta	=	16'h	10e5;
32193	:douta	=	16'h	18e5;
32194	:douta	=	16'h	0883;
32195	:douta	=	16'h	18e6;
32196	:douta	=	16'h	2126;
32197	:douta	=	16'h	10e5;
32198	:douta	=	16'h	10e5;
32199	:douta	=	16'h	10c5;
32200	:douta	=	16'h	10e5;
32201	:douta	=	16'h	1906;
32202	:douta	=	16'h	6c15;
32203	:douta	=	16'h	73f3;
32204	:douta	=	16'h	7c53;
32205	:douta	=	16'h	4aef;
32206	:douta	=	16'h	5310;
32207	:douta	=	16'h	5b50;
32208	:douta	=	16'h	6371;
32209	:douta	=	16'h	7413;
32210	:douta	=	16'h	5330;
32211	:douta	=	16'h	5b91;
32212	:douta	=	16'h	5b71;
32213	:douta	=	16'h	4aef;
32214	:douta	=	16'h	5b71;
32215	:douta	=	16'h	6bd3;
32216	:douta	=	16'h	4b10;
32217	:douta	=	16'h	5352;
32218	:douta	=	16'h	5372;
32219	:douta	=	16'h	5352;
32220	:douta	=	16'h	6c34;
32221	:douta	=	16'h	4b31;
32222	:douta	=	16'h	3a8d;
32223	:douta	=	16'h	42ee;
32224	:douta	=	16'h	c69a;
32225	:douta	=	16'h	9d78;
32226	:douta	=	16'h	8474;
32227	:douta	=	16'h	6269;
32228	:douta	=	16'h	5208;
32229	:douta	=	16'h	49e8;
32230	:douta	=	16'h	41a7;
32231	:douta	=	16'h	49c8;
32232	:douta	=	16'h	41a7;
32233	:douta	=	16'h	41a7;
32234	:douta	=	16'h	41a7;
32235	:douta	=	16'h	41a7;
32236	:douta	=	16'h	49c7;
32237	:douta	=	16'h	41a6;
32238	:douta	=	16'h	41a7;
32239	:douta	=	16'h	49c7;
32240	:douta	=	16'h	41a7;
32241	:douta	=	16'h	39a6;
32242	:douta	=	16'h	41a7;
32243	:douta	=	16'h	4186;
32244	:douta	=	16'h	4186;
32245	:douta	=	16'h	41c7;
32246	:douta	=	16'h	41c7;
32247	:douta	=	16'h	3966;
32248	:douta	=	16'h	49c8;
32249	:douta	=	16'h	49c8;
32250	:douta	=	16'h	49e8;
32251	:douta	=	16'h	49e8;
32252	:douta	=	16'h	49e8;
32253	:douta	=	16'h	49e7;
32254	:douta	=	16'h	49e7;
32255	:douta	=	16'h	5209;
32256	:douta	=	16'h	dd2a;
32257	:douta	=	16'h	d52a;
32258	:douta	=	16'h	51e5;
32259	:douta	=	16'h	3945;
32260	:douta	=	16'h	41a6;
32261	:douta	=	16'h	634e;
32262	:douta	=	16'h	2904;
32263	:douta	=	16'h	2924;
32264	:douta	=	16'h	3124;
32265	:douta	=	16'h	3166;
32266	:douta	=	16'h	320a;
32267	:douta	=	16'h	2188;
32268	:douta	=	16'h	1967;
32269	:douta	=	16'h	3a2b;
32270	:douta	=	16'h	424b;
32271	:douta	=	16'h	422b;
32272	:douta	=	16'h	3a0a;
32273	:douta	=	16'h	420a;
32274	:douta	=	16'h	31a8;
32275	:douta	=	16'h	3a2a;
32276	:douta	=	16'h	4a8c;
32277	:douta	=	16'h	3a2b;
32278	:douta	=	16'h	428c;
32279	:douta	=	16'h	4acd;
32280	:douta	=	16'h	4acd;
32281	:douta	=	16'h	52ed;
32282	:douta	=	16'h	5b4f;
32283	:douta	=	16'h	6390;
32284	:douta	=	16'h	63b0;
32285	:douta	=	16'h	6bb1;
32286	:douta	=	16'h	6bb1;
32287	:douta	=	16'h	6bb0;
32288	:douta	=	16'h	6bb0;
32289	:douta	=	16'h	7411;
32290	:douta	=	16'h	73f1;
32291	:douta	=	16'h	5b6f;
32292	:douta	=	16'h	5b6e;
32293	:douta	=	16'h	638f;
32294	:douta	=	16'h	638f;
32295	:douta	=	16'h	6baf;
32296	:douta	=	16'h	6bcf;
32297	:douta	=	16'h	6bcf;
32298	:douta	=	16'h	638f;
32299	:douta	=	16'h	6bcf;
32300	:douta	=	16'h	6bd0;
32301	:douta	=	16'h	73d0;
32302	:douta	=	16'h	63af;
32303	:douta	=	16'h	5b2d;
32304	:douta	=	16'h	5b4d;
32305	:douta	=	16'h	42ec;
32306	:douta	=	16'h	6b6e;
32307	:douta	=	16'h	a470;
32308	:douta	=	16'h	9c50;
32309	:douta	=	16'h	7b8e;
32310	:douta	=	16'h	6b0d;
32311	:douta	=	16'h	62ec;
32312	:douta	=	16'h	398a;
32313	:douta	=	16'h	8b09;
32314	:douta	=	16'h	e675;
32315	:douta	=	16'h	de34;
32316	:douta	=	16'h	e696;
32317	:douta	=	16'h	e675;
32318	:douta	=	16'h	e655;
32319	:douta	=	16'h	eed7;
32320	:douta	=	16'h	e655;
32321	:douta	=	16'h	eeb7;
32322	:douta	=	16'h	de34;
32323	:douta	=	16'h	e634;
32324	:douta	=	16'h	cdb3;
32325	:douta	=	16'h	c593;
32326	:douta	=	16'h	bd54;
32327	:douta	=	16'h	bd73;
32328	:douta	=	16'h	b533;
32329	:douta	=	16'h	9494;
32330	:douta	=	16'h	8c54;
32331	:douta	=	16'h	8433;
32332	:douta	=	16'h	7c12;
32333	:douta	=	16'h	7bd1;
32334	:douta	=	16'h	738f;
32335	:douta	=	16'h	7390;
32336	:douta	=	16'h	7390;
32337	:douta	=	16'h	630e;
32338	:douta	=	16'h	632e;
32339	:douta	=	16'h	6aed;
32340	:douta	=	16'h	4146;
32341	:douta	=	16'h	6a89;
32342	:douta	=	16'h	ccee;
32343	:douta	=	16'h	dd90;
32344	:douta	=	16'h	ee95;
32345	:douta	=	16'h	ee75;
32346	:douta	=	16'h	d5d2;
32347	:douta	=	16'h	ac4e;
32348	:douta	=	16'h	f694;
32349	:douta	=	16'h	de13;
32350	:douta	=	16'h	e5f3;
32351	:douta	=	16'h	b511;
32352	:douta	=	16'h	b4b1;
32353	:douta	=	16'h	c531;
32354	:douta	=	16'h	a472;
32355	:douta	=	16'h	a492;
32356	:douta	=	16'h	9472;
32357	:douta	=	16'h	7bb0;
32358	:douta	=	16'h	736f;
32359	:douta	=	16'h	7b8f;
32360	:douta	=	16'h	9411;
32361	:douta	=	16'h	736f;
32362	:douta	=	16'h	7b90;
32363	:douta	=	16'h	83af;
32364	:douta	=	16'h	8bf0;
32365	:douta	=	16'h	8baf;
32366	:douta	=	16'h	7b4d;
32367	:douta	=	16'h	7b2d;
32368	:douta	=	16'h	6aec;
32369	:douta	=	16'h	8b6d;
32370	:douta	=	16'h	b40c;
32371	:douta	=	16'h	e632;
32372	:douta	=	16'h	d591;
32373	:douta	=	16'h	e674;
32374	:douta	=	16'h	d5b3;
32375	:douta	=	16'h	de13;
32376	:douta	=	16'h	de14;
32377	:douta	=	16'h	bd33;
32378	:douta	=	16'h	b533;
32379	:douta	=	16'h	b4f4;
32380	:douta	=	16'h	acd4;
32381	:douta	=	16'h	a4d3;
32382	:douta	=	16'h	bd74;
32383	:douta	=	16'h	bd54;
32384	:douta	=	16'h	bd54;
32385	:douta	=	16'h	b513;
32386	:douta	=	16'h	b513;
32387	:douta	=	16'h	9cb3;
32388	:douta	=	16'h	9452;
32389	:douta	=	16'h	8c32;
32390	:douta	=	16'h	8c31;
32391	:douta	=	16'h	8411;
32392	:douta	=	16'h	83f1;
32393	:douta	=	16'h	8c32;
32394	:douta	=	16'h	7bd1;
32395	:douta	=	16'h	7bb0;
32396	:douta	=	16'h	736f;
32397	:douta	=	16'h	6b4f;
32398	:douta	=	16'h	6b4f;
32399	:douta	=	16'h	528d;
32400	:douta	=	16'h	6aed;
32401	:douta	=	16'h	e614;
32402	:douta	=	16'h	d592;
32403	:douta	=	16'h	de14;
32404	:douta	=	16'h	d5b3;
32405	:douta	=	16'h	c554;
32406	:douta	=	16'h	a4d4;
32407	:douta	=	16'h	8c74;
32408	:douta	=	16'h	7c33;
32409	:douta	=	16'h	6b90;
32410	:douta	=	16'h	6370;
32411	:douta	=	16'h	52ce;
32412	:douta	=	16'h	5b0f;
32413	:douta	=	16'h	52ce;
32414	:douta	=	16'h	4aae;
32415	:douta	=	16'h	4aad;
32416	:douta	=	16'h	426c;
32417	:douta	=	16'h	320b;
32418	:douta	=	16'h	3a2c;
32419	:douta	=	16'h	39ea;
32420	:douta	=	16'h	31eb;
32421	:douta	=	16'h	21a9;
32422	:douta	=	16'h	4a4b;
32423	:douta	=	16'h	ac70;
32424	:douta	=	16'h	9494;
32425	:douta	=	16'h	5b30;
32426	:douta	=	16'h	424d;
32427	:douta	=	16'h	7414;
32428	:douta	=	16'h	42ae;
32429	:douta	=	16'h	322c;
32430	:douta	=	16'h	3a6d;
32431	:douta	=	16'h	3a4e;
32432	:douta	=	16'h	3a8e;
32433	:douta	=	16'h	324d;
32434	:douta	=	16'h	29cb;
32435	:douta	=	16'h	2a0b;
32436	:douta	=	16'h	324e;
32437	:douta	=	16'h	1989;
32438	:douta	=	16'h	7414;
32439	:douta	=	16'h	1948;
32440	:douta	=	16'h	322c;
32441	:douta	=	16'h	29cb;
32442	:douta	=	16'h	2189;
32443	:douta	=	16'h	29ca;
32444	:douta	=	16'h	1907;
32445	:douta	=	16'h	1927;
32446	:douta	=	16'h	2147;
32447	:douta	=	16'h	1968;
32448	:douta	=	16'h	10a4;
32449	:douta	=	16'h	2167;
32450	:douta	=	16'h	10a4;
32451	:douta	=	16'h	10e5;
32452	:douta	=	16'h	1906;
32453	:douta	=	16'h	10e5;
32454	:douta	=	16'h	10c5;
32455	:douta	=	16'h	10e5;
32456	:douta	=	16'h	10e5;
32457	:douta	=	16'h	10e5;
32458	:douta	=	16'h	3a4c;
32459	:douta	=	16'h	63b3;
32460	:douta	=	16'h	4aef;
32461	:douta	=	16'h	5b71;
32462	:douta	=	16'h	5b31;
32463	:douta	=	16'h	428d;
32464	:douta	=	16'h	6391;
32465	:douta	=	16'h	5b51;
32466	:douta	=	16'h	6bd2;
32467	:douta	=	16'h	8454;
32468	:douta	=	16'h	5b71;
32469	:douta	=	16'h	5331;
32470	:douta	=	16'h	5372;
32471	:douta	=	16'h	63d3;
32472	:douta	=	16'h	63b3;
32473	:douta	=	16'h	4af0;
32474	:douta	=	16'h	328e;
32475	:douta	=	16'h	4b31;
32476	:douta	=	16'h	42f0;
32477	:douta	=	16'h	21ec;
32478	:douta	=	16'h	5bb3;
32479	:douta	=	16'h	4332;
32480	:douta	=	16'h	5352;
32481	:douta	=	16'h	c639;
32482	:douta	=	16'h	ae3b;
32483	:douta	=	16'h	3189;
32484	:douta	=	16'h	628a;
32485	:douta	=	16'h	5208;
32486	:douta	=	16'h	49e7;
32487	:douta	=	16'h	41a7;
32488	:douta	=	16'h	41e7;
32489	:douta	=	16'h	49a7;
32490	:douta	=	16'h	41a7;
32491	:douta	=	16'h	49c7;
32492	:douta	=	16'h	41a7;
32493	:douta	=	16'h	49c7;
32494	:douta	=	16'h	41a7;
32495	:douta	=	16'h	41c7;
32496	:douta	=	16'h	41a7;
32497	:douta	=	16'h	3986;
32498	:douta	=	16'h	39a6;
32499	:douta	=	16'h	41a7;
32500	:douta	=	16'h	49e7;
32501	:douta	=	16'h	3986;
32502	:douta	=	16'h	39a6;
32503	:douta	=	16'h	41a7;
32504	:douta	=	16'h	49e8;
32505	:douta	=	16'h	49e8;
32506	:douta	=	16'h	49c8;
32507	:douta	=	16'h	49c8;
32508	:douta	=	16'h	49e8;
32509	:douta	=	16'h	49e8;
32510	:douta	=	16'h	49c8;
32511	:douta	=	16'h	49e8;
32512	:douta	=	16'h	dd2b;
32513	:douta	=	16'h	f5ab;
32514	:douta	=	16'h	8ba8;
32515	:douta	=	16'h	3965;
32516	:douta	=	16'h	30e3;
32517	:douta	=	16'h	630d;
32518	:douta	=	16'h	28c2;
32519	:douta	=	16'h	3124;
32520	:douta	=	16'h	3145;
32521	:douta	=	16'h	2924;
32522	:douta	=	16'h	3a2b;
32523	:douta	=	16'h	2187;
32524	:douta	=	16'h	1967;
32525	:douta	=	16'h	3a2b;
32526	:douta	=	16'h	3a2b;
32527	:douta	=	16'h	3a0a;
32528	:douta	=	16'h	31e9;
32529	:douta	=	16'h	31c9;
32530	:douta	=	16'h	31a8;
32531	:douta	=	16'h	422a;
32532	:douta	=	16'h	3a2a;
32533	:douta	=	16'h	3a4b;
32534	:douta	=	16'h	424b;
32535	:douta	=	16'h	4aac;
32536	:douta	=	16'h	52cd;
32537	:douta	=	16'h	52ed;
32538	:douta	=	16'h	636f;
32539	:douta	=	16'h	6390;
32540	:douta	=	16'h	6370;
32541	:douta	=	16'h	6370;
32542	:douta	=	16'h	636f;
32543	:douta	=	16'h	6bd0;
32544	:douta	=	16'h	6bb0;
32545	:douta	=	16'h	6bb1;
32546	:douta	=	16'h	6bf1;
32547	:douta	=	16'h	5b2e;
32548	:douta	=	16'h	636f;
32549	:douta	=	16'h	5b6e;
32550	:douta	=	16'h	636e;
32551	:douta	=	16'h	5b6e;
32552	:douta	=	16'h	5b6e;
32553	:douta	=	16'h	638f;
32554	:douta	=	16'h	638f;
32555	:douta	=	16'h	638e;
32556	:douta	=	16'h	638e;
32557	:douta	=	16'h	530d;
32558	:douta	=	16'h	5b2d;
32559	:douta	=	16'h	530c;
32560	:douta	=	16'h	530d;
32561	:douta	=	16'h	4acc;
32562	:douta	=	16'h	4acb;
32563	:douta	=	16'h	4acb;
32564	:douta	=	16'h	4acb;
32565	:douta	=	16'h	632d;
32566	:douta	=	16'h	736e;
32567	:douta	=	16'h	4a8c;
32568	:douta	=	16'h	ff37;
32569	:douta	=	16'h	de34;
32570	:douta	=	16'h	eeb6;
32571	:douta	=	16'h	eeb6;
32572	:douta	=	16'h	eeb7;
32573	:douta	=	16'h	eeb6;
32574	:douta	=	16'h	eeb6;
32575	:douta	=	16'h	eed7;
32576	:douta	=	16'h	cd93;
32577	:douta	=	16'h	d5b3;
32578	:douta	=	16'h	d5d4;
32579	:douta	=	16'h	c573;
32580	:douta	=	16'h	b4f3;
32581	:douta	=	16'h	acd4;
32582	:douta	=	16'h	b514;
32583	:douta	=	16'h	ad14;
32584	:douta	=	16'h	a4f4;
32585	:douta	=	16'h	9cb4;
32586	:douta	=	16'h	8433;
32587	:douta	=	16'h	8412;
32588	:douta	=	16'h	7bd1;
32589	:douta	=	16'h	73b0;
32590	:douta	=	16'h	6b4f;
32591	:douta	=	16'h	6b2e;
32592	:douta	=	16'h	630d;
32593	:douta	=	16'h	6b2e;
32594	:douta	=	16'h	62cd;
32595	:douta	=	16'h	72ca;
32596	:douta	=	16'h	c50d;
32597	:douta	=	16'h	c4ee;
32598	:douta	=	16'h	e633;
32599	:douta	=	16'h	ddf2;
32600	:douta	=	16'h	eeb6;
32601	:douta	=	16'h	e655;
32602	:douta	=	16'h	ddf2;
32603	:douta	=	16'h	83d0;
32604	:douta	=	16'h	5aee;
32605	:douta	=	16'h	d571;
32606	:douta	=	16'h	b490;
32607	:douta	=	16'h	9c91;
32608	:douta	=	16'h	83d1;
32609	:douta	=	16'h	73b0;
32610	:douta	=	16'h	83f2;
32611	:douta	=	16'h	83d1;
32612	:douta	=	16'h	8c11;
32613	:douta	=	16'h	83d0;
32614	:douta	=	16'h	83af;
32615	:douta	=	16'h	7b8f;
32616	:douta	=	16'h	736e;
32617	:douta	=	16'h	6b0d;
32618	:douta	=	16'h	6aec;
32619	:douta	=	16'h	62ed;
32620	:douta	=	16'h	422a;
32621	:douta	=	16'h	31a9;
32622	:douta	=	16'h	524c;
32623	:douta	=	16'h	9bec;
32624	:douta	=	16'h	c4ae;
32625	:douta	=	16'h	e5f3;
32626	:douta	=	16'h	ee96;
32627	:douta	=	16'h	f6d7;
32628	:douta	=	16'h	cd51;
32629	:douta	=	16'h	d5d2;
32630	:douta	=	16'h	de35;
32631	:douta	=	16'h	de13;
32632	:douta	=	16'h	d592;
32633	:douta	=	16'h	b514;
32634	:douta	=	16'h	8c53;
32635	:douta	=	16'h	9453;
32636	:douta	=	16'h	9c93;
32637	:douta	=	16'h	9432;
32638	:douta	=	16'h	9432;
32639	:douta	=	16'h	9452;
32640	:douta	=	16'h	8c32;
32641	:douta	=	16'h	8c31;
32642	:douta	=	16'h	8c31;
32643	:douta	=	16'h	9472;
32644	:douta	=	16'h	a4d4;
32645	:douta	=	16'h	9492;
32646	:douta	=	16'h	8c11;
32647	:douta	=	16'h	8432;
32648	:douta	=	16'h	9453;
32649	:douta	=	16'h	8412;
32650	:douta	=	16'h	7bcf;
32651	:douta	=	16'h	736e;
32652	:douta	=	16'h	6aee;
32653	:douta	=	16'h	9c0f;
32654	:douta	=	16'h	d5b3;
32655	:douta	=	16'h	eeb5;
32656	:douta	=	16'h	e655;
32657	:douta	=	16'h	ddf4;
32658	:douta	=	16'h	bd34;
32659	:douta	=	16'h	acd4;
32660	:douta	=	16'h	9494;
32661	:douta	=	16'h	9c94;
32662	:douta	=	16'h	8c53;
32663	:douta	=	16'h	8433;
32664	:douta	=	16'h	73d1;
32665	:douta	=	16'h	6b6f;
32666	:douta	=	16'h	5aee;
32667	:douta	=	16'h	630e;
32668	:douta	=	16'h	632f;
32669	:douta	=	16'h	630f;
32670	:douta	=	16'h	4a8d;
32671	:douta	=	16'h	4a8d;
32672	:douta	=	16'h	4a8d;
32673	:douta	=	16'h	424c;
32674	:douta	=	16'h	3a4c;
32675	:douta	=	16'h	29a9;
32676	:douta	=	16'h	39ea;
32677	:douta	=	16'h	b491;
32678	:douta	=	16'h	acb2;
32679	:douta	=	16'h	7bd2;
32680	:douta	=	16'h	734f;
32681	:douta	=	16'h	5b0f;
32682	:douta	=	16'h	6350;
32683	:douta	=	16'h	5b50;
32684	:douta	=	16'h	4ace;
32685	:douta	=	16'h	42ae;
32686	:douta	=	16'h	3a6c;
32687	:douta	=	16'h	3a4c;
32688	:douta	=	16'h	2a0c;
32689	:douta	=	16'h	42ae;
32690	:douta	=	16'h	2a0c;
32691	:douta	=	16'h	21cb;
32692	:douta	=	16'h	7bd1;
32693	:douta	=	16'h	a4f5;
32694	:douta	=	16'h	5331;
32695	:douta	=	16'h	3a4d;
32696	:douta	=	16'h	4aef;
32697	:douta	=	16'h	42cf;
32698	:douta	=	16'h	42ce;
32699	:douta	=	16'h	320c;
32700	:douta	=	16'h	320c;
32701	:douta	=	16'h	31eb;
32702	:douta	=	16'h	2989;
32703	:douta	=	16'h	10e5;
32704	:douta	=	16'h	320b;
32705	:douta	=	16'h	4af1;
32706	:douta	=	16'h	29ca;
32707	:douta	=	16'h	10c4;
32708	:douta	=	16'h	18e5;
32709	:douta	=	16'h	10e5;
32710	:douta	=	16'h	10c5;
32711	:douta	=	16'h	10e5;
32712	:douta	=	16'h	1906;
32713	:douta	=	16'h	1906;
32714	:douta	=	16'h	18e5;
32715	:douta	=	16'h	0884;
32716	:douta	=	16'h	5330;
32717	:douta	=	16'h	0000;
32718	:douta	=	16'h	29a9;
32719	:douta	=	16'h	6bb1;
32720	:douta	=	16'h	42ce;
32721	:douta	=	16'h	5b71;
32722	:douta	=	16'h	6bf2;
32723	:douta	=	16'h	5b72;
32724	:douta	=	16'h	5b72;
32725	:douta	=	16'h	8495;
32726	:douta	=	16'h	7c56;
32727	:douta	=	16'h	5b72;
32728	:douta	=	16'h	63b3;
32729	:douta	=	16'h	5351;
32730	:douta	=	16'h	5bb3;
32731	:douta	=	16'h	4b31;
32732	:douta	=	16'h	6bd3;
32733	:douta	=	16'h	63f4;
32734	:douta	=	16'h	6c36;
32735	:douta	=	16'h	6c56;
32736	:douta	=	16'h	53f6;
32737	:douta	=	16'h	4b73;
32738	:douta	=	16'h	94f5;
32739	:douta	=	16'h	adda;
32740	:douta	=	16'h	11cb;
32741	:douta	=	16'h	5394;
32742	:douta	=	16'h	5a27;
32743	:douta	=	16'h	5227;
32744	:douta	=	16'h	49c8;
32745	:douta	=	16'h	49e7;
32746	:douta	=	16'h	41a7;
32747	:douta	=	16'h	49c7;
32748	:douta	=	16'h	4186;
32749	:douta	=	16'h	41a6;
32750	:douta	=	16'h	41a7;
32751	:douta	=	16'h	41a7;
32752	:douta	=	16'h	41a7;
32753	:douta	=	16'h	41a7;
32754	:douta	=	16'h	39a6;
32755	:douta	=	16'h	41a7;
32756	:douta	=	16'h	41a7;
32757	:douta	=	16'h	49e7;
32758	:douta	=	16'h	49e7;
32759	:douta	=	16'h	4a08;
32760	:douta	=	16'h	49e8;
32761	:douta	=	16'h	49e8;
32762	:douta	=	16'h	49e8;
32763	:douta	=	16'h	49e8;
32764	:douta	=	16'h	49e8;
32765	:douta	=	16'h	49e8;
32766	:douta	=	16'h	49e8;
32767	:douta	=	16'h	5208;
32768	:douta	=	16'h	dd2b;
32769	:douta	=	16'h	f5ab;
32770	:douta	=	16'h	ac68;
32771	:douta	=	16'h	3944;
32772	:douta	=	16'h	30e3;
32773	:douta	=	16'h	528a;
32774	:douta	=	16'h	30e2;
32775	:douta	=	16'h	3144;
32776	:douta	=	16'h	3124;
32777	:douta	=	16'h	28e4;
32778	:douta	=	16'h	3a0a;
32779	:douta	=	16'h	1946;
32780	:douta	=	16'h	2147;
32781	:douta	=	16'h	3a2b;
32782	:douta	=	16'h	320b;
32783	:douta	=	16'h	3a0a;
32784	:douta	=	16'h	31c9;
32785	:douta	=	16'h	2987;
32786	:douta	=	16'h	31a8;
32787	:douta	=	16'h	39e9;
32788	:douta	=	16'h	3a0a;
32789	:douta	=	16'h	424b;
32790	:douta	=	16'h	426c;
32791	:douta	=	16'h	4aad;
32792	:douta	=	16'h	4aac;
32793	:douta	=	16'h	4aac;
32794	:douta	=	16'h	5b2f;
32795	:douta	=	16'h	636f;
32796	:douta	=	16'h	6370;
32797	:douta	=	16'h	6390;
32798	:douta	=	16'h	6390;
32799	:douta	=	16'h	6bb1;
32800	:douta	=	16'h	6bd1;
32801	:douta	=	16'h	63b0;
32802	:douta	=	16'h	6390;
32803	:douta	=	16'h	532e;
32804	:douta	=	16'h	532e;
32805	:douta	=	16'h	532e;
32806	:douta	=	16'h	5b2e;
32807	:douta	=	16'h	5b4e;
32808	:douta	=	16'h	532e;
32809	:douta	=	16'h	4aec;
32810	:douta	=	16'h	532d;
32811	:douta	=	16'h	5b4e;
32812	:douta	=	16'h	4aec;
32813	:douta	=	16'h	52ec;
32814	:douta	=	16'h	52ec;
32815	:douta	=	16'h	4acb;
32816	:douta	=	16'h	4acc;
32817	:douta	=	16'h	4acb;
32818	:douta	=	16'h	4acb;
32819	:douta	=	16'h	52ec;
32820	:douta	=	16'h	52ec;
32821	:douta	=	16'h	4acc;
32822	:douta	=	16'h	52ec;
32823	:douta	=	16'h	4aac;
32824	:douta	=	16'h	f696;
32825	:douta	=	16'h	f718;
32826	:douta	=	16'h	eeb7;
32827	:douta	=	16'h	eed7;
32828	:douta	=	16'h	eeb7;
32829	:douta	=	16'h	eeb7;
32830	:douta	=	16'h	eed7;
32831	:douta	=	16'h	ee96;
32832	:douta	=	16'h	c572;
32833	:douta	=	16'h	bd32;
32834	:douta	=	16'h	d5b4;
32835	:douta	=	16'h	cd73;
32836	:douta	=	16'h	ad14;
32837	:douta	=	16'h	a4b2;
32838	:douta	=	16'h	9c92;
32839	:douta	=	16'h	9cb4;
32840	:douta	=	16'h	a4f4;
32841	:douta	=	16'h	9cb4;
32842	:douta	=	16'h	9473;
32843	:douta	=	16'h	8c74;
32844	:douta	=	16'h	8411;
32845	:douta	=	16'h	7bf1;
32846	:douta	=	16'h	738f;
32847	:douta	=	16'h	734e;
32848	:douta	=	16'h	6b4e;
32849	:douta	=	16'h	62cd;
32850	:douta	=	16'h	4168;
32851	:douta	=	16'h	c4cc;
32852	:douta	=	16'h	ddf3;
32853	:douta	=	16'h	e613;
32854	:douta	=	16'h	f6d7;
32855	:douta	=	16'h	e675;
32856	:douta	=	16'h	e675;
32857	:douta	=	16'h	ee95;
32858	:douta	=	16'h	cd71;
32859	:douta	=	16'h	6b6e;
32860	:douta	=	16'h	6b70;
32861	:douta	=	16'h	cd51;
32862	:douta	=	16'h	c511;
32863	:douta	=	16'h	9452;
32864	:douta	=	16'h	9432;
32865	:douta	=	16'h	83d1;
32866	:douta	=	16'h	83f2;
32867	:douta	=	16'h	7bb0;
32868	:douta	=	16'h	83b0;
32869	:douta	=	16'h	7b6f;
32870	:douta	=	16'h	83af;
32871	:douta	=	16'h	7b8f;
32872	:douta	=	16'h	7b8f;
32873	:douta	=	16'h	734e;
32874	:douta	=	16'h	6aec;
32875	:douta	=	16'h	62ab;
32876	:douta	=	16'h	422b;
32877	:douta	=	16'h	39ea;
32878	:douta	=	16'h	ac0d;
32879	:douta	=	16'h	ddb0;
32880	:douta	=	16'h	e633;
32881	:douta	=	16'h	ddf3;
32882	:douta	=	16'h	e696;
32883	:douta	=	16'h	cd72;
32884	:douta	=	16'h	d5f4;
32885	:douta	=	16'h	cd92;
32886	:douta	=	16'h	cd52;
32887	:douta	=	16'h	c554;
32888	:douta	=	16'h	c532;
32889	:douta	=	16'h	acf3;
32890	:douta	=	16'h	a4d3;
32891	:douta	=	16'h	8433;
32892	:douta	=	16'h	7bf2;
32893	:douta	=	16'h	a4d4;
32894	:douta	=	16'h	9453;
32895	:douta	=	16'h	9451;
32896	:douta	=	16'h	9432;
32897	:douta	=	16'h	9472;
32898	:douta	=	16'h	83d0;
32899	:douta	=	16'h	9451;
32900	:douta	=	16'h	9c52;
32901	:douta	=	16'h	9452;
32902	:douta	=	16'h	9c93;
32903	:douta	=	16'h	8c30;
32904	:douta	=	16'h	8c11;
32905	:douta	=	16'h	83d0;
32906	:douta	=	16'h	6acc;
32907	:douta	=	16'h	7b6e;
32908	:douta	=	16'h	bd12;
32909	:douta	=	16'h	ee75;
32910	:douta	=	16'h	eeb6;
32911	:douta	=	16'h	d5d4;
32912	:douta	=	16'h	d5d5;
32913	:douta	=	16'h	bd74;
32914	:douta	=	16'h	bd35;
32915	:douta	=	16'h	b515;
32916	:douta	=	16'h	94b5;
32917	:douta	=	16'h	94b4;
32918	:douta	=	16'h	8432;
32919	:douta	=	16'h	7bd1;
32920	:douta	=	16'h	7390;
32921	:douta	=	16'h	632e;
32922	:douta	=	16'h	632e;
32923	:douta	=	16'h	630e;
32924	:douta	=	16'h	6b50;
32925	:douta	=	16'h	6b4f;
32926	:douta	=	16'h	4aad;
32927	:douta	=	16'h	4aad;
32928	:douta	=	16'h	4a6d;
32929	:douta	=	16'h	4a6c;
32930	:douta	=	16'h	3a0b;
32931	:douta	=	16'h	5aed;
32932	:douta	=	16'h	9c52;
32933	:douta	=	16'h	cd53;
32934	:douta	=	16'h	8c13;
32935	:douta	=	16'h	7bd2;
32936	:douta	=	16'h	736f;
32937	:douta	=	16'h	634f;
32938	:douta	=	16'h	5b2f;
32939	:douta	=	16'h	530f;
32940	:douta	=	16'h	4aad;
32941	:douta	=	16'h	428d;
32942	:douta	=	16'h	428d;
32943	:douta	=	16'h	3a2c;
32944	:douta	=	16'h	322b;
32945	:douta	=	16'h	4ace;
32946	:douta	=	16'h	21aa;
32947	:douta	=	16'h	630e;
32948	:douta	=	16'h	acd4;
32949	:douta	=	16'h	8c73;
32950	:douta	=	16'h	5351;
32951	:douta	=	16'h	4aaf;
32952	:douta	=	16'h	5310;
32953	:douta	=	16'h	4aae;
32954	:douta	=	16'h	4acf;
32955	:douta	=	16'h	324d;
32956	:douta	=	16'h	322c;
32957	:douta	=	16'h	29eb;
32958	:douta	=	16'h	2189;
32959	:douta	=	16'h	1947;
32960	:douta	=	16'h	21a9;
32961	:douta	=	16'h	3a2d;
32962	:douta	=	16'h	4af0;
32963	:douta	=	16'h	10e5;
32964	:douta	=	16'h	1083;
32965	:douta	=	16'h	10e5;
32966	:douta	=	16'h	10c5;
32967	:douta	=	16'h	10e5;
32968	:douta	=	16'h	1905;
32969	:douta	=	16'h	10e5;
32970	:douta	=	16'h	10e5;
32971	:douta	=	16'h	10c4;
32972	:douta	=	16'h	1906;
32973	:douta	=	16'h	0042;
32974	:douta	=	16'h	0884;
32975	:douta	=	16'h	8cd6;
32976	:douta	=	16'h	5b2f;
32977	:douta	=	16'h	6bd2;
32978	:douta	=	16'h	7414;
32979	:douta	=	16'h	42ce;
32980	:douta	=	16'h	7414;
32981	:douta	=	16'h	6bd3;
32982	:douta	=	16'h	73f4;
32983	:douta	=	16'h	428f;
32984	:douta	=	16'h	5b92;
32985	:douta	=	16'h	7435;
32986	:douta	=	16'h	5352;
32987	:douta	=	16'h	5bd4;
32988	:douta	=	16'h	7456;
32989	:douta	=	16'h	6c15;
32990	:douta	=	16'h	5bd5;
32991	:douta	=	16'h	6c56;
32992	:douta	=	16'h	6c57;
32993	:douta	=	16'h	3b34;
32994	:douta	=	16'h	74f9;
32995	:douta	=	16'h	c67a;
32996	:douta	=	16'h	74f9;
32997	:douta	=	16'h	43b6;
32998	:douta	=	16'h	21ea;
32999	:douta	=	16'h	41c7;
33000	:douta	=	16'h	49e7;
33001	:douta	=	16'h	41a7;
33002	:douta	=	16'h	49c7;
33003	:douta	=	16'h	49e7;
33004	:douta	=	16'h	41a7;
33005	:douta	=	16'h	3986;
33006	:douta	=	16'h	49a7;
33007	:douta	=	16'h	41c7;
33008	:douta	=	16'h	41a7;
33009	:douta	=	16'h	41a7;
33010	:douta	=	16'h	39a6;
33011	:douta	=	16'h	49e8;
33012	:douta	=	16'h	49e7;
33013	:douta	=	16'h	49e8;
33014	:douta	=	16'h	49e8;
33015	:douta	=	16'h	5229;
33016	:douta	=	16'h	49c8;
33017	:douta	=	16'h	49c8;
33018	:douta	=	16'h	49e8;
33019	:douta	=	16'h	49e8;
33020	:douta	=	16'h	49e8;
33021	:douta	=	16'h	5208;
33022	:douta	=	16'h	49e8;
33023	:douta	=	16'h	5228;
33024	:douta	=	16'h	dd4c;
33025	:douta	=	16'h	e54a;
33026	:douta	=	16'h	edab;
33027	:douta	=	16'h	28c4;
33028	:douta	=	16'h	3924;
33029	:douta	=	16'h	3945;
33030	:douta	=	16'h	49e7;
33031	:douta	=	16'h	3103;
33032	:douta	=	16'h	3124;
33033	:douta	=	16'h	3124;
33034	:douta	=	16'h	2946;
33035	:douta	=	16'h	2147;
33036	:douta	=	16'h	2147;
33037	:douta	=	16'h	1926;
33038	:douta	=	16'h	3a2b;
33039	:douta	=	16'h	31c9;
33040	:douta	=	16'h	2988;
33041	:douta	=	16'h	31a8;
33042	:douta	=	16'h	2987;
33043	:douta	=	16'h	2987;
33044	:douta	=	16'h	2987;
33045	:douta	=	16'h	3a2a;
33046	:douta	=	16'h	3a6b;
33047	:douta	=	16'h	4a8c;
33048	:douta	=	16'h	4a8c;
33049	:douta	=	16'h	4a8c;
33050	:douta	=	16'h	4acd;
33051	:douta	=	16'h	530e;
33052	:douta	=	16'h	636f;
33053	:douta	=	16'h	6390;
33054	:douta	=	16'h	6390;
33055	:douta	=	16'h	6bb1;
33056	:douta	=	16'h	6390;
33057	:douta	=	16'h	6bd1;
33058	:douta	=	16'h	6bf1;
33059	:douta	=	16'h	5b4e;
33060	:douta	=	16'h	5b6f;
33061	:douta	=	16'h	5b6f;
33062	:douta	=	16'h	532e;
33063	:douta	=	16'h	5b6e;
33064	:douta	=	16'h	5b6e;
33065	:douta	=	16'h	5b4e;
33066	:douta	=	16'h	5b4e;
33067	:douta	=	16'h	5b4e;
33068	:douta	=	16'h	52ec;
33069	:douta	=	16'h	4acb;
33070	:douta	=	16'h	4aab;
33071	:douta	=	16'h	4acc;
33072	:douta	=	16'h	4aab;
33073	:douta	=	16'h	532d;
33074	:douta	=	16'h	532d;
33075	:douta	=	16'h	530d;
33076	:douta	=	16'h	532d;
33077	:douta	=	16'h	52ec;
33078	:douta	=	16'h	530c;
33079	:douta	=	16'h	5b2e;
33080	:douta	=	16'h	42cc;
33081	:douta	=	16'h	734c;
33082	:douta	=	16'h	ff38;
33083	:douta	=	16'h	eeb7;
33084	:douta	=	16'h	eeb7;
33085	:douta	=	16'h	e696;
33086	:douta	=	16'h	eed7;
33087	:douta	=	16'h	e655;
33088	:douta	=	16'h	cd93;
33089	:douta	=	16'h	bd12;
33090	:douta	=	16'h	b513;
33091	:douta	=	16'h	c554;
33092	:douta	=	16'h	bd54;
33093	:douta	=	16'h	b535;
33094	:douta	=	16'h	b536;
33095	:douta	=	16'h	9cb4;
33096	:douta	=	16'h	8c72;
33097	:douta	=	16'h	8412;
33098	:douta	=	16'h	7bd1;
33099	:douta	=	16'h	738f;
33100	:douta	=	16'h	83f1;
33101	:douta	=	16'h	83f2;
33102	:douta	=	16'h	7bb0;
33103	:douta	=	16'h	6b4e;
33104	:douta	=	16'h	49e8;
33105	:douta	=	16'h	9b2a;
33106	:douta	=	16'h	d570;
33107	:douta	=	16'h	ddf3;
33108	:douta	=	16'h	e6b5;
33109	:douta	=	16'h	ee96;
33110	:douta	=	16'h	e654;
33111	:douta	=	16'h	ee95;
33112	:douta	=	16'h	e634;
33113	:douta	=	16'h	e655;
33114	:douta	=	16'h	ddf3;
33115	:douta	=	16'h	a492;
33116	:douta	=	16'h	7c52;
33117	:douta	=	16'h	426d;
33118	:douta	=	16'h	62eb;
33119	:douta	=	16'h	a4b3;
33120	:douta	=	16'h	7bb0;
33121	:douta	=	16'h	7bb0;
33122	:douta	=	16'h	736f;
33123	:douta	=	16'h	734e;
33124	:douta	=	16'h	6b0d;
33125	:douta	=	16'h	7b8f;
33126	:douta	=	16'h	736e;
33127	:douta	=	16'h	732c;
33128	:douta	=	16'h	730c;
33129	:douta	=	16'h	6acc;
33130	:douta	=	16'h	6aec;
33131	:douta	=	16'h	5a8c;
33132	:douta	=	16'h	a3eb;
33133	:douta	=	16'h	d50e;
33134	:douta	=	16'h	ddf4;
33135	:douta	=	16'h	eed7;
33136	:douta	=	16'h	ee96;
33137	:douta	=	16'h	eeb7;
33138	:douta	=	16'h	ee76;
33139	:douta	=	16'h	b533;
33140	:douta	=	16'h	b513;
33141	:douta	=	16'h	cd93;
33142	:douta	=	16'h	bd33;
33143	:douta	=	16'h	b513;
33144	:douta	=	16'h	9c93;
33145	:douta	=	16'h	9452;
33146	:douta	=	16'h	9452;
33147	:douta	=	16'h	8432;
33148	:douta	=	16'h	83f1;
33149	:douta	=	16'h	52ef;
33150	:douta	=	16'h	5b50;
33151	:douta	=	16'h	6b6f;
33152	:douta	=	16'h	8bf0;
33153	:douta	=	16'h	8c30;
33154	:douta	=	16'h	83cf;
33155	:douta	=	16'h	83af;
33156	:douta	=	16'h	8bae;
33157	:douta	=	16'h	8c10;
33158	:douta	=	16'h	7b8e;
33159	:douta	=	16'h	836e;
33160	:douta	=	16'h	836d;
33161	:douta	=	16'h	c552;
33162	:douta	=	16'h	ee75;
33163	:douta	=	16'h	d5b3;
33164	:douta	=	16'h	c573;
33165	:douta	=	16'h	acd3;
33166	:douta	=	16'h	a493;
33167	:douta	=	16'h	acd4;
33168	:douta	=	16'h	a4d4;
33169	:douta	=	16'h	ad15;
33170	:douta	=	16'h	94b4;
33171	:douta	=	16'h	8433;
33172	:douta	=	16'h	7bd1;
33173	:douta	=	16'h	7bd1;
33174	:douta	=	16'h	7bd1;
33175	:douta	=	16'h	7bb0;
33176	:douta	=	16'h	736f;
33177	:douta	=	16'h	6b0e;
33178	:douta	=	16'h	62ed;
33179	:douta	=	16'h	630e;
33180	:douta	=	16'h	62cd;
33181	:douta	=	16'h	630e;
33182	:douta	=	16'h	52cd;
33183	:douta	=	16'h	52ad;
33184	:douta	=	16'h	4a4c;
33185	:douta	=	16'h	9451;
33186	:douta	=	16'h	c554;
33187	:douta	=	16'h	acd3;
33188	:douta	=	16'h	9473;
33189	:douta	=	16'h	8412;
33190	:douta	=	16'h	7370;
33191	:douta	=	16'h	6b6f;
33192	:douta	=	16'h	6b4f;
33193	:douta	=	16'h	630e;
33194	:douta	=	16'h	5b0e;
33195	:douta	=	16'h	52cd;
33196	:douta	=	16'h	52ce;
33197	:douta	=	16'h	424c;
33198	:douta	=	16'h	428d;
33199	:douta	=	16'h	324c;
33200	:douta	=	16'h	324b;
33201	:douta	=	16'h	52ae;
33202	:douta	=	16'h	a4d5;
33203	:douta	=	16'h	9453;
33204	:douta	=	16'h	8413;
33205	:douta	=	16'h	7bf3;
33206	:douta	=	16'h	5b0f;
33207	:douta	=	16'h	530f;
33208	:douta	=	16'h	52ef;
33209	:douta	=	16'h	42ae;
33210	:douta	=	16'h	4aae;
33211	:douta	=	16'h	426d;
33212	:douta	=	16'h	320b;
33213	:douta	=	16'h	29ca;
33214	:douta	=	16'h	29ca;
33215	:douta	=	16'h	2168;
33216	:douta	=	16'h	31ea;
33217	:douta	=	16'h	320b;
33218	:douta	=	16'h	29a9;
33219	:douta	=	16'h	29ca;
33220	:douta	=	16'h	322b;
33221	:douta	=	16'h	1906;
33222	:douta	=	16'h	10e5;
33223	:douta	=	16'h	1906;
33224	:douta	=	16'h	10e5;
33225	:douta	=	16'h	10c5;
33226	:douta	=	16'h	18e5;
33227	:douta	=	16'h	10a4;
33228	:douta	=	16'h	10a4;
33229	:douta	=	16'h	1926;
33230	:douta	=	16'h	2127;
33231	:douta	=	16'h	0083;
33232	:douta	=	16'h	94d6;
33233	:douta	=	16'h	84b5;
33234	:douta	=	16'h	4b10;
33235	:douta	=	16'h	73f3;
33236	:douta	=	16'h	42d0;
33237	:douta	=	16'h	8cd6;
33238	:douta	=	16'h	5392;
33239	:douta	=	16'h	5331;
33240	:douta	=	16'h	63d4;
33241	:douta	=	16'h	63f5;
33242	:douta	=	16'h	63d4;
33243	:douta	=	16'h	63f4;
33244	:douta	=	16'h	63f4;
33245	:douta	=	16'h	4332;
33246	:douta	=	16'h	63f5;
33247	:douta	=	16'h	5bf5;
33248	:douta	=	16'h	5c15;
33249	:douta	=	16'h	7cb8;
33250	:douta	=	16'h	5bb4;
33251	:douta	=	16'h	53b4;
33252	:douta	=	16'h	5bd4;
33253	:douta	=	16'h	8518;
33254	:douta	=	16'h	8d9c;
33255	:douta	=	16'h	755b;
33256	:douta	=	16'h	2b13;
33257	:douta	=	16'h	49e8;
33258	:douta	=	16'h	4986;
33259	:douta	=	16'h	41a7;
33260	:douta	=	16'h	49e8;
33261	:douta	=	16'h	41a6;
33262	:douta	=	16'h	41a6;
33263	:douta	=	16'h	41a6;
33264	:douta	=	16'h	49c7;
33265	:douta	=	16'h	49c7;
33266	:douta	=	16'h	49e7;
33267	:douta	=	16'h	49e7;
33268	:douta	=	16'h	49e8;
33269	:douta	=	16'h	5228;
33270	:douta	=	16'h	5228;
33271	:douta	=	16'h	5208;
33272	:douta	=	16'h	5208;
33273	:douta	=	16'h	5249;
33274	:douta	=	16'h	5208;
33275	:douta	=	16'h	5208;
33276	:douta	=	16'h	5249;
33277	:douta	=	16'h	5228;
33278	:douta	=	16'h	5228;
33279	:douta	=	16'h	5228;
33280	:douta	=	16'h	dd4c;
33281	:douta	=	16'h	dd4a;
33282	:douta	=	16'h	f5ec;
33283	:douta	=	16'h	20a3;
33284	:douta	=	16'h	3965;
33285	:douta	=	16'h	30e3;
33286	:douta	=	16'h	52cb;
33287	:douta	=	16'h	30c2;
33288	:douta	=	16'h	3124;
33289	:douta	=	16'h	3104;
33290	:douta	=	16'h	3125;
33291	:douta	=	16'h	1967;
33292	:douta	=	16'h	2167;
33293	:douta	=	16'h	1946;
33294	:douta	=	16'h	29a9;
33295	:douta	=	16'h	29a9;
33296	:douta	=	16'h	2968;
33297	:douta	=	16'h	2967;
33298	:douta	=	16'h	2988;
33299	:douta	=	16'h	29a8;
33300	:douta	=	16'h	2987;
33301	:douta	=	16'h	3a4b;
33302	:douta	=	16'h	3a4b;
33303	:douta	=	16'h	426c;
33304	:douta	=	16'h	428c;
33305	:douta	=	16'h	4aac;
33306	:douta	=	16'h	4aad;
33307	:douta	=	16'h	52ee;
33308	:douta	=	16'h	5b4f;
33309	:douta	=	16'h	5b4f;
33310	:douta	=	16'h	5b4f;
33311	:douta	=	16'h	636f;
33312	:douta	=	16'h	6bd1;
33313	:douta	=	16'h	6bd1;
33314	:douta	=	16'h	6bf1;
33315	:douta	=	16'h	5b4e;
33316	:douta	=	16'h	5b4e;
33317	:douta	=	16'h	5b4e;
33318	:douta	=	16'h	636f;
33319	:douta	=	16'h	5b2e;
33320	:douta	=	16'h	5b4e;
33321	:douta	=	16'h	636f;
33322	:douta	=	16'h	5b6f;
33323	:douta	=	16'h	63af;
33324	:douta	=	16'h	532d;
33325	:douta	=	16'h	532e;
33326	:douta	=	16'h	4aab;
33327	:douta	=	16'h	428b;
33328	:douta	=	16'h	4acb;
33329	:douta	=	16'h	530c;
33330	:douta	=	16'h	5b2e;
33331	:douta	=	16'h	52ed;
33332	:douta	=	16'h	530d;
33333	:douta	=	16'h	530d;
33334	:douta	=	16'h	4acc;
33335	:douta	=	16'h	530c;
33336	:douta	=	16'h	5b6e;
33337	:douta	=	16'h	42ac;
33338	:douta	=	16'h	ddb4;
33339	:douta	=	16'h	ee76;
33340	:douta	=	16'h	ee96;
33341	:douta	=	16'h	e676;
33342	:douta	=	16'h	eeb6;
33343	:douta	=	16'h	de35;
33344	:douta	=	16'h	cdb3;
33345	:douta	=	16'h	c573;
33346	:douta	=	16'h	a4b3;
33347	:douta	=	16'h	acd3;
33348	:douta	=	16'h	bd55;
33349	:douta	=	16'h	ad15;
33350	:douta	=	16'h	a4d5;
33351	:douta	=	16'h	a515;
33352	:douta	=	16'h	a4d5;
33353	:douta	=	16'h	8c73;
33354	:douta	=	16'h	7bd1;
33355	:douta	=	16'h	738f;
33356	:douta	=	16'h	738f;
33357	:douta	=	16'h	738f;
33358	:douta	=	16'h	83f1;
33359	:douta	=	16'h	3146;
33360	:douta	=	16'h	59c5;
33361	:douta	=	16'h	dd91;
33362	:douta	=	16'h	ee75;
33363	:douta	=	16'h	ee76;
33364	:douta	=	16'h	eed7;
33365	:douta	=	16'h	e675;
33366	:douta	=	16'h	e675;
33367	:douta	=	16'h	e675;
33368	:douta	=	16'h	d5d3;
33369	:douta	=	16'h	de13;
33370	:douta	=	16'h	d593;
33371	:douta	=	16'h	a4b2;
33372	:douta	=	16'h	8c53;
33373	:douta	=	16'h	7c54;
33374	:douta	=	16'h	3aaf;
33375	:douta	=	16'h	62cc;
33376	:douta	=	16'h	8c11;
33377	:douta	=	16'h	7b8e;
33378	:douta	=	16'h	736f;
33379	:douta	=	16'h	736f;
33380	:douta	=	16'h	62ec;
33381	:douta	=	16'h	6b0d;
33382	:douta	=	16'h	6b2d;
33383	:douta	=	16'h	62cc;
33384	:douta	=	16'h	6b0d;
33385	:douta	=	16'h	732d;
33386	:douta	=	16'h	62cd;
33387	:douta	=	16'h	72eb;
33388	:douta	=	16'h	d52f;
33389	:douta	=	16'h	ddd2;
33390	:douta	=	16'h	e675;
33391	:douta	=	16'h	ee98;
33392	:douta	=	16'h	ee96;
33393	:douta	=	16'h	e656;
33394	:douta	=	16'h	de35;
33395	:douta	=	16'h	cd94;
33396	:douta	=	16'h	8452;
33397	:douta	=	16'h	a4f3;
33398	:douta	=	16'h	a4b3;
33399	:douta	=	16'h	a493;
33400	:douta	=	16'h	a4d4;
33401	:douta	=	16'h	9453;
33402	:douta	=	16'h	8c32;
33403	:douta	=	16'h	9453;
33404	:douta	=	16'h	8c72;
33405	:douta	=	16'h	6b70;
33406	:douta	=	16'h	5330;
33407	:douta	=	16'h	5330;
33408	:douta	=	16'h	5b2f;
33409	:douta	=	16'h	630f;
33410	:douta	=	16'h	736f;
33411	:douta	=	16'h	632d;
33412	:douta	=	16'h	528c;
33413	:douta	=	16'h	4a2b;
33414	:douta	=	16'h	7b6d;
33415	:douta	=	16'h	ac70;
33416	:douta	=	16'h	f6d6;
33417	:douta	=	16'h	ddf4;
33418	:douta	=	16'h	ee97;
33419	:douta	=	16'h	f6b6;
33420	:douta	=	16'h	ddf5;
33421	:douta	=	16'h	b4d4;
33422	:douta	=	16'h	9c94;
33423	:douta	=	16'h	9473;
33424	:douta	=	16'h	9454;
33425	:douta	=	16'h	9c94;
33426	:douta	=	16'h	9474;
33427	:douta	=	16'h	8c53;
33428	:douta	=	16'h	8412;
33429	:douta	=	16'h	83f1;
33430	:douta	=	16'h	7bd1;
33431	:douta	=	16'h	7b90;
33432	:douta	=	16'h	736f;
33433	:douta	=	16'h	6b2e;
33434	:douta	=	16'h	732e;
33435	:douta	=	16'h	630d;
33436	:douta	=	16'h	630e;
33437	:douta	=	16'h	52ad;
33438	:douta	=	16'h	426b;
33439	:douta	=	16'h	528c;
33440	:douta	=	16'h	9432;
33441	:douta	=	16'h	c596;
33442	:douta	=	16'h	b4f4;
33443	:douta	=	16'h	9452;
33444	:douta	=	16'h	8c32;
33445	:douta	=	16'h	8c31;
33446	:douta	=	16'h	7390;
33447	:douta	=	16'h	7390;
33448	:douta	=	16'h	630e;
33449	:douta	=	16'h	5aed;
33450	:douta	=	16'h	5aee;
33451	:douta	=	16'h	52cd;
33452	:douta	=	16'h	4aad;
33453	:douta	=	16'h	428d;
33454	:douta	=	16'h	428d;
33455	:douta	=	16'h	320b;
33456	:douta	=	16'h	3a2b;
33457	:douta	=	16'h	9c94;
33458	:douta	=	16'h	8433;
33459	:douta	=	16'h	7c12;
33460	:douta	=	16'h	7bd2;
33461	:douta	=	16'h	7bf2;
33462	:douta	=	16'h	5b0f;
33463	:douta	=	16'h	4ace;
33464	:douta	=	16'h	42ce;
33465	:douta	=	16'h	428e;
33466	:douta	=	16'h	428e;
33467	:douta	=	16'h	3a6d;
33468	:douta	=	16'h	322c;
33469	:douta	=	16'h	320b;
33470	:douta	=	16'h	29a9;
33471	:douta	=	16'h	2188;
33472	:douta	=	16'h	42ae;
33473	:douta	=	16'h	5b30;
33474	:douta	=	16'h	426d;
33475	:douta	=	16'h	29eb;
33476	:douta	=	16'h	29ca;
33477	:douta	=	16'h	29ca;
33478	:douta	=	16'h	10e5;
33479	:douta	=	16'h	10e5;
33480	:douta	=	16'h	10c4;
33481	:douta	=	16'h	10c4;
33482	:douta	=	16'h	10e5;
33483	:douta	=	16'h	10c4;
33484	:douta	=	16'h	10c4;
33485	:douta	=	16'h	10e5;
33486	:douta	=	16'h	1906;
33487	:douta	=	16'h	10e6;
33488	:douta	=	16'h	4acd;
33489	:douta	=	16'h	6370;
33490	:douta	=	16'h	7414;
33491	:douta	=	16'h	7c75;
33492	:douta	=	16'h	5b71;
33493	:douta	=	16'h	5b72;
33494	:douta	=	16'h	5351;
33495	:douta	=	16'h	84d8;
33496	:douta	=	16'h	7456;
33497	:douta	=	16'h	6436;
33498	:douta	=	16'h	5bb4;
33499	:douta	=	16'h	63f5;
33500	:douta	=	16'h	6c15;
33501	:douta	=	16'h	84b8;
33502	:douta	=	16'h	5bd5;
33503	:douta	=	16'h	6c77;
33504	:douta	=	16'h	7cd9;
33505	:douta	=	16'h	5bd4;
33506	:douta	=	16'h	6416;
33507	:douta	=	16'h	53d4;
33508	:douta	=	16'h	6c57;
33509	:douta	=	16'h	6c77;
33510	:douta	=	16'h	9579;
33511	:douta	=	16'h	7d39;
33512	:douta	=	16'h	8d9b;
33513	:douta	=	16'h	4bb5;
33514	:douta	=	16'h	422a;
33515	:douta	=	16'h	4165;
33516	:douta	=	16'h	41a6;
33517	:douta	=	16'h	49c7;
33518	:douta	=	16'h	41a6;
33519	:douta	=	16'h	49a7;
33520	:douta	=	16'h	41a7;
33521	:douta	=	16'h	49e7;
33522	:douta	=	16'h	49e7;
33523	:douta	=	16'h	5208;
33524	:douta	=	16'h	5208;
33525	:douta	=	16'h	49e8;
33526	:douta	=	16'h	5208;
33527	:douta	=	16'h	5229;
33528	:douta	=	16'h	5208;
33529	:douta	=	16'h	5229;
33530	:douta	=	16'h	5228;
33531	:douta	=	16'h	5249;
33532	:douta	=	16'h	4a08;
33533	:douta	=	16'h	49e8;
33534	:douta	=	16'h	5229;
33535	:douta	=	16'h	5229;
33536	:douta	=	16'h	dd4b;
33537	:douta	=	16'h	dd2b;
33538	:douta	=	16'h	ed8b;
33539	:douta	=	16'h	41c5;
33540	:douta	=	16'h	3945;
33541	:douta	=	16'h	30e3;
33542	:douta	=	16'h	6b90;
33543	:douta	=	16'h	3124;
33544	:douta	=	16'h	3124;
33545	:douta	=	16'h	3924;
33546	:douta	=	16'h	2904;
33547	:douta	=	16'h	2168;
33548	:douta	=	16'h	1926;
33549	:douta	=	16'h	1926;
33550	:douta	=	16'h	29a9;
33551	:douta	=	16'h	29a9;
33552	:douta	=	16'h	29c9;
33553	:douta	=	16'h	2988;
33554	:douta	=	16'h	2968;
33555	:douta	=	16'h	320b;
33556	:douta	=	16'h	3a4c;
33557	:douta	=	16'h	3a2b;
33558	:douta	=	16'h	3a4c;
33559	:douta	=	16'h	3a4b;
33560	:douta	=	16'h	426c;
33561	:douta	=	16'h	4aad;
33562	:douta	=	16'h	52ee;
33563	:douta	=	16'h	5b2f;
33564	:douta	=	16'h	530e;
33565	:douta	=	16'h	5b4f;
33566	:douta	=	16'h	530e;
33567	:douta	=	16'h	4aed;
33568	:douta	=	16'h	530e;
33569	:douta	=	16'h	5b4f;
33570	:douta	=	16'h	5b4f;
33571	:douta	=	16'h	532e;
33572	:douta	=	16'h	5b4e;
33573	:douta	=	16'h	5b4e;
33574	:douta	=	16'h	534e;
33575	:douta	=	16'h	5b4e;
33576	:douta	=	16'h	5b4e;
33577	:douta	=	16'h	5b6f;
33578	:douta	=	16'h	5b6f;
33579	:douta	=	16'h	638f;
33580	:douta	=	16'h	5b6f;
33581	:douta	=	16'h	5b6e;
33582	:douta	=	16'h	530d;
33583	:douta	=	16'h	4acc;
33584	:douta	=	16'h	4acc;
33585	:douta	=	16'h	530d;
33586	:douta	=	16'h	4acc;
33587	:douta	=	16'h	530d;
33588	:douta	=	16'h	428b;
33589	:douta	=	16'h	4aac;
33590	:douta	=	16'h	52ec;
33591	:douta	=	16'h	530c;
33592	:douta	=	16'h	530d;
33593	:douta	=	16'h	532d;
33594	:douta	=	16'h	530c;
33595	:douta	=	16'h	acb1;
33596	:douta	=	16'h	e614;
33597	:douta	=	16'h	d5f5;
33598	:douta	=	16'h	de35;
33599	:douta	=	16'h	d5f4;
33600	:douta	=	16'h	c5b4;
33601	:douta	=	16'h	bd53;
33602	:douta	=	16'h	b514;
33603	:douta	=	16'h	a4d4;
33604	:douta	=	16'h	9cb5;
33605	:douta	=	16'h	a4f5;
33606	:douta	=	16'h	a515;
33607	:douta	=	16'h	9cd4;
33608	:douta	=	16'h	94b4;
33609	:douta	=	16'h	8411;
33610	:douta	=	16'h	738e;
33611	:douta	=	16'h	734e;
33612	:douta	=	16'h	734e;
33613	:douta	=	16'h	6b2e;
33614	:douta	=	16'h	49a5;
33615	:douta	=	16'h	e5d1;
33616	:douta	=	16'h	cd0d;
33617	:douta	=	16'h	eeb5;
33618	:douta	=	16'h	e613;
33619	:douta	=	16'h	eed7;
33620	:douta	=	16'h	eeb7;
33621	:douta	=	16'h	eeb7;
33622	:douta	=	16'h	de34;
33623	:douta	=	16'h	e635;
33624	:douta	=	16'h	cd73;
33625	:douta	=	16'h	cd73;
33626	:douta	=	16'h	bd52;
33627	:douta	=	16'h	9cb3;
33628	:douta	=	16'h	8c73;
33629	:douta	=	16'h	8453;
33630	:douta	=	16'h	8473;
33631	:douta	=	16'h	6bd3;
33632	:douta	=	16'h	31ea;
33633	:douta	=	16'h	5acd;
33634	:douta	=	16'h	732d;
33635	:douta	=	16'h	6b0d;
33636	:douta	=	16'h	6b0d;
33637	:douta	=	16'h	6acc;
33638	:douta	=	16'h	62cc;
33639	:douta	=	16'h	5a8b;
33640	:douta	=	16'h	4a2a;
33641	:douta	=	16'h	72ea;
33642	:douta	=	16'h	d52e;
33643	:douta	=	16'h	e612;
33644	:douta	=	16'h	eeb6;
33645	:douta	=	16'h	f6f8;
33646	:douta	=	16'h	ac70;
33647	:douta	=	16'h	ee96;
33648	:douta	=	16'h	de54;
33649	:douta	=	16'h	cdb4;
33650	:douta	=	16'h	bd54;
33651	:douta	=	16'h	b514;
33652	:douta	=	16'h	b515;
33653	:douta	=	16'h	8c94;
33654	:douta	=	16'h	9473;
33655	:douta	=	16'h	acd4;
33656	:douta	=	16'h	a4b4;
33657	:douta	=	16'h	9452;
33658	:douta	=	16'h	8411;
33659	:douta	=	16'h	8412;
33660	:douta	=	16'h	8c12;
33661	:douta	=	16'h	83f1;
33662	:douta	=	16'h	7b8f;
33663	:douta	=	16'h	7baf;
33664	:douta	=	16'h	734e;
33665	:douta	=	16'h	734e;
33666	:douta	=	16'h	62ed;
33667	:douta	=	16'h	93ee;
33668	:douta	=	16'h	b4b1;
33669	:douta	=	16'h	e613;
33670	:douta	=	16'h	b4d3;
33671	:douta	=	16'h	c553;
33672	:douta	=	16'h	d5f4;
33673	:douta	=	16'h	c553;
33674	:douta	=	16'h	acd3;
33675	:douta	=	16'h	9c53;
33676	:douta	=	16'h	9453;
33677	:douta	=	16'h	9452;
33678	:douta	=	16'h	9c93;
33679	:douta	=	16'h	a4d4;
33680	:douta	=	16'h	a4b4;
33681	:douta	=	16'h	8c53;
33682	:douta	=	16'h	8432;
33683	:douta	=	16'h	8432;
33684	:douta	=	16'h	83f1;
33685	:douta	=	16'h	736e;
33686	:douta	=	16'h	7bb0;
33687	:douta	=	16'h	734e;
33688	:douta	=	16'h	6b0d;
33689	:douta	=	16'h	6b2e;
33690	:douta	=	16'h	6b0e;
33691	:douta	=	16'h	62ac;
33692	:douta	=	16'h	6aed;
33693	:douta	=	16'h	83d0;
33694	:douta	=	16'h	a4b4;
33695	:douta	=	16'h	a493;
33696	:douta	=	16'h	9cb3;
33697	:douta	=	16'h	9c94;
33698	:douta	=	16'h	9453;
33699	:douta	=	16'h	83d1;
33700	:douta	=	16'h	83d0;
33701	:douta	=	16'h	734f;
33702	:douta	=	16'h	736f;
33703	:douta	=	16'h	630e;
33704	:douta	=	16'h	630e;
33705	:douta	=	16'h	5b0d;
33706	:douta	=	16'h	5acd;
33707	:douta	=	16'h	52ad;
33708	:douta	=	16'h	4a8c;
33709	:douta	=	16'h	424c;
33710	:douta	=	16'h	630d;
33711	:douta	=	16'h	acd4;
33712	:douta	=	16'h	a4b5;
33713	:douta	=	16'h	8c73;
33714	:douta	=	16'h	8c33;
33715	:douta	=	16'h	8452;
33716	:douta	=	16'h	8413;
33717	:douta	=	16'h	7bf2;
33718	:douta	=	16'h	632f;
33719	:douta	=	16'h	4a8d;
33720	:douta	=	16'h	4a8d;
33721	:douta	=	16'h	52ce;
33722	:douta	=	16'h	4aad;
33723	:douta	=	16'h	3a4d;
33724	:douta	=	16'h	320b;
33725	:douta	=	16'h	320b;
33726	:douta	=	16'h	3a2b;
33727	:douta	=	16'h	5b72;
33728	:douta	=	16'h	6b4e;
33729	:douta	=	16'h	6bf3;
33730	:douta	=	16'h	3a4e;
33731	:douta	=	16'h	530f;
33732	:douta	=	16'h	5310;
33733	:douta	=	16'h	2189;
33734	:douta	=	16'h	2168;
33735	:douta	=	16'h	29aa;
33736	:douta	=	16'h	18e6;
33737	:douta	=	16'h	0884;
33738	:douta	=	16'h	18e5;
33739	:douta	=	16'h	08c4;
33740	:douta	=	16'h	10e5;
33741	:douta	=	16'h	18e5;
33742	:douta	=	16'h	10e5;
33743	:douta	=	16'h	10e6;
33744	:douta	=	16'h	1107;
33745	:douta	=	16'h	6371;
33746	:douta	=	16'h	6bb3;
33747	:douta	=	16'h	6bf3;
33748	:douta	=	16'h	7c75;
33749	:douta	=	16'h	6c35;
33750	:douta	=	16'h	9d59;
33751	:douta	=	16'h	7435;
33752	:douta	=	16'h	63f5;
33753	:douta	=	16'h	7456;
33754	:douta	=	16'h	63f5;
33755	:douta	=	16'h	6c56;
33756	:douta	=	16'h	7456;
33757	:douta	=	16'h	5bb4;
33758	:douta	=	16'h	5bf5;
33759	:douta	=	16'h	7497;
33760	:douta	=	16'h	5bd4;
33761	:douta	=	16'h	5394;
33762	:douta	=	16'h	6c77;
33763	:douta	=	16'h	5bd4;
33764	:douta	=	16'h	53b4;
33765	:douta	=	16'h	4b93;
33766	:douta	=	16'h	6436;
33767	:douta	=	16'h	74b8;
33768	:douta	=	16'h	53f6;
33769	:douta	=	16'h	8d7a;
33770	:douta	=	16'h	7c97;
33771	:douta	=	16'h	959c;
33772	:douta	=	16'h	73f3;
33773	:douta	=	16'h	3924;
33774	:douta	=	16'h	49e7;
33775	:douta	=	16'h	49e7;
33776	:douta	=	16'h	49e7;
33777	:douta	=	16'h	49e8;
33778	:douta	=	16'h	5228;
33779	:douta	=	16'h	5208;
33780	:douta	=	16'h	5229;
33781	:douta	=	16'h	5249;
33782	:douta	=	16'h	5228;
33783	:douta	=	16'h	5208;
33784	:douta	=	16'h	5228;
33785	:douta	=	16'h	5208;
33786	:douta	=	16'h	5208;
33787	:douta	=	16'h	5208;
33788	:douta	=	16'h	5208;
33789	:douta	=	16'h	5228;
33790	:douta	=	16'h	5208;
33791	:douta	=	16'h	5228;
33792	:douta	=	16'h	dd4c;
33793	:douta	=	16'h	dd4b;
33794	:douta	=	16'h	e54b;
33795	:douta	=	16'h	6265;
33796	:douta	=	16'h	3965;
33797	:douta	=	16'h	3924;
33798	:douta	=	16'h	6b6f;
33799	:douta	=	16'h	41a6;
33800	:douta	=	16'h	3944;
33801	:douta	=	16'h	3144;
33802	:douta	=	16'h	2904;
33803	:douta	=	16'h	2988;
33804	:douta	=	16'h	1946;
33805	:douta	=	16'h	29a9;
33806	:douta	=	16'h	29a9;
33807	:douta	=	16'h	2168;
33808	:douta	=	16'h	2988;
33809	:douta	=	16'h	2988;
33810	:douta	=	16'h	2988;
33811	:douta	=	16'h	3a2c;
33812	:douta	=	16'h	3a6c;
33813	:douta	=	16'h	3a2b;
33814	:douta	=	16'h	3a4c;
33815	:douta	=	16'h	322b;
33816	:douta	=	16'h	3a2b;
33817	:douta	=	16'h	426c;
33818	:douta	=	16'h	530e;
33819	:douta	=	16'h	532e;
33820	:douta	=	16'h	530e;
33821	:douta	=	16'h	530e;
33822	:douta	=	16'h	530e;
33823	:douta	=	16'h	4aed;
33824	:douta	=	16'h	532e;
33825	:douta	=	16'h	5b4f;
33826	:douta	=	16'h	638f;
33827	:douta	=	16'h	530e;
33828	:douta	=	16'h	532d;
33829	:douta	=	16'h	534e;
33830	:douta	=	16'h	534e;
33831	:douta	=	16'h	534e;
33832	:douta	=	16'h	5b4e;
33833	:douta	=	16'h	5b4e;
33834	:douta	=	16'h	5b6f;
33835	:douta	=	16'h	638f;
33836	:douta	=	16'h	5b6e;
33837	:douta	=	16'h	534e;
33838	:douta	=	16'h	5b4e;
33839	:douta	=	16'h	5b2d;
33840	:douta	=	16'h	4acc;
33841	:douta	=	16'h	532d;
33842	:douta	=	16'h	530d;
33843	:douta	=	16'h	52ec;
33844	:douta	=	16'h	52ec;
33845	:douta	=	16'h	4acc;
33846	:douta	=	16'h	4aab;
33847	:douta	=	16'h	4acc;
33848	:douta	=	16'h	4acb;
33849	:douta	=	16'h	4acb;
33850	:douta	=	16'h	5b4d;
33851	:douta	=	16'h	4aed;
33852	:douta	=	16'h	7b8f;
33853	:douta	=	16'h	ddb3;
33854	:douta	=	16'h	ddf4;
33855	:douta	=	16'h	cdb3;
33856	:douta	=	16'h	b533;
33857	:douta	=	16'h	bd53;
33858	:douta	=	16'h	b535;
33859	:douta	=	16'h	acf4;
33860	:douta	=	16'h	a4d4;
33861	:douta	=	16'h	8c74;
33862	:douta	=	16'h	9453;
33863	:douta	=	16'h	9493;
33864	:douta	=	16'h	8c53;
33865	:douta	=	16'h	7bf1;
33866	:douta	=	16'h	736e;
33867	:douta	=	16'h	736e;
33868	:douta	=	16'h	62cc;
33869	:douta	=	16'h	5209;
33870	:douta	=	16'h	8ae7;
33871	:douta	=	16'h	ee73;
33872	:douta	=	16'h	c50e;
33873	:douta	=	16'h	e653;
33874	:douta	=	16'h	ddb1;
33875	:douta	=	16'h	eeb7;
33876	:douta	=	16'h	e676;
33877	:douta	=	16'h	e676;
33878	:douta	=	16'h	de35;
33879	:douta	=	16'h	d5f3;
33880	:douta	=	16'h	bd13;
33881	:douta	=	16'h	bd33;
33882	:douta	=	16'h	acd3;
33883	:douta	=	16'h	9473;
33884	:douta	=	16'h	8c53;
33885	:douta	=	16'h	8412;
33886	:douta	=	16'h	8412;
33887	:douta	=	16'h	5b2e;
33888	:douta	=	16'h	424c;
33889	:douta	=	16'h	29ca;
33890	:douta	=	16'h	7b4e;
33891	:douta	=	16'h	7b6e;
33892	:douta	=	16'h	6b2c;
33893	:douta	=	16'h	6b0c;
33894	:douta	=	16'h	6aec;
33895	:douta	=	16'h	524b;
33896	:douta	=	16'h	628b;
33897	:douta	=	16'h	bcad;
33898	:douta	=	16'h	e614;
33899	:douta	=	16'h	eeb6;
33900	:douta	=	16'h	de55;
33901	:douta	=	16'h	e675;
33902	:douta	=	16'h	a4b3;
33903	:douta	=	16'h	de14;
33904	:douta	=	16'h	cd54;
33905	:douta	=	16'h	b534;
33906	:douta	=	16'h	ad14;
33907	:douta	=	16'h	acf4;
33908	:douta	=	16'h	ad15;
33909	:douta	=	16'h	9cf5;
33910	:douta	=	16'h	7bf1;
33911	:douta	=	16'h	8c33;
33912	:douta	=	16'h	9c93;
33913	:douta	=	16'h	8c32;
33914	:douta	=	16'h	83d1;
33915	:douta	=	16'h	83d0;
33916	:douta	=	16'h	83f1;
33917	:douta	=	16'h	83d0;
33918	:douta	=	16'h	736e;
33919	:douta	=	16'h	7b8f;
33920	:douta	=	16'h	736e;
33921	:douta	=	16'h	62cc;
33922	:douta	=	16'h	7b4d;
33923	:douta	=	16'h	f696;
33924	:douta	=	16'h	ee96;
33925	:douta	=	16'h	bd33;
33926	:douta	=	16'h	9434;
33927	:douta	=	16'h	cd74;
33928	:douta	=	16'h	de15;
33929	:douta	=	16'h	d5d4;
33930	:douta	=	16'h	bd55;
33931	:douta	=	16'h	b535;
33932	:douta	=	16'h	9452;
33933	:douta	=	16'h	8410;
33934	:douta	=	16'h	8c11;
33935	:douta	=	16'h	8c11;
33936	:douta	=	16'h	8c11;
33937	:douta	=	16'h	83f0;
33938	:douta	=	16'h	83d0;
33939	:douta	=	16'h	7b90;
33940	:douta	=	16'h	7bb0;
33941	:douta	=	16'h	734e;
33942	:douta	=	16'h	736f;
33943	:douta	=	16'h	7b6f;
33944	:douta	=	16'h	734e;
33945	:douta	=	16'h	5a8c;
33946	:douta	=	16'h	528c;
33947	:douta	=	16'h	7b8f;
33948	:douta	=	16'h	acd4;
33949	:douta	=	16'h	bd15;
33950	:douta	=	16'h	9cb3;
33951	:douta	=	16'h	9472;
33952	:douta	=	16'h	8c32;
33953	:douta	=	16'h	9453;
33954	:douta	=	16'h	8412;
33955	:douta	=	16'h	7bb0;
33956	:douta	=	16'h	7bb0;
33957	:douta	=	16'h	7b8f;
33958	:douta	=	16'h	736f;
33959	:douta	=	16'h	6b2e;
33960	:douta	=	16'h	630e;
33961	:douta	=	16'h	630d;
33962	:douta	=	16'h	52cd;
33963	:douta	=	16'h	52ad;
33964	:douta	=	16'h	528d;
33965	:douta	=	16'h	acb1;
33966	:douta	=	16'h	cd94;
33967	:douta	=	16'h	a4d3;
33968	:douta	=	16'h	9c94;
33969	:douta	=	16'h	9474;
33970	:douta	=	16'h	8433;
33971	:douta	=	16'h	7bf2;
33972	:douta	=	16'h	7390;
33973	:douta	=	16'h	6b70;
33974	:douta	=	16'h	5b2f;
33975	:douta	=	16'h	52ce;
33976	:douta	=	16'h	4ace;
33977	:douta	=	16'h	4a8d;
33978	:douta	=	16'h	426d;
33979	:douta	=	16'h	428d;
33980	:douta	=	16'h	428d;
33981	:douta	=	16'h	3a2c;
33982	:douta	=	16'h	322d;
33983	:douta	=	16'h	426d;
33984	:douta	=	16'h	c5b7;
33985	:douta	=	16'h	4b30;
33986	:douta	=	16'h	428e;
33987	:douta	=	16'h	6bb1;
33988	:douta	=	16'h	5b30;
33989	:douta	=	16'h	29a9;
33990	:douta	=	16'h	29a9;
33991	:douta	=	16'h	2168;
33992	:douta	=	16'h	31ca;
33993	:douta	=	16'h	29a9;
33994	:douta	=	16'h	1083;
33995	:douta	=	16'h	10e5;
33996	:douta	=	16'h	18e5;
33997	:douta	=	16'h	1905;
33998	:douta	=	16'h	1905;
33999	:douta	=	16'h	10e5;
34000	:douta	=	16'h	10e6;
34001	:douta	=	16'h	428c;
34002	:douta	=	16'h	84b6;
34003	:douta	=	16'h	7c75;
34004	:douta	=	16'h	7435;
34005	:douta	=	16'h	7c76;
34006	:douta	=	16'h	63f4;
34007	:douta	=	16'h	5bb4;
34008	:douta	=	16'h	6c35;
34009	:douta	=	16'h	5bf5;
34010	:douta	=	16'h	84b7;
34011	:douta	=	16'h	9559;
34012	:douta	=	16'h	63f4;
34013	:douta	=	16'h	7c96;
34014	:douta	=	16'h	84d8;
34015	:douta	=	16'h	4b73;
34016	:douta	=	16'h	5bd4;
34017	:douta	=	16'h	53b4;
34018	:douta	=	16'h	6415;
34019	:douta	=	16'h	5bd5;
34020	:douta	=	16'h	5394;
34021	:douta	=	16'h	4b53;
34022	:douta	=	16'h	6c56;
34023	:douta	=	16'h	6477;
34024	:douta	=	16'h	6cb9;
34025	:douta	=	16'h	4311;
34026	:douta	=	16'h	1948;
34027	:douta	=	16'h	5b70;
34028	:douta	=	16'h	6c55;
34029	:douta	=	16'h	8c32;
34030	:douta	=	16'h	49c7;
34031	:douta	=	16'h	49e8;
34032	:douta	=	16'h	5208;
34033	:douta	=	16'h	49e7;
34034	:douta	=	16'h	5208;
34035	:douta	=	16'h	5229;
34036	:douta	=	16'h	5229;
34037	:douta	=	16'h	49e8;
34038	:douta	=	16'h	4a08;
34039	:douta	=	16'h	5228;
34040	:douta	=	16'h	49e8;
34041	:douta	=	16'h	4a08;
34042	:douta	=	16'h	49e8;
34043	:douta	=	16'h	5228;
34044	:douta	=	16'h	49e8;
34045	:douta	=	16'h	49e8;
34046	:douta	=	16'h	5208;
34047	:douta	=	16'h	5208;
34048	:douta	=	16'h	dd4b;
34049	:douta	=	16'h	dd4b;
34050	:douta	=	16'h	e54b;
34051	:douta	=	16'h	ac29;
34052	:douta	=	16'h	4165;
34053	:douta	=	16'h	3945;
34054	:douta	=	16'h	632e;
34055	:douta	=	16'h	630d;
34056	:douta	=	16'h	3944;
34057	:douta	=	16'h	3924;
34058	:douta	=	16'h	3104;
34059	:douta	=	16'h	10e4;
34060	:douta	=	16'h	1083;
34061	:douta	=	16'h	10a4;
34062	:douta	=	16'h	2125;
34063	:douta	=	16'h	2125;
34064	:douta	=	16'h	1905;
34065	:douta	=	16'h	1905;
34066	:douta	=	16'h	1906;
34067	:douta	=	16'h	31eb;
34068	:douta	=	16'h	322b;
34069	:douta	=	16'h	322b;
34070	:douta	=	16'h	3a2c;
34071	:douta	=	16'h	320b;
34072	:douta	=	16'h	320a;
34073	:douta	=	16'h	3a2b;
34074	:douta	=	16'h	4aad;
34075	:douta	=	16'h	4ace;
34076	:douta	=	16'h	4aee;
34077	:douta	=	16'h	532f;
34078	:douta	=	16'h	530e;
34079	:douta	=	16'h	532f;
34080	:douta	=	16'h	532f;
34081	:douta	=	16'h	5b4f;
34082	:douta	=	16'h	5b6f;
34083	:douta	=	16'h	4acd;
34084	:douta	=	16'h	532e;
34085	:douta	=	16'h	4aed;
34086	:douta	=	16'h	4aed;
34087	:douta	=	16'h	530d;
34088	:douta	=	16'h	530d;
34089	:douta	=	16'h	4b0d;
34090	:douta	=	16'h	532e;
34091	:douta	=	16'h	534e;
34092	:douta	=	16'h	5b6e;
34093	:douta	=	16'h	5b6f;
34094	:douta	=	16'h	428b;
34095	:douta	=	16'h	4aac;
34096	:douta	=	16'h	530d;
34097	:douta	=	16'h	532d;
34098	:douta	=	16'h	5b4e;
34099	:douta	=	16'h	636f;
34100	:douta	=	16'h	5b6f;
34101	:douta	=	16'h	5b2d;
34102	:douta	=	16'h	5b2e;
34103	:douta	=	16'h	5b4e;
34104	:douta	=	16'h	636f;
34105	:douta	=	16'h	6bd0;
34106	:douta	=	16'h	5b2e;
34107	:douta	=	16'h	6bf1;
34108	:douta	=	16'h	63d0;
34109	:douta	=	16'h	4b2f;
34110	:douta	=	16'h	5b6e;
34111	:douta	=	16'h	acd2;
34112	:douta	=	16'h	bcf2;
34113	:douta	=	16'h	acb2;
34114	:douta	=	16'h	acb2;
34115	:douta	=	16'h	acd3;
34116	:douta	=	16'h	9cb4;
34117	:douta	=	16'h	8c73;
34118	:douta	=	16'h	8c53;
34119	:douta	=	16'h	736e;
34120	:douta	=	16'h	6b2d;
34121	:douta	=	16'h	62cd;
34122	:douta	=	16'h	630d;
34123	:douta	=	16'h	4a2b;
34124	:douta	=	16'h	936a;
34125	:douta	=	16'h	bc6b;
34126	:douta	=	16'h	f6b5;
34127	:douta	=	16'h	d571;
34128	:douta	=	16'h	ee75;
34129	:douta	=	16'h	bd10;
34130	:douta	=	16'h	ac4e;
34131	:douta	=	16'h	eeb7;
34132	:douta	=	16'h	ddd2;
34133	:douta	=	16'h	ddd2;
34134	:douta	=	16'h	cdb3;
34135	:douta	=	16'h	cdb4;
34136	:douta	=	16'h	bd54;
34137	:douta	=	16'h	acf4;
34138	:douta	=	16'h	a4b4;
34139	:douta	=	16'h	9493;
34140	:douta	=	16'h	8c53;
34141	:douta	=	16'h	7bd1;
34142	:douta	=	16'h	73b0;
34143	:douta	=	16'h	734e;
34144	:douta	=	16'h	6b2d;
34145	:douta	=	16'h	6b2e;
34146	:douta	=	16'h	526d;
34147	:douta	=	16'h	422b;
34148	:douta	=	16'h	39ea;
34149	:douta	=	16'h	2189;
34150	:douta	=	16'h	4209;
34151	:douta	=	16'h	ac0c;
34152	:douta	=	16'h	d56f;
34153	:douta	=	16'h	e654;
34154	:douta	=	16'h	eeb7;
34155	:douta	=	16'h	ee75;
34156	:douta	=	16'h	d5d5;
34157	:douta	=	16'h	c533;
34158	:douta	=	16'h	ad14;
34159	:douta	=	16'h	a4d4;
34160	:douta	=	16'h	bd54;
34161	:douta	=	16'h	8432;
34162	:douta	=	16'h	9452;
34163	:douta	=	16'h	9473;
34164	:douta	=	16'h	8c32;
34165	:douta	=	16'h	8433;
34166	:douta	=	16'h	8c52;
34167	:douta	=	16'h	8432;
34168	:douta	=	16'h	734e;
34169	:douta	=	16'h	83f0;
34170	:douta	=	16'h	8c31;
34171	:douta	=	16'h	83b0;
34172	:douta	=	16'h	7bb0;
34173	:douta	=	16'h	7b6f;
34174	:douta	=	16'h	5a8c;
34175	:douta	=	16'h	6b0c;
34176	:douta	=	16'h	bd11;
34177	:douta	=	16'h	e5d4;
34178	:douta	=	16'h	ddf4;
34179	:douta	=	16'h	bd12;
34180	:douta	=	16'h	d593;
34181	:douta	=	16'h	9495;
34182	:douta	=	16'h	63b1;
34183	:douta	=	16'h	a4b3;
34184	:douta	=	16'h	9c73;
34185	:douta	=	16'h	9c74;
34186	:douta	=	16'h	8c12;
34187	:douta	=	16'h	8c12;
34188	:douta	=	16'h	8bf1;
34189	:douta	=	16'h	9452;
34190	:douta	=	16'h	8c31;
34191	:douta	=	16'h	83f0;
34192	:douta	=	16'h	7bcf;
34193	:douta	=	16'h	7b6e;
34194	:douta	=	16'h	7b6e;
34195	:douta	=	16'h	7b4d;
34196	:douta	=	16'h	732c;
34197	:douta	=	16'h	730c;
34198	:douta	=	16'h	628a;
34199	:douta	=	16'h	732d;
34200	:douta	=	16'h	83af;
34201	:douta	=	16'h	b535;
34202	:douta	=	16'h	bd75;
34203	:douta	=	16'h	a4b4;
34204	:douta	=	16'h	9474;
34205	:douta	=	16'h	9453;
34206	:douta	=	16'h	8c12;
34207	:douta	=	16'h	8bf1;
34208	:douta	=	16'h	8411;
34209	:douta	=	16'h	83d0;
34210	:douta	=	16'h	83f1;
34211	:douta	=	16'h	83d0;
34212	:douta	=	16'h	7b90;
34213	:douta	=	16'h	7b6f;
34214	:douta	=	16'h	734f;
34215	:douta	=	16'h	6b2f;
34216	:douta	=	16'h	5aed;
34217	:douta	=	16'h	52cc;
34218	:douta	=	16'h	632f;
34219	:douta	=	16'h	73d0;
34220	:douta	=	16'h	9474;
34221	:douta	=	16'h	8412;
34222	:douta	=	16'h	8412;
34223	:douta	=	16'h	83f1;
34224	:douta	=	16'h	83f1;
34225	:douta	=	16'h	7bd1;
34226	:douta	=	16'h	7390;
34227	:douta	=	16'h	7390;
34228	:douta	=	16'h	6b6f;
34229	:douta	=	16'h	6b4f;
34230	:douta	=	16'h	5ace;
34231	:douta	=	16'h	52cd;
34232	:douta	=	16'h	5aee;
34233	:douta	=	16'h	4aad;
34234	:douta	=	16'h	4aad;
34235	:douta	=	16'h	4a8d;
34236	:douta	=	16'h	4a8d;
34237	:douta	=	16'h	5aee;
34238	:douta	=	16'h	d5b4;
34239	:douta	=	16'h	c575;
34240	:douta	=	16'h	7433;
34241	:douta	=	16'h	6bb2;
34242	:douta	=	16'h	6bb1;
34243	:douta	=	16'h	63b2;
34244	:douta	=	16'h	428e;
34245	:douta	=	16'h	4aae;
34246	:douta	=	16'h	2189;
34247	:douta	=	16'h	2189;
34248	:douta	=	16'h	2168;
34249	:douta	=	16'h	1906;
34250	:douta	=	16'h	320c;
34251	:douta	=	16'h	1906;
34252	:douta	=	16'h	18e5;
34253	:douta	=	16'h	10e5;
34254	:douta	=	16'h	10e5;
34255	:douta	=	16'h	10c5;
34256	:douta	=	16'h	10e5;
34257	:douta	=	16'h	10e5;
34258	:douta	=	16'h	21a9;
34259	:douta	=	16'h	5312;
34260	:douta	=	16'h	84d6;
34261	:douta	=	16'h	5bf3;
34262	:douta	=	16'h	6c15;
34263	:douta	=	16'h	8cf7;
34264	:douta	=	16'h	6c15;
34265	:douta	=	16'h	63f4;
34266	:douta	=	16'h	7c96;
34267	:douta	=	16'h	5393;
34268	:douta	=	16'h	6c55;
34269	:douta	=	16'h	8d39;
34270	:douta	=	16'h	5bd4;
34271	:douta	=	16'h	7cb7;
34272	:douta	=	16'h	6c56;
34273	:douta	=	16'h	6c35;
34274	:douta	=	16'h	7cb8;
34275	:douta	=	16'h	6c37;
34276	:douta	=	16'h	5393;
34277	:douta	=	16'h	6c57;
34278	:douta	=	16'h	6c56;
34279	:douta	=	16'h	855b;
34280	:douta	=	16'h	4b11;
34281	:douta	=	16'h	21c9;
34282	:douta	=	16'h	29ea;
34283	:douta	=	16'h	29ca;
34284	:douta	=	16'h	29eb;
34285	:douta	=	16'h	1947;
34286	:douta	=	16'h	5acc;
34287	:douta	=	16'h	5a69;
34288	:douta	=	16'h	5228;
34289	:douta	=	16'h	4a28;
34290	:douta	=	16'h	49e8;
34291	:douta	=	16'h	5228;
34292	:douta	=	16'h	4a08;
34293	:douta	=	16'h	5229;
34294	:douta	=	16'h	49e7;
34295	:douta	=	16'h	5228;
34296	:douta	=	16'h	5228;
34297	:douta	=	16'h	5208;
34298	:douta	=	16'h	5228;
34299	:douta	=	16'h	49e8;
34300	:douta	=	16'h	4a08;
34301	:douta	=	16'h	4a08;
34302	:douta	=	16'h	4a08;
34303	:douta	=	16'h	49c7;
34304	:douta	=	16'h	e56c;
34305	:douta	=	16'h	dd4b;
34306	:douta	=	16'h	dd4b;
34307	:douta	=	16'h	ccea;
34308	:douta	=	16'h	3945;
34309	:douta	=	16'h	3965;
34310	:douta	=	16'h	5acb;
34311	:douta	=	16'h	6b6f;
34312	:douta	=	16'h	3945;
34313	:douta	=	16'h	3924;
34314	:douta	=	16'h	3124;
34315	:douta	=	16'h	10a3;
34316	:douta	=	16'h	10c4;
34317	:douta	=	16'h	10c4;
34318	:douta	=	16'h	1083;
34319	:douta	=	16'h	1083;
34320	:douta	=	16'h	10a3;
34321	:douta	=	16'h	1083;
34322	:douta	=	16'h	1906;
34323	:douta	=	16'h	320b;
34324	:douta	=	16'h	31eb;
34325	:douta	=	16'h	322b;
34326	:douta	=	16'h	3a2c;
34327	:douta	=	16'h	31ea;
34328	:douta	=	16'h	320b;
34329	:douta	=	16'h	3a4c;
34330	:douta	=	16'h	428d;
34331	:douta	=	16'h	42ad;
34332	:douta	=	16'h	4aee;
34333	:douta	=	16'h	532f;
34334	:douta	=	16'h	532f;
34335	:douta	=	16'h	532f;
34336	:douta	=	16'h	530e;
34337	:douta	=	16'h	532f;
34338	:douta	=	16'h	532f;
34339	:douta	=	16'h	42cd;
34340	:douta	=	16'h	4aed;
34341	:douta	=	16'h	4b0d;
34342	:douta	=	16'h	4b0d;
34343	:douta	=	16'h	532e;
34344	:douta	=	16'h	532e;
34345	:douta	=	16'h	4aed;
34346	:douta	=	16'h	532e;
34347	:douta	=	16'h	532e;
34348	:douta	=	16'h	4b0d;
34349	:douta	=	16'h	532d;
34350	:douta	=	16'h	530d;
34351	:douta	=	16'h	4aac;
34352	:douta	=	16'h	52ed;
34353	:douta	=	16'h	52ec;
34354	:douta	=	16'h	530d;
34355	:douta	=	16'h	5b2e;
34356	:douta	=	16'h	5b4e;
34357	:douta	=	16'h	5b4e;
34358	:douta	=	16'h	638f;
34359	:douta	=	16'h	638f;
34360	:douta	=	16'h	638f;
34361	:douta	=	16'h	636f;
34362	:douta	=	16'h	636f;
34363	:douta	=	16'h	63d0;
34364	:douta	=	16'h	63b0;
34365	:douta	=	16'h	63af;
34366	:douta	=	16'h	5bb0;
34367	:douta	=	16'h	638f;
34368	:douta	=	16'h	9c50;
34369	:douta	=	16'h	acb1;
34370	:douta	=	16'h	a491;
34371	:douta	=	16'h	a492;
34372	:douta	=	16'h	8c51;
34373	:douta	=	16'h	8411;
34374	:douta	=	16'h	7bb0;
34375	:douta	=	16'h	736e;
34376	:douta	=	16'h	732e;
34377	:douta	=	16'h	6b2c;
34378	:douta	=	16'h	4a0a;
34379	:douta	=	16'h	6a8a;
34380	:douta	=	16'h	d52f;
34381	:douta	=	16'h	c4ed;
34382	:douta	=	16'h	eeb7;
34383	:douta	=	16'h	e634;
34384	:douta	=	16'h	f6f7;
34385	:douta	=	16'h	bd10;
34386	:douta	=	16'h	ac4e;
34387	:douta	=	16'h	ee75;
34388	:douta	=	16'h	cd92;
34389	:douta	=	16'h	d573;
34390	:douta	=	16'h	cd73;
34391	:douta	=	16'h	c532;
34392	:douta	=	16'h	b514;
34393	:douta	=	16'h	acf4;
34394	:douta	=	16'h	9cb3;
34395	:douta	=	16'h	8c73;
34396	:douta	=	16'h	8452;
34397	:douta	=	16'h	7bf1;
34398	:douta	=	16'h	73b0;
34399	:douta	=	16'h	6b6e;
34400	:douta	=	16'h	734e;
34401	:douta	=	16'h	6b2d;
34402	:douta	=	16'h	6b0d;
34403	:douta	=	16'h	6acd;
34404	:douta	=	16'h	5aac;
34405	:douta	=	16'h	5a49;
34406	:douta	=	16'h	a3cb;
34407	:douta	=	16'h	ddf3;
34408	:douta	=	16'h	eeb6;
34409	:douta	=	16'h	cd72;
34410	:douta	=	16'h	ee96;
34411	:douta	=	16'h	de14;
34412	:douta	=	16'h	bd74;
34413	:douta	=	16'h	b554;
34414	:douta	=	16'h	8c34;
34415	:douta	=	16'h	a4f4;
34416	:douta	=	16'h	acf5;
34417	:douta	=	16'h	8c33;
34418	:douta	=	16'h	632f;
34419	:douta	=	16'h	8c31;
34420	:douta	=	16'h	83d0;
34421	:douta	=	16'h	83af;
34422	:douta	=	16'h	8bf1;
34423	:douta	=	16'h	8bf1;
34424	:douta	=	16'h	732e;
34425	:douta	=	16'h	734e;
34426	:douta	=	16'h	83f0;
34427	:douta	=	16'h	83b0;
34428	:douta	=	16'h	83d0;
34429	:douta	=	16'h	630d;
34430	:douta	=	16'h	8bce;
34431	:douta	=	16'h	bcd0;
34432	:douta	=	16'h	f6b5;
34433	:douta	=	16'h	a493;
34434	:douta	=	16'h	e636;
34435	:douta	=	16'h	bd12;
34436	:douta	=	16'h	c533;
34437	:douta	=	16'h	9cd5;
34438	:douta	=	16'h	8454;
34439	:douta	=	16'h	5b10;
34440	:douta	=	16'h	a4b3;
34441	:douta	=	16'h	9c53;
34442	:douta	=	16'h	8bf2;
34443	:douta	=	16'h	8bf1;
34444	:douta	=	16'h	8bf0;
34445	:douta	=	16'h	838e;
34446	:douta	=	16'h	7b8e;
34447	:douta	=	16'h	7b8e;
34448	:douta	=	16'h	7b6e;
34449	:douta	=	16'h	7b6e;
34450	:douta	=	16'h	732d;
34451	:douta	=	16'h	732d;
34452	:douta	=	16'h	6aec;
34453	:douta	=	16'h	62aa;
34454	:douta	=	16'h	8bd0;
34455	:douta	=	16'h	ad14;
34456	:douta	=	16'h	b535;
34457	:douta	=	16'h	8c32;
34458	:douta	=	16'h	83f1;
34459	:douta	=	16'h	8c32;
34460	:douta	=	16'h	8c32;
34461	:douta	=	16'h	8c32;
34462	:douta	=	16'h	83f1;
34463	:douta	=	16'h	7b90;
34464	:douta	=	16'h	7b90;
34465	:douta	=	16'h	7b6f;
34466	:douta	=	16'h	736e;
34467	:douta	=	16'h	7bd0;
34468	:douta	=	16'h	7bb0;
34469	:douta	=	16'h	6b4e;
34470	:douta	=	16'h	5ace;
34471	:douta	=	16'h	5aad;
34472	:douta	=	16'h	632e;
34473	:douta	=	16'h	83d1;
34474	:douta	=	16'h	9cb5;
34475	:douta	=	16'h	9474;
34476	:douta	=	16'h	8c53;
34477	:douta	=	16'h	a494;
34478	:douta	=	16'h	a493;
34479	:douta	=	16'h	8c32;
34480	:douta	=	16'h	8c32;
34481	:douta	=	16'h	83f1;
34482	:douta	=	16'h	6b4e;
34483	:douta	=	16'h	6b4f;
34484	:douta	=	16'h	6b4f;
34485	:douta	=	16'h	632e;
34486	:douta	=	16'h	630f;
34487	:douta	=	16'h	5aee;
34488	:douta	=	16'h	5acd;
34489	:douta	=	16'h	52cd;
34490	:douta	=	16'h	4a6c;
34491	:douta	=	16'h	4a8c;
34492	:douta	=	16'h	9451;
34493	:douta	=	16'h	cdb4;
34494	:douta	=	16'h	b534;
34495	:douta	=	16'h	94b5;
34496	:douta	=	16'h	8434;
34497	:douta	=	16'h	7c54;
34498	:douta	=	16'h	7433;
34499	:douta	=	16'h	5330;
34500	:douta	=	16'h	4aae;
34501	:douta	=	16'h	5331;
34502	:douta	=	16'h	29a9;
34503	:douta	=	16'h	320b;
34504	:douta	=	16'h	2189;
34505	:douta	=	16'h	29eb;
34506	:douta	=	16'h	18e5;
34507	:douta	=	16'h	428e;
34508	:douta	=	16'h	29c9;
34509	:douta	=	16'h	1906;
34510	:douta	=	16'h	10e5;
34511	:douta	=	16'h	10e5;
34512	:douta	=	16'h	10e6;
34513	:douta	=	16'h	1926;
34514	:douta	=	16'h	10c4;
34515	:douta	=	16'h	29a9;
34516	:douta	=	16'h	7496;
34517	:douta	=	16'h	7435;
34518	:douta	=	16'h	9517;
34519	:douta	=	16'h	5394;
34520	:douta	=	16'h	6c15;
34521	:douta	=	16'h	7455;
34522	:douta	=	16'h	63f4;
34523	:douta	=	16'h	6c55;
34524	:douta	=	16'h	9539;
34525	:douta	=	16'h	7cb8;
34526	:douta	=	16'h	84b7;
34527	:douta	=	16'h	6c35;
34528	:douta	=	16'h	4b32;
34529	:douta	=	16'h	6c56;
34530	:douta	=	16'h	5bd4;
34531	:douta	=	16'h	7cb8;
34532	:douta	=	16'h	53d4;
34533	:douta	=	16'h	7457;
34534	:douta	=	16'h	6457;
34535	:douta	=	16'h	6436;
34536	:douta	=	16'h	2188;
34537	:douta	=	16'h	2189;
34538	:douta	=	16'h	29aa;
34539	:douta	=	16'h	29a9;
34540	:douta	=	16'h	29ca;
34541	:douta	=	16'h	29c9;
34542	:douta	=	16'h	2168;
34543	:douta	=	16'h	39e9;
34544	:douta	=	16'h	6aaa;
34545	:douta	=	16'h	5a49;
34546	:douta	=	16'h	5208;
34547	:douta	=	16'h	5a49;
34548	:douta	=	16'h	5229;
34549	:douta	=	16'h	5208;
34550	:douta	=	16'h	49e8;
34551	:douta	=	16'h	5208;
34552	:douta	=	16'h	5249;
34553	:douta	=	16'h	5249;
34554	:douta	=	16'h	4a08;
34555	:douta	=	16'h	5208;
34556	:douta	=	16'h	49e8;
34557	:douta	=	16'h	4a08;
34558	:douta	=	16'h	5208;
34559	:douta	=	16'h	49c7;
34560	:douta	=	16'h	e56c;
34561	:douta	=	16'h	dd4b;
34562	:douta	=	16'h	e54c;
34563	:douta	=	16'h	edec;
34564	:douta	=	16'h	28e4;
34565	:douta	=	16'h	4165;
34566	:douta	=	16'h	4985;
34567	:douta	=	16'h	7bd1;
34568	:douta	=	16'h	3903;
34569	:douta	=	16'h	4165;
34570	:douta	=	16'h	28e3;
34571	:douta	=	16'h	10a3;
34572	:douta	=	16'h	10c4;
34573	:douta	=	16'h	1905;
34574	:douta	=	16'h	2146;
34575	:douta	=	16'h	2146;
34576	:douta	=	16'h	2125;
34577	:douta	=	16'h	2105;
34578	:douta	=	16'h	29ca;
34579	:douta	=	16'h	29ea;
34580	:douta	=	16'h	31eb;
34581	:douta	=	16'h	322b;
34582	:douta	=	16'h	3a2b;
34583	:douta	=	16'h	29ea;
34584	:douta	=	16'h	3a4c;
34585	:douta	=	16'h	428d;
34586	:douta	=	16'h	42ae;
34587	:douta	=	16'h	4ace;
34588	:douta	=	16'h	4aae;
34589	:douta	=	16'h	4ace;
34590	:douta	=	16'h	530f;
34591	:douta	=	16'h	530e;
34592	:douta	=	16'h	4aee;
34593	:douta	=	16'h	530e;
34594	:douta	=	16'h	4b0e;
34595	:douta	=	16'h	3a6b;
34596	:douta	=	16'h	42ac;
34597	:douta	=	16'h	4aad;
34598	:douta	=	16'h	4b0d;
34599	:douta	=	16'h	530e;
34600	:douta	=	16'h	4b0d;
34601	:douta	=	16'h	530e;
34602	:douta	=	16'h	534e;
34603	:douta	=	16'h	4aed;
34604	:douta	=	16'h	4b0d;
34605	:douta	=	16'h	4aed;
34606	:douta	=	16'h	52ed;
34607	:douta	=	16'h	4acc;
34608	:douta	=	16'h	4aac;
34609	:douta	=	16'h	4aac;
34610	:douta	=	16'h	4aac;
34611	:douta	=	16'h	4aac;
34612	:douta	=	16'h	52ed;
34613	:douta	=	16'h	5b2e;
34614	:douta	=	16'h	5b4e;
34615	:douta	=	16'h	636f;
34616	:douta	=	16'h	638f;
34617	:douta	=	16'h	5b6f;
34618	:douta	=	16'h	6bf0;
34619	:douta	=	16'h	63d0;
34620	:douta	=	16'h	63af;
34621	:douta	=	16'h	63d0;
34622	:douta	=	16'h	63d0;
34623	:douta	=	16'h	63d0;
34624	:douta	=	16'h	5bb0;
34625	:douta	=	16'h	536f;
34626	:douta	=	16'h	6bb0;
34627	:douta	=	16'h	7bd0;
34628	:douta	=	16'h	9451;
34629	:douta	=	16'h	9411;
34630	:douta	=	16'h	8c11;
34631	:douta	=	16'h	6b2d;
34632	:douta	=	16'h	6b2d;
34633	:douta	=	16'h	39c8;
34634	:douta	=	16'h	d54f;
34635	:douta	=	16'h	bcae;
34636	:douta	=	16'h	ee95;
34637	:douta	=	16'h	e614;
34638	:douta	=	16'h	cd50;
34639	:douta	=	16'h	f759;
34640	:douta	=	16'h	eeb6;
34641	:douta	=	16'h	b4f1;
34642	:douta	=	16'h	9410;
34643	:douta	=	16'h	e675;
34644	:douta	=	16'h	c552;
34645	:douta	=	16'h	b4d3;
34646	:douta	=	16'h	a4b3;
34647	:douta	=	16'h	9c93;
34648	:douta	=	16'h	83f2;
34649	:douta	=	16'h	83f1;
34650	:douta	=	16'h	7bf1;
34651	:douta	=	16'h	7bd1;
34652	:douta	=	16'h	7bb0;
34653	:douta	=	16'h	734e;
34654	:douta	=	16'h	732e;
34655	:douta	=	16'h	6b2d;
34656	:douta	=	16'h	62ec;
34657	:douta	=	16'h	62cc;
34658	:douta	=	16'h	5aac;
34659	:douta	=	16'h	4a4b;
34660	:douta	=	16'h	9b6b;
34661	:douta	=	16'h	e613;
34662	:douta	=	16'h	ee76;
34663	:douta	=	16'h	e674;
34664	:douta	=	16'h	e635;
34665	:douta	=	16'h	d5f5;
34666	:douta	=	16'h	bd53;
34667	:douta	=	16'h	bd54;
34668	:douta	=	16'h	a4d5;
34669	:douta	=	16'h	a515;
34670	:douta	=	16'h	a516;
34671	:douta	=	16'h	8c94;
34672	:douta	=	16'h	7c33;
34673	:douta	=	16'h	9453;
34674	:douta	=	16'h	94b3;
34675	:douta	=	16'h	632f;
34676	:douta	=	16'h	4ace;
34677	:douta	=	16'h	5b0e;
34678	:douta	=	16'h	7b6f;
34679	:douta	=	16'h	838f;
34680	:douta	=	16'h	8bd0;
34681	:douta	=	16'h	838f;
34682	:douta	=	16'h	62ed;
34683	:douta	=	16'h	5a6c;
34684	:douta	=	16'h	8b6d;
34685	:douta	=	16'h	f6b6;
34686	:douta	=	16'h	acb2;
34687	:douta	=	16'h	e655;
34688	:douta	=	16'h	cd93;
34689	:douta	=	16'h	b514;
34690	:douta	=	16'h	5b50;
34691	:douta	=	16'h	8453;
34692	:douta	=	16'h	8c95;
34693	:douta	=	16'h	94b5;
34694	:douta	=	16'h	8454;
34695	:douta	=	16'h	6b91;
34696	:douta	=	16'h	5b50;
34697	:douta	=	16'h	6371;
34698	:douta	=	16'h	83f1;
34699	:douta	=	16'h	9430;
34700	:douta	=	16'h	83ae;
34701	:douta	=	16'h	732d;
34702	:douta	=	16'h	730d;
34703	:douta	=	16'h	6aec;
34704	:douta	=	16'h	6aec;
34705	:douta	=	16'h	5249;
34706	:douta	=	16'h	8bf0;
34707	:douta	=	16'h	8c11;
34708	:douta	=	16'h	73d0;
34709	:douta	=	16'h	6b70;
34710	:douta	=	16'h	7bf2;
34711	:douta	=	16'h	8412;
34712	:douta	=	16'h	8bf1;
34713	:douta	=	16'h	7baf;
34714	:douta	=	16'h	83b0;
34715	:douta	=	16'h	736f;
34716	:douta	=	16'h	6b2f;
34717	:douta	=	16'h	736f;
34718	:douta	=	16'h	83b0;
34719	:douta	=	16'h	7b8f;
34720	:douta	=	16'h	7b8f;
34721	:douta	=	16'h	62ee;
34722	:douta	=	16'h	62ee;
34723	:douta	=	16'h	6b4e;
34724	:douta	=	16'h	736f;
34725	:douta	=	16'h	a493;
34726	:douta	=	16'h	c593;
34727	:douta	=	16'h	cdd4;
34728	:douta	=	16'h	bd35;
34729	:douta	=	16'h	a4d4;
34730	:douta	=	16'h	9473;
34731	:douta	=	16'h	8c53;
34732	:douta	=	16'h	8433;
34733	:douta	=	16'h	8c53;
34734	:douta	=	16'h	9c94;
34735	:douta	=	16'h	8c52;
34736	:douta	=	16'h	8431;
34737	:douta	=	16'h	73b0;
34738	:douta	=	16'h	6b6f;
34739	:douta	=	16'h	7390;
34740	:douta	=	16'h	73b1;
34741	:douta	=	16'h	73b0;
34742	:douta	=	16'h	6b6f;
34743	:douta	=	16'h	632e;
34744	:douta	=	16'h	632e;
34745	:douta	=	16'h	7b6e;
34746	:douta	=	16'h	acf3;
34747	:douta	=	16'h	d5d5;
34748	:douta	=	16'h	cdb5;
34749	:douta	=	16'h	c554;
34750	:douta	=	16'h	ad15;
34751	:douta	=	16'h	9cf5;
34752	:douta	=	16'h	8c95;
34753	:douta	=	16'h	8474;
34754	:douta	=	16'h	7c35;
34755	:douta	=	16'h	6bb2;
34756	:douta	=	16'h	6372;
34757	:douta	=	16'h	4b10;
34758	:douta	=	16'h	4af0;
34759	:douta	=	16'h	3a2c;
34760	:douta	=	16'h	42ae;
34761	:douta	=	16'h	3a8d;
34762	:douta	=	16'h	29ca;
34763	:douta	=	16'h	2168;
34764	:douta	=	16'h	1948;
34765	:douta	=	16'h	5b31;
34766	:douta	=	16'h	29ca;
34767	:douta	=	16'h	2126;
34768	:douta	=	16'h	2147;
34769	:douta	=	16'h	2168;
34770	:douta	=	16'h	10c5;
34771	:douta	=	16'h	1905;
34772	:douta	=	16'h	0000;
34773	:douta	=	16'h	5b93;
34774	:douta	=	16'h	7cb7;
34775	:douta	=	16'h	8cf6;
34776	:douta	=	16'h	9d79;
34777	:douta	=	16'h	6c14;
34778	:douta	=	16'h	9d59;
34779	:douta	=	16'h	8cf8;
34780	:douta	=	16'h	7cb7;
34781	:douta	=	16'h	84d8;
34782	:douta	=	16'h	5373;
34783	:douta	=	16'h	7c75;
34784	:douta	=	16'h	7cb7;
34785	:douta	=	16'h	5bb4;
34786	:douta	=	16'h	5bb4;
34787	:douta	=	16'h	5bf5;
34788	:douta	=	16'h	8519;
34789	:douta	=	16'h	84f9;
34790	:douta	=	16'h	4311;
34791	:douta	=	16'h	1926;
34792	:douta	=	16'h	320b;
34793	:douta	=	16'h	29ca;
34794	:douta	=	16'h	29a9;
34795	:douta	=	16'h	21a9;
34796	:douta	=	16'h	2188;
34797	:douta	=	16'h	31c9;
34798	:douta	=	16'h	29c9;
34799	:douta	=	16'h	29c9;
34800	:douta	=	16'h	21aa;
34801	:douta	=	16'h	320a;
34802	:douta	=	16'h	6aaa;
34803	:douta	=	16'h	49c7;
34804	:douta	=	16'h	49e8;
34805	:douta	=	16'h	5249;
34806	:douta	=	16'h	5249;
34807	:douta	=	16'h	5229;
34808	:douta	=	16'h	5229;
34809	:douta	=	16'h	5228;
34810	:douta	=	16'h	5208;
34811	:douta	=	16'h	49e8;
34812	:douta	=	16'h	5208;
34813	:douta	=	16'h	49e8;
34814	:douta	=	16'h	49e8;
34815	:douta	=	16'h	49e8;
34816	:douta	=	16'h	e56c;
34817	:douta	=	16'h	dd4b;
34818	:douta	=	16'h	dd4b;
34819	:douta	=	16'h	f5cc;
34820	:douta	=	16'h	28e4;
34821	:douta	=	16'h	3945;
34822	:douta	=	16'h	3923;
34823	:douta	=	16'h	7b90;
34824	:douta	=	16'h	3923;
34825	:douta	=	16'h	3965;
34826	:douta	=	16'h	20e4;
34827	:douta	=	16'h	0861;
34828	:douta	=	16'h	08a2;
34829	:douta	=	16'h	10a4;
34830	:douta	=	16'h	2105;
34831	:douta	=	16'h	10c4;
34832	:douta	=	16'h	1084;
34833	:douta	=	16'h	1083;
34834	:douta	=	16'h	1948;
34835	:douta	=	16'h	320b;
34836	:douta	=	16'h	29ea;
34837	:douta	=	16'h	320b;
34838	:douta	=	16'h	3a2c;
34839	:douta	=	16'h	29aa;
34840	:douta	=	16'h	320b;
34841	:douta	=	16'h	3a4c;
34842	:douta	=	16'h	42ad;
34843	:douta	=	16'h	42ad;
34844	:douta	=	16'h	4aee;
34845	:douta	=	16'h	4aee;
34846	:douta	=	16'h	4b0e;
34847	:douta	=	16'h	4ace;
34848	:douta	=	16'h	4ace;
34849	:douta	=	16'h	530e;
34850	:douta	=	16'h	4acd;
34851	:douta	=	16'h	3a6c;
34852	:douta	=	16'h	428c;
34853	:douta	=	16'h	42ac;
34854	:douta	=	16'h	4acd;
34855	:douta	=	16'h	4b0e;
34856	:douta	=	16'h	4aed;
34857	:douta	=	16'h	4aed;
34858	:douta	=	16'h	532e;
34859	:douta	=	16'h	4b0e;
34860	:douta	=	16'h	4acd;
34861	:douta	=	16'h	4acd;
34862	:douta	=	16'h	4aac;
34863	:douta	=	16'h	428b;
34864	:douta	=	16'h	52ed;
34865	:douta	=	16'h	4aac;
34866	:douta	=	16'h	4aac;
34867	:douta	=	16'h	4aac;
34868	:douta	=	16'h	426b;
34869	:douta	=	16'h	530d;
34870	:douta	=	16'h	4acc;
34871	:douta	=	16'h	5b2e;
34872	:douta	=	16'h	5b2e;
34873	:douta	=	16'h	636f;
34874	:douta	=	16'h	63f0;
34875	:douta	=	16'h	5b6f;
34876	:douta	=	16'h	63b0;
34877	:douta	=	16'h	63af;
34878	:douta	=	16'h	63b0;
34879	:douta	=	16'h	63af;
34880	:douta	=	16'h	63b0;
34881	:douta	=	16'h	5b6f;
34882	:douta	=	16'h	5b90;
34883	:douta	=	16'h	5b90;
34884	:douta	=	16'h	6b8f;
34885	:douta	=	16'h	8bd0;
34886	:douta	=	16'h	8410;
34887	:douta	=	16'h	734e;
34888	:douta	=	16'h	422c;
34889	:douta	=	16'h	7ae9;
34890	:douta	=	16'h	d613;
34891	:douta	=	16'h	ac2b;
34892	:douta	=	16'h	f739;
34893	:douta	=	16'h	e675;
34894	:douta	=	16'h	ac6f;
34895	:douta	=	16'h	fef7;
34896	:douta	=	16'h	ee75;
34897	:douta	=	16'h	bd32;
34898	:douta	=	16'h	8bf1;
34899	:douta	=	16'h	d5d3;
34900	:douta	=	16'h	bd51;
34901	:douta	=	16'h	acd2;
34902	:douta	=	16'h	9c93;
34903	:douta	=	16'h	8c53;
34904	:douta	=	16'h	73b0;
34905	:douta	=	16'h	7b6f;
34906	:douta	=	16'h	736e;
34907	:douta	=	16'h	736f;
34908	:douta	=	16'h	734e;
34909	:douta	=	16'h	6b2d;
34910	:douta	=	16'h	6b0d;
34911	:douta	=	16'h	6b2d;
34912	:douta	=	16'h	62ec;
34913	:douta	=	16'h	62ec;
34914	:douta	=	16'h	420a;
34915	:douta	=	16'h	832b;
34916	:douta	=	16'h	ee12;
34917	:douta	=	16'h	ac91;
34918	:douta	=	16'h	e614;
34919	:douta	=	16'h	cdd3;
34920	:douta	=	16'h	bd33;
34921	:douta	=	16'h	c574;
34922	:douta	=	16'h	acf4;
34923	:douta	=	16'h	acf4;
34924	:douta	=	16'h	a515;
34925	:douta	=	16'h	94b5;
34926	:douta	=	16'h	9cd5;
34927	:douta	=	16'h	8474;
34928	:douta	=	16'h	8453;
34929	:douta	=	16'h	73d1;
34930	:douta	=	16'h	8432;
34931	:douta	=	16'h	83f1;
34932	:douta	=	16'h	5b0e;
34933	:douta	=	16'h	4aad;
34934	:douta	=	16'h	424c;
34935	:douta	=	16'h	4a8c;
34936	:douta	=	16'h	52ac;
34937	:douta	=	16'h	4a2c;
34938	:douta	=	16'h	524b;
34939	:douta	=	16'h	d572;
34940	:douta	=	16'h	f674;
34941	:douta	=	16'h	e614;
34942	:douta	=	16'h	73d2;
34943	:douta	=	16'h	b4f3;
34944	:douta	=	16'h	ad13;
34945	:douta	=	16'h	a4b4;
34946	:douta	=	16'h	7c95;
34947	:douta	=	16'h	6b91;
34948	:douta	=	16'h	6bd2;
34949	:douta	=	16'h	8412;
34950	:douta	=	16'h	7bd1;
34951	:douta	=	16'h	7b90;
34952	:douta	=	16'h	7390;
34953	:douta	=	16'h	7391;
34954	:douta	=	16'h	5b2f;
34955	:douta	=	16'h	630e;
34956	:douta	=	16'h	734d;
34957	:douta	=	16'h	62cc;
34958	:douta	=	16'h	5aac;
34959	:douta	=	16'h	420a;
34960	:douta	=	16'h	39a8;
34961	:douta	=	16'h	734e;
34962	:douta	=	16'h	ad15;
34963	:douta	=	16'h	9cb4;
34964	:douta	=	16'h	8454;
34965	:douta	=	16'h	7c54;
34966	:douta	=	16'h	7bf3;
34967	:douta	=	16'h	7bf2;
34968	:douta	=	16'h	8411;
34969	:douta	=	16'h	7b90;
34970	:douta	=	16'h	738f;
34971	:douta	=	16'h	7baf;
34972	:douta	=	16'h	6b2e;
34973	:douta	=	16'h	62ed;
34974	:douta	=	16'h	632e;
34975	:douta	=	16'h	6b4e;
34976	:douta	=	16'h	52ac;
34977	:douta	=	16'h	8c10;
34978	:douta	=	16'h	8bf0;
34979	:douta	=	16'h	b4f3;
34980	:douta	=	16'h	d5b4;
34981	:douta	=	16'h	9432;
34982	:douta	=	16'h	73b1;
34983	:douta	=	16'h	83f1;
34984	:douta	=	16'h	9c73;
34985	:douta	=	16'h	9c93;
34986	:douta	=	16'h	9493;
34987	:douta	=	16'h	8452;
34988	:douta	=	16'h	83f2;
34989	:douta	=	16'h	8432;
34990	:douta	=	16'h	9453;
34991	:douta	=	16'h	9453;
34992	:douta	=	16'h	8c12;
34993	:douta	=	16'h	73b0;
34994	:douta	=	16'h	6b4f;
34995	:douta	=	16'h	632e;
34996	:douta	=	16'h	632e;
34997	:douta	=	16'h	6b4f;
34998	:douta	=	16'h	5aee;
34999	:douta	=	16'h	630d;
35000	:douta	=	16'h	62ed;
35001	:douta	=	16'h	8bce;
35002	:douta	=	16'h	ac90;
35003	:douta	=	16'h	bd74;
35004	:douta	=	16'h	b534;
35005	:douta	=	16'h	b534;
35006	:douta	=	16'h	a515;
35007	:douta	=	16'h	9cd5;
35008	:douta	=	16'h	8cb5;
35009	:douta	=	16'h	7c54;
35010	:douta	=	16'h	73f3;
35011	:douta	=	16'h	6392;
35012	:douta	=	16'h	5b71;
35013	:douta	=	16'h	5b31;
35014	:douta	=	16'h	4ad0;
35015	:douta	=	16'h	320c;
35016	:douta	=	16'h	4acf;
35017	:douta	=	16'h	3a8e;
35018	:douta	=	16'h	21aa;
35019	:douta	=	16'h	29a9;
35020	:douta	=	16'h	29a9;
35021	:douta	=	16'h	4aad;
35022	:douta	=	16'h	6370;
35023	:douta	=	16'h	10e5;
35024	:douta	=	16'h	1927;
35025	:douta	=	16'h	2168;
35026	:douta	=	16'h	1946;
35027	:douta	=	16'h	10e5;
35028	:douta	=	16'h	10e5;
35029	:douta	=	16'h	08c6;
35030	:douta	=	16'h	7455;
35031	:douta	=	16'h	7c96;
35032	:douta	=	16'h	6bf3;
35033	:douta	=	16'h	9d58;
35034	:douta	=	16'h	9518;
35035	:douta	=	16'h	84b6;
35036	:douta	=	16'h	84b7;
35037	:douta	=	16'h	5bd3;
35038	:douta	=	16'h	7455;
35039	:douta	=	16'h	84d8;
35040	:douta	=	16'h	6c35;
35041	:douta	=	16'h	6c56;
35042	:douta	=	16'h	6c56;
35043	:douta	=	16'h	32b0;
35044	:douta	=	16'h	7497;
35045	:douta	=	16'h	53f5;
35046	:douta	=	16'h	31c9;
35047	:douta	=	16'h	2167;
35048	:douta	=	16'h	29c9;
35049	:douta	=	16'h	29a9;
35050	:douta	=	16'h	2188;
35051	:douta	=	16'h	29ca;
35052	:douta	=	16'h	29ea;
35053	:douta	=	16'h	320a;
35054	:douta	=	16'h	320b;
35055	:douta	=	16'h	3a4c;
35056	:douta	=	16'h	3a4c;
35057	:douta	=	16'h	2a2c;
35058	:douta	=	16'h	422a;
35059	:douta	=	16'h	5207;
35060	:douta	=	16'h	49e7;
35061	:douta	=	16'h	5228;
35062	:douta	=	16'h	5208;
35063	:douta	=	16'h	5229;
35064	:douta	=	16'h	5208;
35065	:douta	=	16'h	4a08;
35066	:douta	=	16'h	5208;
35067	:douta	=	16'h	5229;
35068	:douta	=	16'h	5208;
35069	:douta	=	16'h	49e8;
35070	:douta	=	16'h	49e8;
35071	:douta	=	16'h	5208;
35072	:douta	=	16'h	e56c;
35073	:douta	=	16'h	e56c;
35074	:douta	=	16'h	dd4c;
35075	:douta	=	16'h	e54b;
35076	:douta	=	16'h	5a47;
35077	:douta	=	16'h	3924;
35078	:douta	=	16'h	4144;
35079	:douta	=	16'h	628a;
35080	:douta	=	16'h	49c6;
35081	:douta	=	16'h	1861;
35082	:douta	=	16'h	4a4b;
35083	:douta	=	16'h	52ac;
35084	:douta	=	16'h	2105;
35085	:douta	=	16'h	31c8;
35086	:douta	=	16'h	0883;
35087	:douta	=	16'h	7b0c;
35088	:douta	=	16'h	a4b5;
35089	:douta	=	16'h	9d16;
35090	:douta	=	16'h	a598;
35091	:douta	=	16'h	29c9;
35092	:douta	=	16'h	29aa;
35093	:douta	=	16'h	320b;
35094	:douta	=	16'h	322b;
35095	:douta	=	16'h	29ca;
35096	:douta	=	16'h	322b;
35097	:douta	=	16'h	3a4c;
35098	:douta	=	16'h	428d;
35099	:douta	=	16'h	3a6d;
35100	:douta	=	16'h	42cd;
35101	:douta	=	16'h	4aee;
35102	:douta	=	16'h	42ce;
35103	:douta	=	16'h	4aee;
35104	:douta	=	16'h	4ace;
35105	:douta	=	16'h	4ace;
35106	:douta	=	16'h	42ad;
35107	:douta	=	16'h	322a;
35108	:douta	=	16'h	3a4b;
35109	:douta	=	16'h	3a6b;
35110	:douta	=	16'h	3a8c;
35111	:douta	=	16'h	428c;
35112	:douta	=	16'h	428c;
35113	:douta	=	16'h	4acd;
35114	:douta	=	16'h	532e;
35115	:douta	=	16'h	4b0e;
35116	:douta	=	16'h	4b0e;
35117	:douta	=	16'h	4aed;
35118	:douta	=	16'h	42ac;
35119	:douta	=	16'h	428b;
35120	:douta	=	16'h	4acc;
35121	:douta	=	16'h	4aac;
35122	:douta	=	16'h	4aac;
35123	:douta	=	16'h	52ed;
35124	:douta	=	16'h	52ed;
35125	:douta	=	16'h	4acc;
35126	:douta	=	16'h	5b2e;
35127	:douta	=	16'h	530d;
35128	:douta	=	16'h	5b6f;
35129	:douta	=	16'h	534e;
35130	:douta	=	16'h	5b6f;
35131	:douta	=	16'h	5b8f;
35132	:douta	=	16'h	5b6f;
35133	:douta	=	16'h	5b8f;
35134	:douta	=	16'h	63b0;
35135	:douta	=	16'h	5b8f;
35136	:douta	=	16'h	5b6f;
35137	:douta	=	16'h	63b0;
35138	:douta	=	16'h	63d0;
35139	:douta	=	16'h	63d0;
35140	:douta	=	16'h	6bd1;
35141	:douta	=	16'h	5b8f;
35142	:douta	=	16'h	6bd0;
35143	:douta	=	16'h	634f;
35144	:douta	=	16'h	cd52;
35145	:douta	=	16'h	bcd1;
35146	:douta	=	16'h	c571;
35147	:douta	=	16'h	c4f0;
35148	:douta	=	16'h	eeb6;
35149	:douta	=	16'h	f6b6;
35150	:douta	=	16'h	d5f4;
35151	:douta	=	16'h	c511;
35152	:douta	=	16'h	ddf3;
35153	:douta	=	16'h	cd52;
35154	:douta	=	16'h	a492;
35155	:douta	=	16'h	acb2;
35156	:douta	=	16'h	bd32;
35157	:douta	=	16'h	9c92;
35158	:douta	=	16'h	9473;
35159	:douta	=	16'h	8c53;
35160	:douta	=	16'h	7bd1;
35161	:douta	=	16'h	6b2e;
35162	:douta	=	16'h	732e;
35163	:douta	=	16'h	62ec;
35164	:douta	=	16'h	62ec;
35165	:douta	=	16'h	62cc;
35166	:douta	=	16'h	62cb;
35167	:douta	=	16'h	5a6a;
35168	:douta	=	16'h	526a;
35169	:douta	=	16'h	524a;
35170	:douta	=	16'h	dd50;
35171	:douta	=	16'h	e635;
35172	:douta	=	16'h	e655;
35173	:douta	=	16'h	7414;
35174	:douta	=	16'h	ad15;
35175	:douta	=	16'h	bd75;
35176	:douta	=	16'h	a4f5;
35177	:douta	=	16'h	94d5;
35178	:douta	=	16'h	9cf5;
35179	:douta	=	16'h	94d5;
35180	:douta	=	16'h	94b5;
35181	:douta	=	16'h	94b5;
35182	:douta	=	16'h	8453;
35183	:douta	=	16'h	8432;
35184	:douta	=	16'h	7c12;
35185	:douta	=	16'h	736f;
35186	:douta	=	16'h	732f;
35187	:douta	=	16'h	7b90;
35188	:douta	=	16'h	736f;
35189	:douta	=	16'h	7b6f;
35190	:douta	=	16'h	734d;
35191	:douta	=	16'h	62cd;
35192	:douta	=	16'h	62ad;
35193	:douta	=	16'h	d52f;
35194	:douta	=	16'h	e614;
35195	:douta	=	16'h	cd93;
35196	:douta	=	16'h	c572;
35197	:douta	=	16'h	a4d4;
35198	:douta	=	16'h	8c74;
35199	:douta	=	16'h	8c33;
35200	:douta	=	16'h	a4b4;
35201	:douta	=	16'h	8434;
35202	:douta	=	16'h	7bd2;
35203	:douta	=	16'h	73f1;
35204	:douta	=	16'h	6b4f;
35205	:douta	=	16'h	4a8d;
35206	:douta	=	16'h	5aef;
35207	:douta	=	16'h	7b8f;
35208	:douta	=	16'h	62cc;
35209	:douta	=	16'h	6acc;
35210	:douta	=	16'h	6b0d;
35211	:douta	=	16'h	732e;
35212	:douta	=	16'h	732d;
35213	:douta	=	16'h	5aab;
35214	:douta	=	16'h	6b2d;
35215	:douta	=	16'h	8bf1;
35216	:douta	=	16'h	9c93;
35217	:douta	=	16'h	7bf1;
35218	:douta	=	16'h	73b0;
35219	:douta	=	16'h	7b8f;
35220	:douta	=	16'h	6b2e;
35221	:douta	=	16'h	5aed;
35222	:douta	=	16'h	5aee;
35223	:douta	=	16'h	73b0;
35224	:douta	=	16'h	6b90;
35225	:douta	=	16'h	7bb0;
35226	:douta	=	16'h	83d0;
35227	:douta	=	16'h	734e;
35228	:douta	=	16'h	6b2e;
35229	:douta	=	16'h	52ac;
35230	:douta	=	16'h	5acd;
35231	:douta	=	16'h	9410;
35232	:douta	=	16'h	9cb4;
35233	:douta	=	16'h	ac93;
35234	:douta	=	16'h	bcf3;
35235	:douta	=	16'h	b4d3;
35236	:douta	=	16'h	9c94;
35237	:douta	=	16'h	8c53;
35238	:douta	=	16'h	7c12;
35239	:douta	=	16'h	8412;
35240	:douta	=	16'h	8c53;
35241	:douta	=	16'h	8412;
35242	:douta	=	16'h	7b90;
35243	:douta	=	16'h	7bd1;
35244	:douta	=	16'h	7bd1;
35245	:douta	=	16'h	7b90;
35246	:douta	=	16'h	6b0d;
35247	:douta	=	16'h	6b2e;
35248	:douta	=	16'h	6b4f;
35249	:douta	=	16'h	6b6f;
35250	:douta	=	16'h	6b4f;
35251	:douta	=	16'h	630e;
35252	:douta	=	16'h	52ac;
35253	:douta	=	16'h	9410;
35254	:douta	=	16'h	d5f4;
35255	:douta	=	16'h	e676;
35256	:douta	=	16'h	e697;
35257	:douta	=	16'h	e677;
35258	:douta	=	16'h	e676;
35259	:douta	=	16'h	de36;
35260	:douta	=	16'h	bd75;
35261	:douta	=	16'h	a515;
35262	:douta	=	16'h	94b5;
35263	:douta	=	16'h	8c74;
35264	:douta	=	16'h	8c74;
35265	:douta	=	16'h	73f2;
35266	:douta	=	16'h	6bb2;
35267	:douta	=	16'h	6391;
35268	:douta	=	16'h	5b31;
35269	:douta	=	16'h	5b30;
35270	:douta	=	16'h	5b51;
35271	:douta	=	16'h	5b30;
35272	:douta	=	16'h	3a4e;
35273	:douta	=	16'h	324d;
35274	:douta	=	16'h	324c;
35275	:douta	=	16'h	428e;
35276	:douta	=	16'h	2a0c;
35277	:douta	=	16'h	52ee;
35278	:douta	=	16'h	1928;
35279	:douta	=	16'h	2146;
35280	:douta	=	16'h	1905;
35281	:douta	=	16'h	18e4;
35282	:douta	=	16'h	1905;
35283	:douta	=	16'h	10c4;
35284	:douta	=	16'h	10e5;
35285	:douta	=	16'h	2168;
35286	:douta	=	16'h	0063;
35287	:douta	=	16'h	84d7;
35288	:douta	=	16'h	9d78;
35289	:douta	=	16'h	8495;
35290	:douta	=	16'h	84d6;
35291	:douta	=	16'h	7435;
35292	:douta	=	16'h	5b73;
35293	:douta	=	16'h	63f4;
35294	:douta	=	16'h	5bd4;
35295	:douta	=	16'h	7456;
35296	:douta	=	16'h	84d7;
35297	:douta	=	16'h	7476;
35298	:douta	=	16'h	6c35;
35299	:douta	=	16'h	9d9a;
35300	:douta	=	16'h	3aad;
35301	:douta	=	16'h	29a8;
35302	:douta	=	16'h	31ca;
35303	:douta	=	16'h	29a9;
35304	:douta	=	16'h	31ea;
35305	:douta	=	16'h	39eb;
35306	:douta	=	16'h	3a2b;
35307	:douta	=	16'h	3a0b;
35308	:douta	=	16'h	3a6c;
35309	:douta	=	16'h	3a4c;
35310	:douta	=	16'h	326d;
35311	:douta	=	16'h	3a8d;
35312	:douta	=	16'h	42cf;
35313	:douta	=	16'h	4b31;
35314	:douta	=	16'h	5bd3;
35315	:douta	=	16'h	6477;
35316	:douta	=	16'h	634f;
35317	:douta	=	16'h	51e7;
35318	:douta	=	16'h	49c7;
35319	:douta	=	16'h	3987;
35320	:douta	=	16'h	41a7;
35321	:douta	=	16'h	3987;
35322	:douta	=	16'h	41a7;
35323	:douta	=	16'h	49c7;
35324	:douta	=	16'h	49e7;
35325	:douta	=	16'h	4a08;
35326	:douta	=	16'h	49e8;
35327	:douta	=	16'h	49e8;
35328	:douta	=	16'h	e56d;
35329	:douta	=	16'h	e56c;
35330	:douta	=	16'h	dd4c;
35331	:douta	=	16'h	e54b;
35332	:douta	=	16'h	7b28;
35333	:douta	=	16'h	3104;
35334	:douta	=	16'h	4985;
35335	:douta	=	16'h	51c6;
35336	:douta	=	16'h	5a6a;
35337	:douta	=	16'h	2903;
35338	:douta	=	16'h	7391;
35339	:douta	=	16'h	8c13;
35340	:douta	=	16'h	73b0;
35341	:douta	=	16'h	62ee;
35342	:douta	=	16'h	5a6a;
35343	:douta	=	16'h	8b8e;
35344	:douta	=	16'h	9432;
35345	:douta	=	16'h	9495;
35346	:douta	=	16'h	ad99;
35347	:douta	=	16'h	29ca;
35348	:douta	=	16'h	2169;
35349	:douta	=	16'h	320b;
35350	:douta	=	16'h	322c;
35351	:douta	=	16'h	29a9;
35352	:douta	=	16'h	320b;
35353	:douta	=	16'h	3a4c;
35354	:douta	=	16'h	3a8d;
35355	:douta	=	16'h	3a4c;
35356	:douta	=	16'h	42ae;
35357	:douta	=	16'h	42ad;
35358	:douta	=	16'h	3a8d;
35359	:douta	=	16'h	4b0f;
35360	:douta	=	16'h	4aee;
35361	:douta	=	16'h	42ad;
35362	:douta	=	16'h	428d;
35363	:douta	=	16'h	2a0a;
35364	:douta	=	16'h	324b;
35365	:douta	=	16'h	322b;
35366	:douta	=	16'h	3a6b;
35367	:douta	=	16'h	3a6b;
35368	:douta	=	16'h	42ac;
35369	:douta	=	16'h	3a6b;
35370	:douta	=	16'h	42ac;
35371	:douta	=	16'h	4acd;
35372	:douta	=	16'h	4b0e;
35373	:douta	=	16'h	4aed;
35374	:douta	=	16'h	42ac;
35375	:douta	=	16'h	3a6b;
35376	:douta	=	16'h	4a8c;
35377	:douta	=	16'h	3a4a;
35378	:douta	=	16'h	428b;
35379	:douta	=	16'h	4aac;
35380	:douta	=	16'h	52ed;
35381	:douta	=	16'h	530d;
35382	:douta	=	16'h	52ed;
35383	:douta	=	16'h	530d;
35384	:douta	=	16'h	5b4e;
35385	:douta	=	16'h	532e;
35386	:douta	=	16'h	534e;
35387	:douta	=	16'h	532e;
35388	:douta	=	16'h	532e;
35389	:douta	=	16'h	5b8f;
35390	:douta	=	16'h	63b0;
35391	:douta	=	16'h	5b6f;
35392	:douta	=	16'h	5b6f;
35393	:douta	=	16'h	5b6f;
35394	:douta	=	16'h	6bd0;
35395	:douta	=	16'h	63b0;
35396	:douta	=	16'h	6390;
35397	:douta	=	16'h	6bf0;
35398	:douta	=	16'h	7411;
35399	:douta	=	16'h	536f;
35400	:douta	=	16'h	73f0;
35401	:douta	=	16'h	ee34;
35402	:douta	=	16'h	e675;
35403	:douta	=	16'h	d5b2;
35404	:douta	=	16'h	ee96;
35405	:douta	=	16'h	ddf3;
35406	:douta	=	16'h	e675;
35407	:douta	=	16'h	93f0;
35408	:douta	=	16'h	c512;
35409	:douta	=	16'h	c533;
35410	:douta	=	16'h	acd2;
35411	:douta	=	16'h	8432;
35412	:douta	=	16'h	b4f2;
35413	:douta	=	16'h	a492;
35414	:douta	=	16'h	9453;
35415	:douta	=	16'h	8411;
35416	:douta	=	16'h	738f;
35417	:douta	=	16'h	736f;
35418	:douta	=	16'h	62ec;
35419	:douta	=	16'h	732d;
35420	:douta	=	16'h	6b2c;
35421	:douta	=	16'h	6aec;
35422	:douta	=	16'h	5aaa;
35423	:douta	=	16'h	5a8b;
35424	:douta	=	16'h	836c;
35425	:douta	=	16'h	a40c;
35426	:douta	=	16'h	ee96;
35427	:douta	=	16'h	de56;
35428	:douta	=	16'h	de15;
35429	:douta	=	16'h	7413;
35430	:douta	=	16'h	7c13;
35431	:douta	=	16'h	bd54;
35432	:douta	=	16'h	9cd4;
35433	:douta	=	16'h	94d5;
35434	:douta	=	16'h	9495;
35435	:douta	=	16'h	94d5;
35436	:douta	=	16'h	94b5;
35437	:douta	=	16'h	8cb4;
35438	:douta	=	16'h	7bf2;
35439	:douta	=	16'h	7bf1;
35440	:douta	=	16'h	7bb0;
35441	:douta	=	16'h	734f;
35442	:douta	=	16'h	6b0d;
35443	:douta	=	16'h	6b2d;
35444	:douta	=	16'h	734f;
35445	:douta	=	16'h	7b8f;
35446	:douta	=	16'h	528c;
35447	:douta	=	16'h	4a4c;
35448	:douta	=	16'h	b46f;
35449	:douta	=	16'h	c530;
35450	:douta	=	16'h	cd51;
35451	:douta	=	16'h	a494;
35452	:douta	=	16'h	a4b4;
35453	:douta	=	16'h	a4b4;
35454	:douta	=	16'h	8453;
35455	:douta	=	16'h	6bb1;
35456	:douta	=	16'h	9c93;
35457	:douta	=	16'h	8433;
35458	:douta	=	16'h	7390;
35459	:douta	=	16'h	62ee;
35460	:douta	=	16'h	632f;
35461	:douta	=	16'h	632f;
35462	:douta	=	16'h	4aad;
35463	:douta	=	16'h	6b2e;
35464	:douta	=	16'h	7b4e;
35465	:douta	=	16'h	6acc;
35466	:douta	=	16'h	5a6b;
35467	:douta	=	16'h	526b;
35468	:douta	=	16'h	5a8b;
35469	:douta	=	16'h	9452;
35470	:douta	=	16'h	9c94;
35471	:douta	=	16'h	73d0;
35472	:douta	=	16'h	7b6f;
35473	:douta	=	16'h	7b8e;
35474	:douta	=	16'h	734d;
35475	:douta	=	16'h	734d;
35476	:douta	=	16'h	732d;
35477	:douta	=	16'h	6aec;
35478	:douta	=	16'h	4a8b;
35479	:douta	=	16'h	52ac;
35480	:douta	=	16'h	5aed;
35481	:douta	=	16'h	632e;
35482	:douta	=	16'h	7baf;
35483	:douta	=	16'h	732e;
35484	:douta	=	16'h	4a6c;
35485	:douta	=	16'h	62cd;
35486	:douta	=	16'h	bd32;
35487	:douta	=	16'h	ee35;
35488	:douta	=	16'h	9493;
35489	:douta	=	16'h	8413;
35490	:douta	=	16'h	8c32;
35491	:douta	=	16'h	a4d4;
35492	:douta	=	16'h	9c94;
35493	:douta	=	16'h	83f1;
35494	:douta	=	16'h	6b6f;
35495	:douta	=	16'h	6b4f;
35496	:douta	=	16'h	7bd1;
35497	:douta	=	16'h	7bb0;
35498	:douta	=	16'h	5aee;
35499	:douta	=	16'h	52cd;
35500	:douta	=	16'h	632e;
35501	:douta	=	16'h	738f;
35502	:douta	=	16'h	7bb0;
35503	:douta	=	16'h	734e;
35504	:douta	=	16'h	632e;
35505	:douta	=	16'h	424c;
35506	:douta	=	16'h	7b8f;
35507	:douta	=	16'h	8c10;
35508	:douta	=	16'h	8bef;
35509	:douta	=	16'h	b4d1;
35510	:douta	=	16'h	d616;
35511	:douta	=	16'h	e678;
35512	:douta	=	16'h	de36;
35513	:douta	=	16'h	cdb6;
35514	:douta	=	16'h	cdb5;
35515	:douta	=	16'h	bd74;
35516	:douta	=	16'h	94d5;
35517	:douta	=	16'h	94b5;
35518	:douta	=	16'h	8454;
35519	:douta	=	16'h	8454;
35520	:douta	=	16'h	73d1;
35521	:douta	=	16'h	73b1;
35522	:douta	=	16'h	6b91;
35523	:douta	=	16'h	6371;
35524	:douta	=	16'h	6371;
35525	:douta	=	16'h	6391;
35526	:douta	=	16'h	5330;
35527	:douta	=	16'h	4acf;
35528	:douta	=	16'h	3a4d;
35529	:douta	=	16'h	3a6d;
35530	:douta	=	16'h	3a6e;
35531	:douta	=	16'h	21aa;
35532	:douta	=	16'h	52ed;
35533	:douta	=	16'h	426d;
35534	:douta	=	16'h	2148;
35535	:douta	=	16'h	428c;
35536	:douta	=	16'h	10e4;
35537	:douta	=	16'h	1926;
35538	:douta	=	16'h	10c5;
35539	:douta	=	16'h	10c4;
35540	:douta	=	16'h	18e5;
35541	:douta	=	16'h	2167;
35542	:douta	=	16'h	1927;
35543	:douta	=	16'h	7413;
35544	:douta	=	16'h	9d79;
35545	:douta	=	16'h	94f6;
35546	:douta	=	16'h	6bd4;
35547	:douta	=	16'h	7414;
35548	:douta	=	16'h	7434;
35549	:douta	=	16'h	8497;
35550	:douta	=	16'h	63f5;
35551	:douta	=	16'h	8d18;
35552	:douta	=	16'h	8cf8;
35553	:douta	=	16'h	8cf7;
35554	:douta	=	16'h	a5db;
35555	:douta	=	16'h	4b10;
35556	:douta	=	16'h	2126;
35557	:douta	=	16'h	29a9;
35558	:douta	=	16'h	3a2b;
35559	:douta	=	16'h	3a2b;
35560	:douta	=	16'h	424b;
35561	:douta	=	16'h	42ad;
35562	:douta	=	16'h	426c;
35563	:douta	=	16'h	5bb2;
35564	:douta	=	16'h	63d3;
35565	:douta	=	16'h	5391;
35566	:douta	=	16'h	5bf4;
35567	:douta	=	16'h	6435;
35568	:douta	=	16'h	5bb3;
35569	:douta	=	16'h	5bd3;
35570	:douta	=	16'h	5c36;
35571	:douta	=	16'h	42cf;
35572	:douta	=	16'h	5b92;
35573	:douta	=	16'h	6a88;
35574	:douta	=	16'h	49c6;
35575	:douta	=	16'h	3986;
35576	:douta	=	16'h	49c7;
35577	:douta	=	16'h	3966;
35578	:douta	=	16'h	41c7;
35579	:douta	=	16'h	49e7;
35580	:douta	=	16'h	49e7;
35581	:douta	=	16'h	49e7;
35582	:douta	=	16'h	49e8;
35583	:douta	=	16'h	49c7;
35584	:douta	=	16'h	e58d;
35585	:douta	=	16'h	e56c;
35586	:douta	=	16'h	e56c;
35587	:douta	=	16'h	dd4b;
35588	:douta	=	16'h	c509;
35589	:douta	=	16'h	49c5;
35590	:douta	=	16'h	51c5;
35591	:douta	=	16'h	5164;
35592	:douta	=	16'h	83ad;
35593	:douta	=	16'h	9432;
35594	:douta	=	16'h	bd98;
35595	:douta	=	16'h	83f2;
35596	:douta	=	16'h	7bf1;
35597	:douta	=	16'h	734f;
35598	:douta	=	16'h	8b4d;
35599	:douta	=	16'h	a410;
35600	:douta	=	16'h	ad57;
35601	:douta	=	16'h	ad78;
35602	:douta	=	16'h	9d17;
35603	:douta	=	16'h	21ca;
35604	:douta	=	16'h	29eb;
35605	:douta	=	16'h	322c;
35606	:douta	=	16'h	320c;
35607	:douta	=	16'h	2189;
35608	:douta	=	16'h	320b;
35609	:douta	=	16'h	3a4c;
35610	:douta	=	16'h	42ae;
35611	:douta	=	16'h	3a6d;
35612	:douta	=	16'h	3a8d;
35613	:douta	=	16'h	3a6c;
35614	:douta	=	16'h	3a6d;
35615	:douta	=	16'h	42ae;
35616	:douta	=	16'h	428d;
35617	:douta	=	16'h	4ace;
35618	:douta	=	16'h	42ad;
35619	:douta	=	16'h	324b;
35620	:douta	=	16'h	322a;
35621	:douta	=	16'h	322b;
35622	:douta	=	16'h	3a4b;
35623	:douta	=	16'h	3a6b;
35624	:douta	=	16'h	3a8c;
35625	:douta	=	16'h	3a6b;
35626	:douta	=	16'h	428c;
35627	:douta	=	16'h	3a6b;
35628	:douta	=	16'h	3a8c;
35629	:douta	=	16'h	42cd;
35630	:douta	=	16'h	4b0e;
35631	:douta	=	16'h	4b0e;
35632	:douta	=	16'h	3a6b;
35633	:douta	=	16'h	31e9;
35634	:douta	=	16'h	322a;
35635	:douta	=	16'h	4a8c;
35636	:douta	=	16'h	4aac;
35637	:douta	=	16'h	424b;
35638	:douta	=	16'h	530d;
35639	:douta	=	16'h	530e;
35640	:douta	=	16'h	5b4e;
35641	:douta	=	16'h	5b4f;
35642	:douta	=	16'h	5b6f;
35643	:douta	=	16'h	5b6f;
35644	:douta	=	16'h	534e;
35645	:douta	=	16'h	42ac;
35646	:douta	=	16'h	532e;
35647	:douta	=	16'h	5b6f;
35648	:douta	=	16'h	5b4f;
35649	:douta	=	16'h	5b8f;
35650	:douta	=	16'h	6390;
35651	:douta	=	16'h	6390;
35652	:douta	=	16'h	63b0;
35653	:douta	=	16'h	63d1;
35654	:douta	=	16'h	6c11;
35655	:douta	=	16'h	5b70;
35656	:douta	=	16'h	63af;
35657	:douta	=	16'h	4b2e;
35658	:douta	=	16'h	cd71;
35659	:douta	=	16'h	c510;
35660	:douta	=	16'h	d5b4;
35661	:douta	=	16'h	bcf2;
35662	:douta	=	16'h	bd33;
35663	:douta	=	16'h	acb2;
35664	:douta	=	16'h	9c93;
35665	:douta	=	16'h	c533;
35666	:douta	=	16'h	acd2;
35667	:douta	=	16'h	8432;
35668	:douta	=	16'h	9c93;
35669	:douta	=	16'h	9473;
35670	:douta	=	16'h	7bf1;
35671	:douta	=	16'h	83d0;
35672	:douta	=	16'h	7baf;
35673	:douta	=	16'h	7b90;
35674	:douta	=	16'h	6b2e;
35675	:douta	=	16'h	6b0d;
35676	:douta	=	16'h	6b0c;
35677	:douta	=	16'h	62cc;
35678	:douta	=	16'h	62ed;
35679	:douta	=	16'h	8b29;
35680	:douta	=	16'h	d5f3;
35681	:douta	=	16'h	de55;
35682	:douta	=	16'h	e655;
35683	:douta	=	16'h	de35;
35684	:douta	=	16'h	bd75;
35685	:douta	=	16'h	9d16;
35686	:douta	=	16'h	84b5;
35687	:douta	=	16'h	8c74;
35688	:douta	=	16'h	b556;
35689	:douta	=	16'h	94b5;
35690	:douta	=	16'h	8454;
35691	:douta	=	16'h	8c94;
35692	:douta	=	16'h	8c94;
35693	:douta	=	16'h	8c53;
35694	:douta	=	16'h	7370;
35695	:douta	=	16'h	734e;
35696	:douta	=	16'h	734e;
35697	:douta	=	16'h	734f;
35698	:douta	=	16'h	7b6f;
35699	:douta	=	16'h	8390;
35700	:douta	=	16'h	52ac;
35701	:douta	=	16'h	730d;
35702	:douta	=	16'h	ddb2;
35703	:douta	=	16'h	d5b3;
35704	:douta	=	16'h	d593;
35705	:douta	=	16'h	bd75;
35706	:douta	=	16'h	b533;
35707	:douta	=	16'h	bd55;
35708	:douta	=	16'h	a4b4;
35709	:douta	=	16'h	ad35;
35710	:douta	=	16'h	9495;
35711	:douta	=	16'h	8434;
35712	:douta	=	16'h	6371;
35713	:douta	=	16'h	6bb1;
35714	:douta	=	16'h	7bb1;
35715	:douta	=	16'h	736f;
35716	:douta	=	16'h	62cd;
35717	:douta	=	16'h	39eb;
35718	:douta	=	16'h	31ca;
35719	:douta	=	16'h	420a;
35720	:douta	=	16'h	31a8;
35721	:douta	=	16'h	31a8;
35722	:douta	=	16'h	526c;
35723	:douta	=	16'h	7bb0;
35724	:douta	=	16'h	a4b5;
35725	:douta	=	16'h	7bd1;
35726	:douta	=	16'h	7370;
35727	:douta	=	16'h	732e;
35728	:douta	=	16'h	62ed;
35729	:douta	=	16'h	5a8b;
35730	:douta	=	16'h	732d;
35731	:douta	=	16'h	732d;
35732	:douta	=	16'h	734d;
35733	:douta	=	16'h	730c;
35734	:douta	=	16'h	422a;
35735	:douta	=	16'h	31c9;
35736	:douta	=	16'h	31a8;
35737	:douta	=	16'h	39c9;
35738	:douta	=	16'h	420c;
35739	:douta	=	16'h	cdb4;
35740	:douta	=	16'h	d595;
35741	:douta	=	16'h	b514;
35742	:douta	=	16'h	a4b4;
35743	:douta	=	16'h	9cb5;
35744	:douta	=	16'h	9474;
35745	:douta	=	16'h	9494;
35746	:douta	=	16'h	8c74;
35747	:douta	=	16'h	7bd1;
35748	:douta	=	16'h	7b8f;
35749	:douta	=	16'h	734e;
35750	:douta	=	16'h	734e;
35751	:douta	=	16'h	6b0e;
35752	:douta	=	16'h	5acc;
35753	:douta	=	16'h	62ed;
35754	:douta	=	16'h	630d;
35755	:douta	=	16'h	5aed;
35756	:douta	=	16'h	422b;
35757	:douta	=	16'h	31ca;
35758	:douta	=	16'h	3a2b;
35759	:douta	=	16'h	62ac;
35760	:douta	=	16'h	836d;
35761	:douta	=	16'h	ee75;
35762	:douta	=	16'h	eeb7;
35763	:douta	=	16'h	e697;
35764	:douta	=	16'h	de57;
35765	:douta	=	16'h	cdf7;
35766	:douta	=	16'h	cdf6;
35767	:douta	=	16'h	c5b6;
35768	:douta	=	16'h	bd76;
35769	:douta	=	16'h	ad15;
35770	:douta	=	16'h	ad15;
35771	:douta	=	16'h	ad15;
35772	:douta	=	16'h	9c94;
35773	:douta	=	16'h	8452;
35774	:douta	=	16'h	7bd1;
35775	:douta	=	16'h	6b91;
35776	:douta	=	16'h	6b91;
35777	:douta	=	16'h	6b90;
35778	:douta	=	16'h	6b90;
35779	:douta	=	16'h	6b91;
35780	:douta	=	16'h	6b91;
35781	:douta	=	16'h	5b30;
35782	:douta	=	16'h	52ef;
35783	:douta	=	16'h	4ace;
35784	:douta	=	16'h	4aae;
35785	:douta	=	16'h	3a2c;
35786	:douta	=	16'h	62eb;
35787	:douta	=	16'h	c574;
35788	:douta	=	16'h	6b92;
35789	:douta	=	16'h	21aa;
35790	:douta	=	16'h	2168;
35791	:douta	=	16'h	18c5;
35792	:douta	=	16'h	5b50;
35793	:douta	=	16'h	31c9;
35794	:douta	=	16'h	10a4;
35795	:douta	=	16'h	10c4;
35796	:douta	=	16'h	18e5;
35797	:douta	=	16'h	18e5;
35798	:douta	=	16'h	10e5;
35799	:douta	=	16'h	0083;
35800	:douta	=	16'h	63b2;
35801	:douta	=	16'h	63b2;
35802	:douta	=	16'h	8cd7;
35803	:douta	=	16'h	9d58;
35804	:douta	=	16'h	6c15;
35805	:douta	=	16'h	84b5;
35806	:douta	=	16'h	6c16;
35807	:douta	=	16'h	9d58;
35808	:douta	=	16'h	a599;
35809	:douta	=	16'h	7c76;
35810	:douta	=	16'h	4b10;
35811	:douta	=	16'h	5330;
35812	:douta	=	16'h	63f2;
35813	:douta	=	16'h	6414;
35814	:douta	=	16'h	6c34;
35815	:douta	=	16'h	6c14;
35816	:douta	=	16'h	7cf7;
35817	:douta	=	16'h	6c77;
35818	:douta	=	16'h	855a;
35819	:douta	=	16'h	6bf3;
35820	:douta	=	16'h	5b50;
35821	:douta	=	16'h	630c;
35822	:douta	=	16'h	5a47;
35823	:douta	=	16'h	6247;
35824	:douta	=	16'h	6a25;
35825	:douta	=	16'h	6a46;
35826	:douta	=	16'h	69e4;
35827	:douta	=	16'h	61e4;
35828	:douta	=	16'h	61e4;
35829	:douta	=	16'h	59e5;
35830	:douta	=	16'h	6a47;
35831	:douta	=	16'h	5a28;
35832	:douta	=	16'h	41a7;
35833	:douta	=	16'h	49e8;
35834	:douta	=	16'h	49e7;
35835	:douta	=	16'h	41a7;
35836	:douta	=	16'h	49c7;
35837	:douta	=	16'h	49c7;
35838	:douta	=	16'h	49c7;
35839	:douta	=	16'h	41c7;
35840	:douta	=	16'h	e58d;
35841	:douta	=	16'h	e58d;
35842	:douta	=	16'h	e56d;
35843	:douta	=	16'h	e56c;
35844	:douta	=	16'h	e58c;
35845	:douta	=	16'h	6a86;
35846	:douta	=	16'h	59e6;
35847	:douta	=	16'h	51c5;
35848	:douta	=	16'h	8bae;
35849	:douta	=	16'h	9cb5;
35850	:douta	=	16'h	b516;
35851	:douta	=	16'h	8c32;
35852	:douta	=	16'h	9452;
35853	:douta	=	16'h	6b0d;
35854	:douta	=	16'h	a40f;
35855	:douta	=	16'h	ac51;
35856	:douta	=	16'h	b557;
35857	:douta	=	16'h	b577;
35858	:douta	=	16'h	9d17;
35859	:douta	=	16'h	2188;
35860	:douta	=	16'h	29ca;
35861	:douta	=	16'h	322c;
35862	:douta	=	16'h	322c;
35863	:douta	=	16'h	2188;
35864	:douta	=	16'h	29aa;
35865	:douta	=	16'h	29eb;
35866	:douta	=	16'h	322c;
35867	:douta	=	16'h	3a4c;
35868	:douta	=	16'h	42ae;
35869	:douta	=	16'h	3a6d;
35870	:douta	=	16'h	3a6d;
35871	:douta	=	16'h	3a8d;
35872	:douta	=	16'h	3a8d;
35873	:douta	=	16'h	4ace;
35874	:douta	=	16'h	428d;
35875	:douta	=	16'h	322a;
35876	:douta	=	16'h	322b;
35877	:douta	=	16'h	2a0a;
35878	:douta	=	16'h	322a;
35879	:douta	=	16'h	324b;
35880	:douta	=	16'h	3a6b;
35881	:douta	=	16'h	3a8c;
35882	:douta	=	16'h	3a6c;
35883	:douta	=	16'h	3a6c;
35884	:douta	=	16'h	428c;
35885	:douta	=	16'h	42ad;
35886	:douta	=	16'h	4b0e;
35887	:douta	=	16'h	4b2e;
35888	:douta	=	16'h	530e;
35889	:douta	=	16'h	320a;
35890	:douta	=	16'h	3a2a;
35891	:douta	=	16'h	322a;
35892	:douta	=	16'h	3a4a;
35893	:douta	=	16'h	426b;
35894	:douta	=	16'h	530d;
35895	:douta	=	16'h	4acd;
35896	:douta	=	16'h	5b6f;
35897	:douta	=	16'h	534e;
35898	:douta	=	16'h	63b0;
35899	:douta	=	16'h	534e;
35900	:douta	=	16'h	4b0d;
35901	:douta	=	16'h	4aed;
35902	:douta	=	16'h	5b4f;
35903	:douta	=	16'h	5b4f;
35904	:douta	=	16'h	5b6f;
35905	:douta	=	16'h	6390;
35906	:douta	=	16'h	6390;
35907	:douta	=	16'h	6390;
35908	:douta	=	16'h	6390;
35909	:douta	=	16'h	6c11;
35910	:douta	=	16'h	63b1;
35911	:douta	=	16'h	6390;
35912	:douta	=	16'h	638f;
35913	:douta	=	16'h	63b0;
35914	:douta	=	16'h	6b6f;
35915	:douta	=	16'h	7bce;
35916	:douta	=	16'h	bcf1;
35917	:douta	=	16'h	b4d2;
35918	:douta	=	16'h	b4f2;
35919	:douta	=	16'h	9c51;
35920	:douta	=	16'h	a472;
35921	:douta	=	16'h	acb3;
35922	:douta	=	16'h	acd3;
35923	:douta	=	16'h	8433;
35924	:douta	=	16'h	8412;
35925	:douta	=	16'h	8c32;
35926	:douta	=	16'h	83f0;
35927	:douta	=	16'h	7bd0;
35928	:douta	=	16'h	7baf;
35929	:douta	=	16'h	734e;
35930	:douta	=	16'h	7b6f;
35931	:douta	=	16'h	6b0c;
35932	:douta	=	16'h	6b0d;
35933	:douta	=	16'h	5a6b;
35934	:douta	=	16'h	8bad;
35935	:douta	=	16'h	d591;
35936	:douta	=	16'h	d5d4;
35937	:douta	=	16'h	eeb7;
35938	:douta	=	16'h	de15;
35939	:douta	=	16'h	cdb4;
35940	:douta	=	16'h	ad15;
35941	:douta	=	16'h	9d15;
35942	:douta	=	16'h	94d6;
35943	:douta	=	16'h	6371;
35944	:douta	=	16'h	9494;
35945	:douta	=	16'h	94b4;
35946	:douta	=	16'h	73d1;
35947	:douta	=	16'h	73d0;
35948	:douta	=	16'h	8453;
35949	:douta	=	16'h	8453;
35950	:douta	=	16'h	7bb0;
35951	:douta	=	16'h	736e;
35952	:douta	=	16'h	736e;
35953	:douta	=	16'h	736f;
35954	:douta	=	16'h	736e;
35955	:douta	=	16'h	62ed;
35956	:douta	=	16'h	8bce;
35957	:douta	=	16'h	bcd0;
35958	:douta	=	16'h	ee55;
35959	:douta	=	16'h	cdb4;
35960	:douta	=	16'h	acf3;
35961	:douta	=	16'h	8c53;
35962	:douta	=	16'h	6bb2;
35963	:douta	=	16'h	8413;
35964	:douta	=	16'h	8c53;
35965	:douta	=	16'h	8c74;
35966	:douta	=	16'h	8433;
35967	:douta	=	16'h	7bf3;
35968	:douta	=	16'h	6b91;
35969	:douta	=	16'h	634f;
35970	:douta	=	16'h	6b6f;
35971	:douta	=	16'h	7391;
35972	:douta	=	16'h	7391;
35973	:douta	=	16'h	62cc;
35974	:douta	=	16'h	5a8b;
35975	:douta	=	16'h	4a2a;
35976	:douta	=	16'h	5a8b;
35977	:douta	=	16'h	734f;
35978	:douta	=	16'h	6b71;
35979	:douta	=	16'h	6370;
35980	:douta	=	16'h	9432;
35981	:douta	=	16'h	7bb0;
35982	:douta	=	16'h	7b90;
35983	:douta	=	16'h	6aec;
35984	:douta	=	16'h	62cc;
35985	:douta	=	16'h	524a;
35986	:douta	=	16'h	526b;
35987	:douta	=	16'h	5a8b;
35988	:douta	=	16'h	732c;
35989	:douta	=	16'h	7b2d;
35990	:douta	=	16'h	6acb;
35991	:douta	=	16'h	31c9;
35992	:douta	=	16'h	422a;
35993	:douta	=	16'h	6370;
35994	:douta	=	16'h	8413;
35995	:douta	=	16'h	acd3;
35996	:douta	=	16'h	acf5;
35997	:douta	=	16'h	acf5;
35998	:douta	=	16'h	9cb5;
35999	:douta	=	16'h	a4d5;
36000	:douta	=	16'h	8c73;
36001	:douta	=	16'h	8412;
36002	:douta	=	16'h	8433;
36003	:douta	=	16'h	8432;
36004	:douta	=	16'h	7bf2;
36005	:douta	=	16'h	736f;
36006	:douta	=	16'h	6b0d;
36007	:douta	=	16'h	6aed;
36008	:douta	=	16'h	62cd;
36009	:douta	=	16'h	5a8c;
36010	:douta	=	16'h	5acd;
36011	:douta	=	16'h	5aee;
36012	:douta	=	16'h	4a6c;
36013	:douta	=	16'h	6b0d;
36014	:douta	=	16'h	838e;
36015	:douta	=	16'h	93ee;
36016	:douta	=	16'h	ac6f;
36017	:douta	=	16'h	b512;
36018	:douta	=	16'h	de36;
36019	:douta	=	16'h	d617;
36020	:douta	=	16'h	bd96;
36021	:douta	=	16'h	bd76;
36022	:douta	=	16'h	b536;
36023	:douta	=	16'h	b556;
36024	:douta	=	16'h	bd76;
36025	:douta	=	16'h	ad36;
36026	:douta	=	16'h	ad15;
36027	:douta	=	16'h	9494;
36028	:douta	=	16'h	8432;
36029	:douta	=	16'h	7bf2;
36030	:douta	=	16'h	6b90;
36031	:douta	=	16'h	6b90;
36032	:douta	=	16'h	6b90;
36033	:douta	=	16'h	73d1;
36034	:douta	=	16'h	73f2;
36035	:douta	=	16'h	6b91;
36036	:douta	=	16'h	6350;
36037	:douta	=	16'h	5b50;
36038	:douta	=	16'h	52ce;
36039	:douta	=	16'h	52cf;
36040	:douta	=	16'h	31c9;
36041	:douta	=	16'h	4a09;
36042	:douta	=	16'h	e634;
36043	:douta	=	16'h	8c52;
36044	:douta	=	16'h	4acf;
36045	:douta	=	16'h	1968;
36046	:douta	=	16'h	39ea;
36047	:douta	=	16'h	1906;
36048	:douta	=	16'h	2987;
36049	:douta	=	16'h	52ce;
36050	:douta	=	16'h	0863;
36051	:douta	=	16'h	18c4;
36052	:douta	=	16'h	18e4;
36053	:douta	=	16'h	1906;
36054	:douta	=	16'h	10e4;
36055	:douta	=	16'h	1947;
36056	:douta	=	16'h	42ce;
36057	:douta	=	16'h	7c55;
36058	:douta	=	16'h	84b6;
36059	:douta	=	16'h	7c96;
36060	:douta	=	16'h	84d7;
36061	:douta	=	16'h	a598;
36062	:douta	=	16'h	84b7;
36063	:douta	=	16'h	9518;
36064	:douta	=	16'h	84b8;
36065	:douta	=	16'h	4310;
36066	:douta	=	16'h	42ee;
36067	:douta	=	16'h	7cf8;
36068	:douta	=	16'h	7d19;
36069	:douta	=	16'h	8539;
36070	:douta	=	16'h	7413;
36071	:douta	=	16'h	6390;
36072	:douta	=	16'h	73d0;
36073	:douta	=	16'h	72ea;
36074	:douta	=	16'h	6a47;
36075	:douta	=	16'h	6a25;
36076	:douta	=	16'h	7246;
36077	:douta	=	16'h	7204;
36078	:douta	=	16'h	7224;
36079	:douta	=	16'h	6a25;
36080	:douta	=	16'h	6a25;
36081	:douta	=	16'h	6a05;
36082	:douta	=	16'h	6a26;
36083	:douta	=	16'h	6205;
36084	:douta	=	16'h	6205;
36085	:douta	=	16'h	59c5;
36086	:douta	=	16'h	59e5;
36087	:douta	=	16'h	728a;
36088	:douta	=	16'h	41c7;
36089	:douta	=	16'h	49e8;
36090	:douta	=	16'h	49e7;
36091	:douta	=	16'h	49e7;
36092	:douta	=	16'h	49e8;
36093	:douta	=	16'h	49e8;
36094	:douta	=	16'h	49e8;
36095	:douta	=	16'h	49e7;
36096	:douta	=	16'h	e58c;
36097	:douta	=	16'h	e58e;
36098	:douta	=	16'h	e56d;
36099	:douta	=	16'h	e56c;
36100	:douta	=	16'h	f60d;
36101	:douta	=	16'h	ac48;
36102	:douta	=	16'h	6206;
36103	:douta	=	16'h	6226;
36104	:douta	=	16'h	49c5;
36105	:douta	=	16'h	cdb7;
36106	:douta	=	16'h	acd4;
36107	:douta	=	16'h	9c53;
36108	:douta	=	16'h	9412;
36109	:douta	=	16'h	83b0;
36110	:douta	=	16'h	c490;
36111	:douta	=	16'h	cd96;
36112	:douta	=	16'h	bd97;
36113	:douta	=	16'h	b577;
36114	:douta	=	16'h	7c75;
36115	:douta	=	16'h	1906;
36116	:douta	=	16'h	1926;
36117	:douta	=	16'h	08a4;
36118	:douta	=	16'h	1947;
36119	:douta	=	16'h	21a9;
36120	:douta	=	16'h	2168;
36121	:douta	=	16'h	2188;
36122	:douta	=	16'h	21a9;
36123	:douta	=	16'h	31eb;
36124	:douta	=	16'h	324c;
36125	:douta	=	16'h	3a6d;
36126	:douta	=	16'h	3a6d;
36127	:douta	=	16'h	3a6c;
36128	:douta	=	16'h	324c;
36129	:douta	=	16'h	29eb;
36130	:douta	=	16'h	3a6c;
36131	:douta	=	16'h	3a4b;
36132	:douta	=	16'h	3a4b;
36133	:douta	=	16'h	3a6c;
36134	:douta	=	16'h	3a6c;
36135	:douta	=	16'h	322b;
36136	:douta	=	16'h	322b;
36137	:douta	=	16'h	322b;
36138	:douta	=	16'h	3a8c;
36139	:douta	=	16'h	324b;
36140	:douta	=	16'h	3a4b;
36141	:douta	=	16'h	428c;
36142	:douta	=	16'h	428c;
36143	:douta	=	16'h	42ac;
36144	:douta	=	16'h	42ac;
36145	:douta	=	16'h	4aed;
36146	:douta	=	16'h	4acd;
36147	:douta	=	16'h	52ee;
36148	:douta	=	16'h	4acd;
36149	:douta	=	16'h	4acd;
36150	:douta	=	16'h	42ac;
36151	:douta	=	16'h	42ac;
36152	:douta	=	16'h	3a6b;
36153	:douta	=	16'h	428c;
36154	:douta	=	16'h	534f;
36155	:douta	=	16'h	532e;
36156	:douta	=	16'h	534f;
36157	:douta	=	16'h	5b6f;
36158	:douta	=	16'h	534e;
36159	:douta	=	16'h	534f;
36160	:douta	=	16'h	5b4f;
36161	:douta	=	16'h	5b6f;
36162	:douta	=	16'h	6390;
36163	:douta	=	16'h	5b6f;
36164	:douta	=	16'h	5b6f;
36165	:douta	=	16'h	63b0;
36166	:douta	=	16'h	63b0;
36167	:douta	=	16'h	5b8f;
36168	:douta	=	16'h	5b8f;
36169	:douta	=	16'h	636f;
36170	:douta	=	16'h	63af;
36171	:douta	=	16'h	6bb0;
36172	:douta	=	16'h	5b4f;
36173	:douta	=	16'h	736f;
36174	:douta	=	16'h	940f;
36175	:douta	=	16'h	9c50;
36176	:douta	=	16'h	9431;
36177	:douta	=	16'h	9430;
36178	:douta	=	16'h	8bf0;
36179	:douta	=	16'h	7bcf;
36180	:douta	=	16'h	7baf;
36181	:douta	=	16'h	7b8f;
36182	:douta	=	16'h	83f1;
36183	:douta	=	16'h	7bb0;
36184	:douta	=	16'h	738f;
36185	:douta	=	16'h	732d;
36186	:douta	=	16'h	6b0d;
36187	:douta	=	16'h	528c;
36188	:douta	=	16'h	5a4a;
36189	:douta	=	16'h	f694;
36190	:douta	=	16'h	d593;
36191	:douta	=	16'h	ee97;
36192	:douta	=	16'h	cdb4;
36193	:douta	=	16'h	e696;
36194	:douta	=	16'h	b555;
36195	:douta	=	16'h	ad36;
36196	:douta	=	16'h	9cf5;
36197	:douta	=	16'h	9cf6;
36198	:douta	=	16'h	94f6;
36199	:douta	=	16'h	7c13;
36200	:douta	=	16'h	532f;
36201	:douta	=	16'h	9cd4;
36202	:douta	=	16'h	8c53;
36203	:douta	=	16'h	7c11;
36204	:douta	=	16'h	6b70;
36205	:douta	=	16'h	632f;
36206	:douta	=	16'h	632f;
36207	:douta	=	16'h	630d;
36208	:douta	=	16'h	6b2e;
36209	:douta	=	16'h	5ace;
36210	:douta	=	16'h	528d;
36211	:douta	=	16'h	bc8f;
36212	:douta	=	16'h	cd52;
36213	:douta	=	16'h	ddd4;
36214	:douta	=	16'h	d5d3;
36215	:douta	=	16'h	d5d4;
36216	:douta	=	16'h	acf3;
36217	:douta	=	16'h	94b4;
36218	:douta	=	16'h	9cd5;
36219	:douta	=	16'h	73f2;
36220	:douta	=	16'h	6371;
36221	:douta	=	16'h	52ae;
36222	:douta	=	16'h	736e;
36223	:douta	=	16'h	83ae;
36224	:douta	=	16'h	732d;
36225	:douta	=	16'h	732e;
36226	:douta	=	16'h	6b0c;
36227	:douta	=	16'h	6b0c;
36228	:douta	=	16'h	730c;
36229	:douta	=	16'h	5a6a;
36230	:douta	=	16'h	62cc;
36231	:douta	=	16'h	8bf1;
36232	:douta	=	16'h	a4b4;
36233	:douta	=	16'h	9473;
36234	:douta	=	16'h	634f;
36235	:douta	=	16'h	632f;
36236	:douta	=	16'h	632f;
36237	:douta	=	16'h	62ac;
36238	:douta	=	16'h	734d;
36239	:douta	=	16'h	6acb;
36240	:douta	=	16'h	62ab;
36241	:douta	=	16'h	62cb;
36242	:douta	=	16'h	62cb;
36243	:douta	=	16'h	5a8a;
36244	:douta	=	16'h	41e9;
36245	:douta	=	16'h	3987;
36246	:douta	=	16'h	83d0;
36247	:douta	=	16'h	e5f5;
36248	:douta	=	16'h	ddb3;
36249	:douta	=	16'h	8c55;
36250	:douta	=	16'h	73d3;
36251	:douta	=	16'h	9454;
36252	:douta	=	16'h	9c93;
36253	:douta	=	16'h	9473;
36254	:douta	=	16'h	8c93;
36255	:douta	=	16'h	7bf2;
36256	:douta	=	16'h	83f2;
36257	:douta	=	16'h	8433;
36258	:douta	=	16'h	83f2;
36259	:douta	=	16'h	736f;
36260	:douta	=	16'h	734f;
36261	:douta	=	16'h	6b0d;
36262	:douta	=	16'h	7b6f;
36263	:douta	=	16'h	734f;
36264	:douta	=	16'h	52ad;
36265	:douta	=	16'h	52ad;
36266	:douta	=	16'h	8c0f;
36267	:douta	=	16'h	bd52;
36268	:douta	=	16'h	ee75;
36269	:douta	=	16'h	ee96;
36270	:douta	=	16'h	e676;
36271	:douta	=	16'h	de36;
36272	:douta	=	16'h	e656;
36273	:douta	=	16'h	bd53;
36274	:douta	=	16'h	a4d3;
36275	:douta	=	16'h	ad14;
36276	:douta	=	16'h	b556;
36277	:douta	=	16'h	b556;
36278	:douta	=	16'h	ad36;
36279	:douta	=	16'h	9494;
36280	:douta	=	16'h	94b4;
36281	:douta	=	16'h	94b4;
36282	:douta	=	16'h	94b4;
36283	:douta	=	16'h	8c73;
36284	:douta	=	16'h	8c53;
36285	:douta	=	16'h	8433;
36286	:douta	=	16'h	8432;
36287	:douta	=	16'h	8412;
36288	:douta	=	16'h	7bd1;
36289	:douta	=	16'h	6b70;
36290	:douta	=	16'h	634f;
36291	:douta	=	16'h	632f;
36292	:douta	=	16'h	5b2f;
36293	:douta	=	16'h	4ace;
36294	:douta	=	16'h	4a2a;
36295	:douta	=	16'h	7b2c;
36296	:douta	=	16'h	e613;
36297	:douta	=	16'h	e635;
36298	:douta	=	16'h	d5b2;
36299	:douta	=	16'h	6bb1;
36300	:douta	=	16'h	42ae;
36301	:douta	=	16'h	52cd;
36302	:douta	=	16'h	636e;
36303	:douta	=	16'h	320b;
36304	:douta	=	16'h	29c9;
36305	:douta	=	16'h	1905;
36306	:douta	=	16'h	3a4c;
36307	:douta	=	16'h	31ea;
36308	:douta	=	16'h	18c4;
36309	:douta	=	16'h	2125;
36310	:douta	=	16'h	2148;
36311	:douta	=	16'h	1084;
36312	:douta	=	16'h	1905;
36313	:douta	=	16'h	63d3;
36314	:douta	=	16'h	7cb7;
36315	:douta	=	16'h	9d7a;
36316	:douta	=	16'h	7456;
36317	:douta	=	16'h	8d18;
36318	:douta	=	16'h	a599;
36319	:douta	=	16'h	63d2;
36320	:douta	=	16'h	428d;
36321	:douta	=	16'h	3187;
36322	:douta	=	16'h	5227;
36323	:douta	=	16'h	5162;
36324	:douta	=	16'h	71e2;
36325	:douta	=	16'h	7203;
36326	:douta	=	16'h	7a44;
36327	:douta	=	16'h	7244;
36328	:douta	=	16'h	7244;
36329	:douta	=	16'h	7265;
36330	:douta	=	16'h	6a25;
36331	:douta	=	16'h	6a25;
36332	:douta	=	16'h	6a45;
36333	:douta	=	16'h	6a25;
36334	:douta	=	16'h	6a25;
36335	:douta	=	16'h	6a25;
36336	:douta	=	16'h	6206;
36337	:douta	=	16'h	6a05;
36338	:douta	=	16'h	61e5;
36339	:douta	=	16'h	61e5;
36340	:douta	=	16'h	59e5;
36341	:douta	=	16'h	59e5;
36342	:douta	=	16'h	59e5;
36343	:douta	=	16'h	49a6;
36344	:douta	=	16'h	7b2e;
36345	:douta	=	16'h	41c7;
36346	:douta	=	16'h	49e8;
36347	:douta	=	16'h	49e8;
36348	:douta	=	16'h	49e8;
36349	:douta	=	16'h	5228;
36350	:douta	=	16'h	49e8;
36351	:douta	=	16'h	3987;
36352	:douta	=	16'h	edae;
36353	:douta	=	16'h	e5ad;
36354	:douta	=	16'h	e56d;
36355	:douta	=	16'h	e56c;
36356	:douta	=	16'h	edac;
36357	:douta	=	16'h	cd0a;
36358	:douta	=	16'h	6226;
36359	:douta	=	16'h	7267;
36360	:douta	=	16'h	4964;
36361	:douta	=	16'h	d5b6;
36362	:douta	=	16'h	bd13;
36363	:douta	=	16'h	9c72;
36364	:douta	=	16'h	9432;
36365	:douta	=	16'h	7b4e;
36366	:douta	=	16'h	dd93;
36367	:douta	=	16'h	d5d5;
36368	:douta	=	16'h	bd97;
36369	:douta	=	16'h	bd98;
36370	:douta	=	16'h	73f3;
36371	:douta	=	16'h	6393;
36372	:douta	=	16'h	6c14;
36373	:douta	=	16'h	29c9;
36374	:douta	=	16'h	1927;
36375	:douta	=	16'h	2188;
36376	:douta	=	16'h	21a9;
36377	:douta	=	16'h	29ca;
36378	:douta	=	16'h	322c;
36379	:douta	=	16'h	2a0b;
36380	:douta	=	16'h	322c;
36381	:douta	=	16'h	322c;
36382	:douta	=	16'h	3a4d;
36383	:douta	=	16'h	320b;
36384	:douta	=	16'h	320b;
36385	:douta	=	16'h	3a4c;
36386	:douta	=	16'h	320b;
36387	:douta	=	16'h	29ca;
36388	:douta	=	16'h	3a4c;
36389	:douta	=	16'h	3a6c;
36390	:douta	=	16'h	3a4c;
36391	:douta	=	16'h	322b;
36392	:douta	=	16'h	3a4c;
36393	:douta	=	16'h	3a6c;
36394	:douta	=	16'h	3a8c;
36395	:douta	=	16'h	3a6b;
36396	:douta	=	16'h	3a6b;
36397	:douta	=	16'h	42ac;
36398	:douta	=	16'h	3a8c;
36399	:douta	=	16'h	42ad;
36400	:douta	=	16'h	42ac;
36401	:douta	=	16'h	4acd;
36402	:douta	=	16'h	530e;
36403	:douta	=	16'h	5b2e;
36404	:douta	=	16'h	5b2e;
36405	:douta	=	16'h	5b4f;
36406	:douta	=	16'h	5b4f;
36407	:douta	=	16'h	5b2f;
36408	:douta	=	16'h	530e;
36409	:douta	=	16'h	4b0e;
36410	:douta	=	16'h	532e;
36411	:douta	=	16'h	4aad;
36412	:douta	=	16'h	4aed;
36413	:douta	=	16'h	530e;
36414	:douta	=	16'h	532e;
36415	:douta	=	16'h	530e;
36416	:douta	=	16'h	534f;
36417	:douta	=	16'h	534f;
36418	:douta	=	16'h	63b0;
36419	:douta	=	16'h	5b6f;
36420	:douta	=	16'h	6390;
36421	:douta	=	16'h	6390;
36422	:douta	=	16'h	6390;
36423	:douta	=	16'h	638f;
36424	:douta	=	16'h	6390;
36425	:douta	=	16'h	636f;
36426	:douta	=	16'h	638f;
36427	:douta	=	16'h	638f;
36428	:douta	=	16'h	6bd0;
36429	:douta	=	16'h	6390;
36430	:douta	=	16'h	73d0;
36431	:douta	=	16'h	8c0f;
36432	:douta	=	16'h	93ef;
36433	:douta	=	16'h	940f;
36434	:douta	=	16'h	8bcf;
36435	:douta	=	16'h	83cf;
36436	:douta	=	16'h	7b8e;
36437	:douta	=	16'h	7b8e;
36438	:douta	=	16'h	7bcf;
36439	:douta	=	16'h	7baf;
36440	:douta	=	16'h	6b2c;
36441	:douta	=	16'h	6b0c;
36442	:douta	=	16'h	528b;
36443	:douta	=	16'h	7b0c;
36444	:douta	=	16'h	cd10;
36445	:douta	=	16'h	eeb7;
36446	:douta	=	16'h	cdd4;
36447	:douta	=	16'h	eeb7;
36448	:douta	=	16'h	bd74;
36449	:douta	=	16'h	e676;
36450	:douta	=	16'h	a536;
36451	:douta	=	16'h	a537;
36452	:douta	=	16'h	a516;
36453	:douta	=	16'h	94d6;
36454	:douta	=	16'h	8c95;
36455	:douta	=	16'h	8c95;
36456	:douta	=	16'h	8413;
36457	:douta	=	16'h	5aee;
36458	:douta	=	16'h	9493;
36459	:douta	=	16'h	7bf1;
36460	:douta	=	16'h	6b6f;
36461	:douta	=	16'h	6b6f;
36462	:douta	=	16'h	6b4f;
36463	:douta	=	16'h	630e;
36464	:douta	=	16'h	62ed;
36465	:douta	=	16'h	5a8c;
36466	:douta	=	16'h	a3ee;
36467	:douta	=	16'h	ee55;
36468	:douta	=	16'h	b4d1;
36469	:douta	=	16'h	cdb3;
36470	:douta	=	16'h	acd3;
36471	:douta	=	16'h	a4f4;
36472	:douta	=	16'h	9cd5;
36473	:douta	=	16'h	94b4;
36474	:douta	=	16'h	9cf6;
36475	:douta	=	16'h	7413;
36476	:douta	=	16'h	634f;
36477	:douta	=	16'h	322d;
36478	:douta	=	16'h	3a0a;
36479	:douta	=	16'h	52ac;
36480	:douta	=	16'h	7b4e;
36481	:douta	=	16'h	7b4e;
36482	:douta	=	16'h	7b4d;
36483	:douta	=	16'h	62cb;
36484	:douta	=	16'h	4a09;
36485	:douta	=	16'h	a40f;
36486	:douta	=	16'h	8c32;
36487	:douta	=	16'h	5ace;
36488	:douta	=	16'h	9412;
36489	:douta	=	16'h	83d1;
36490	:douta	=	16'h	62ed;
36491	:douta	=	16'h	6b0e;
36492	:douta	=	16'h	5a8c;
36493	:douta	=	16'h	29aa;
36494	:douta	=	16'h	4a2b;
36495	:douta	=	16'h	6b0c;
36496	:douta	=	16'h	6aeb;
36497	:douta	=	16'h	4a29;
36498	:douta	=	16'h	41a8;
36499	:douta	=	16'h	3167;
36500	:douta	=	16'h	41e8;
36501	:douta	=	16'h	93cf;
36502	:douta	=	16'h	b556;
36503	:douta	=	16'h	8c74;
36504	:douta	=	16'h	9c94;
36505	:douta	=	16'h	94b6;
36506	:douta	=	16'h	8454;
36507	:douta	=	16'h	73d2;
36508	:douta	=	16'h	9c92;
36509	:douta	=	16'h	7bd1;
36510	:douta	=	16'h	8432;
36511	:douta	=	16'h	8c52;
36512	:douta	=	16'h	73b0;
36513	:douta	=	16'h	7bd1;
36514	:douta	=	16'h	7bd1;
36515	:douta	=	16'h	7bb0;
36516	:douta	=	16'h	736f;
36517	:douta	=	16'h	6b2e;
36518	:douta	=	16'h	528c;
36519	:douta	=	16'h	528c;
36520	:douta	=	16'h	7b6d;
36521	:douta	=	16'h	9c50;
36522	:douta	=	16'h	ee75;
36523	:douta	=	16'h	ee96;
36524	:douta	=	16'h	cdb5;
36525	:douta	=	16'h	b554;
36526	:douta	=	16'h	b535;
36527	:douta	=	16'h	bd75;
36528	:douta	=	16'h	c575;
36529	:douta	=	16'h	cdd6;
36530	:douta	=	16'h	a4b2;
36531	:douta	=	16'h	ad14;
36532	:douta	=	16'h	ad15;
36533	:douta	=	16'h	9cd4;
36534	:douta	=	16'h	a4f5;
36535	:douta	=	16'h	9473;
36536	:douta	=	16'h	8c73;
36537	:douta	=	16'h	9494;
36538	:douta	=	16'h	8c53;
36539	:douta	=	16'h	8433;
36540	:douta	=	16'h	8432;
36541	:douta	=	16'h	8432;
36542	:douta	=	16'h	8432;
36543	:douta	=	16'h	7c12;
36544	:douta	=	16'h	6b70;
36545	:douta	=	16'h	6b90;
36546	:douta	=	16'h	6b50;
36547	:douta	=	16'h	6350;
36548	:douta	=	16'h	52ad;
36549	:douta	=	16'h	5aac;
36550	:douta	=	16'h	ac8e;
36551	:douta	=	16'h	cd92;
36552	:douta	=	16'h	de14;
36553	:douta	=	16'h	cdd3;
36554	:douta	=	16'h	cd73;
36555	:douta	=	16'h	6371;
36556	:douta	=	16'h	324d;
36557	:douta	=	16'h	73d1;
36558	:douta	=	16'h	6350;
36559	:douta	=	16'h	322c;
36560	:douta	=	16'h	324c;
36561	:douta	=	16'h	31ea;
36562	:douta	=	16'h	18e5;
36563	:douta	=	16'h	3a4c;
36564	:douta	=	16'h	1083;
36565	:douta	=	16'h	2147;
36566	:douta	=	16'h	2168;
36567	:douta	=	16'h	10e5;
36568	:douta	=	16'h	10e5;
36569	:douta	=	16'h	29ca;
36570	:douta	=	16'h	6c36;
36571	:douta	=	16'h	6c14;
36572	:douta	=	16'h	63b3;
36573	:douta	=	16'h	4b10;
36574	:douta	=	16'h	9558;
36575	:douta	=	16'h	20a2;
36576	:douta	=	16'h	1860;
36577	:douta	=	16'h	4963;
36578	:douta	=	16'h	61c3;
36579	:douta	=	16'h	7a44;
36580	:douta	=	16'h	7a65;
36581	:douta	=	16'h	7a65;
36582	:douta	=	16'h	7245;
36583	:douta	=	16'h	7245;
36584	:douta	=	16'h	7245;
36585	:douta	=	16'h	7225;
36586	:douta	=	16'h	6a04;
36587	:douta	=	16'h	6a24;
36588	:douta	=	16'h	6a25;
36589	:douta	=	16'h	6a25;
36590	:douta	=	16'h	6a25;
36591	:douta	=	16'h	6205;
36592	:douta	=	16'h	6a05;
36593	:douta	=	16'h	6205;
36594	:douta	=	16'h	61e5;
36595	:douta	=	16'h	61e5;
36596	:douta	=	16'h	59e5;
36597	:douta	=	16'h	59c5;
36598	:douta	=	16'h	59c5;
36599	:douta	=	16'h	4964;
36600	:douta	=	16'h	8bf0;
36601	:douta	=	16'h	838f;
36602	:douta	=	16'h	49e7;
36603	:douta	=	16'h	4a08;
36604	:douta	=	16'h	5209;
36605	:douta	=	16'h	49e8;
36606	:douta	=	16'h	41a7;
36607	:douta	=	16'h	41c7;
36608	:douta	=	16'h	e5ae;
36609	:douta	=	16'h	e58d;
36610	:douta	=	16'h	e56c;
36611	:douta	=	16'h	e56c;
36612	:douta	=	16'h	e56b;
36613	:douta	=	16'h	edcc;
36614	:douta	=	16'h	6205;
36615	:douta	=	16'h	7aa8;
36616	:douta	=	16'h	8aeb;
36617	:douta	=	16'h	cd54;
36618	:douta	=	16'h	b4b2;
36619	:douta	=	16'h	ac92;
36620	:douta	=	16'h	ac71;
36621	:douta	=	16'h	c4b0;
36622	:douta	=	16'h	ee77;
36623	:douta	=	16'h	e676;
36624	:douta	=	16'h	b515;
36625	:douta	=	16'h	b536;
36626	:douta	=	16'h	6bb3;
36627	:douta	=	16'h	7c55;
36628	:douta	=	16'h	7c76;
36629	:douta	=	16'h	8d18;
36630	:douta	=	16'h	322b;
36631	:douta	=	16'h	1927;
36632	:douta	=	16'h	31ea;
36633	:douta	=	16'h	320a;
36634	:douta	=	16'h	322c;
36635	:douta	=	16'h	326d;
36636	:douta	=	16'h	326d;
36637	:douta	=	16'h	3a8d;
36638	:douta	=	16'h	3a8d;
36639	:douta	=	16'h	3a8d;
36640	:douta	=	16'h	322c;
36641	:douta	=	16'h	3a4c;
36642	:douta	=	16'h	3a6d;
36643	:douta	=	16'h	3a4c;
36644	:douta	=	16'h	29ca;
36645	:douta	=	16'h	29ea;
36646	:douta	=	16'h	2a0a;
36647	:douta	=	16'h	3a6c;
36648	:douta	=	16'h	3a4c;
36649	:douta	=	16'h	3a6c;
36650	:douta	=	16'h	42ad;
36651	:douta	=	16'h	3a8c;
36652	:douta	=	16'h	3a8d;
36653	:douta	=	16'h	3a4c;
36654	:douta	=	16'h	324b;
36655	:douta	=	16'h	3a6b;
36656	:douta	=	16'h	42cd;
36657	:douta	=	16'h	530f;
36658	:douta	=	16'h	5b0e;
36659	:douta	=	16'h	636f;
36660	:douta	=	16'h	5b4e;
36661	:douta	=	16'h	636f;
36662	:douta	=	16'h	6370;
36663	:douta	=	16'h	634f;
36664	:douta	=	16'h	534f;
36665	:douta	=	16'h	532e;
36666	:douta	=	16'h	4b0e;
36667	:douta	=	16'h	532e;
36668	:douta	=	16'h	530e;
36669	:douta	=	16'h	5b4f;
36670	:douta	=	16'h	532f;
36671	:douta	=	16'h	534f;
36672	:douta	=	16'h	532e;
36673	:douta	=	16'h	534f;
36674	:douta	=	16'h	534f;
36675	:douta	=	16'h	5b4f;
36676	:douta	=	16'h	5b2f;
36677	:douta	=	16'h	63d1;
36678	:douta	=	16'h	5b6f;
36679	:douta	=	16'h	5b6f;
36680	:douta	=	16'h	5b4f;
36681	:douta	=	16'h	6390;
36682	:douta	=	16'h	5b6f;
36683	:douta	=	16'h	638f;
36684	:douta	=	16'h	638f;
36685	:douta	=	16'h	634e;
36686	:douta	=	16'h	6b90;
36687	:douta	=	16'h	6bd0;
36688	:douta	=	16'h	638f;
36689	:douta	=	16'h	6baf;
36690	:douta	=	16'h	6baf;
36691	:douta	=	16'h	736e;
36692	:douta	=	16'h	734c;
36693	:douta	=	16'h	732d;
36694	:douta	=	16'h	732c;
36695	:douta	=	16'h	72cb;
36696	:douta	=	16'h	5a8a;
36697	:douta	=	16'h	62ab;
36698	:douta	=	16'h	ddb3;
36699	:douta	=	16'h	de55;
36700	:douta	=	16'h	eeb7;
36701	:douta	=	16'h	b514;
36702	:douta	=	16'h	e656;
36703	:douta	=	16'h	c574;
36704	:douta	=	16'h	b555;
36705	:douta	=	16'h	bd76;
36706	:douta	=	16'h	ad36;
36707	:douta	=	16'h	9d17;
36708	:douta	=	16'h	94b6;
36709	:douta	=	16'h	94b6;
36710	:douta	=	16'h	8c75;
36711	:douta	=	16'h	7bf2;
36712	:douta	=	16'h	7bd1;
36713	:douta	=	16'h	7bf1;
36714	:douta	=	16'h	6b4f;
36715	:douta	=	16'h	7bf1;
36716	:douta	=	16'h	73b1;
36717	:douta	=	16'h	6b6f;
36718	:douta	=	16'h	734f;
36719	:douta	=	16'h	4a6c;
36720	:douta	=	16'h	730d;
36721	:douta	=	16'h	e614;
36722	:douta	=	16'h	ddf4;
36723	:douta	=	16'h	d593;
36724	:douta	=	16'h	8c54;
36725	:douta	=	16'h	b4f4;
36726	:douta	=	16'h	94b5;
36727	:douta	=	16'h	9cd5;
36728	:douta	=	16'h	8c95;
36729	:douta	=	16'h	8433;
36730	:douta	=	16'h	7c12;
36731	:douta	=	16'h	6b90;
36732	:douta	=	16'h	6b6f;
36733	:douta	=	16'h	736e;
36734	:douta	=	16'h	528c;
36735	:douta	=	16'h	3a2b;
36736	:douta	=	16'h	29ca;
36737	:douta	=	16'h	29ca;
36738	:douta	=	16'h	29aa;
36739	:douta	=	16'h	93f0;
36740	:douta	=	16'h	b4d4;
36741	:douta	=	16'h	8412;
36742	:douta	=	16'h	73f2;
36743	:douta	=	16'h	424c;
36744	:douta	=	16'h	4a4c;
36745	:douta	=	16'h	732d;
36746	:douta	=	16'h	734e;
36747	:douta	=	16'h	6b0c;
36748	:douta	=	16'h	6b0c;
36749	:douta	=	16'h	72ec;
36750	:douta	=	16'h	5aab;
36751	:douta	=	16'h	522a;
36752	:douta	=	16'h	39e9;
36753	:douta	=	16'h	3987;
36754	:douta	=	16'h	732c;
36755	:douta	=	16'h	c511;
36756	:douta	=	16'h	d593;
36757	:douta	=	16'h	b4d3;
36758	:douta	=	16'h	a4f6;
36759	:douta	=	16'h	73d2;
36760	:douta	=	16'h	6b91;
36761	:douta	=	16'h	8c53;
36762	:douta	=	16'h	8453;
36763	:douta	=	16'h	7bf2;
36764	:douta	=	16'h	73b1;
36765	:douta	=	16'h	9493;
36766	:douta	=	16'h	5b0f;
36767	:douta	=	16'h	3a6d;
36768	:douta	=	16'h	52ce;
36769	:douta	=	16'h	7390;
36770	:douta	=	16'h	734f;
36771	:douta	=	16'h	6b4e;
36772	:douta	=	16'h	630d;
36773	:douta	=	16'h	734f;
36774	:douta	=	16'h	c552;
36775	:douta	=	16'h	d5d4;
36776	:douta	=	16'h	de77;
36777	:douta	=	16'h	de56;
36778	:douta	=	16'h	e676;
36779	:douta	=	16'h	de15;
36780	:douta	=	16'h	c595;
36781	:douta	=	16'h	b555;
36782	:douta	=	16'h	b536;
36783	:douta	=	16'h	8c51;
36784	:douta	=	16'h	8c51;
36785	:douta	=	16'h	8c11;
36786	:douta	=	16'h	8c31;
36787	:douta	=	16'h	9c93;
36788	:douta	=	16'h	ad35;
36789	:douta	=	16'h	a4f5;
36790	:douta	=	16'h	9cf5;
36791	:douta	=	16'h	9474;
36792	:douta	=	16'h	8c73;
36793	:douta	=	16'h	8433;
36794	:douta	=	16'h	8c53;
36795	:douta	=	16'h	83f2;
36796	:douta	=	16'h	7390;
36797	:douta	=	16'h	736f;
36798	:douta	=	16'h	73b0;
36799	:douta	=	16'h	6b90;
36800	:douta	=	16'h	6b90;
36801	:douta	=	16'h	62ed;
36802	:douta	=	16'h	528b;
36803	:douta	=	16'h	6aeb;
36804	:douta	=	16'h	8bee;
36805	:douta	=	16'h	ad10;
36806	:douta	=	16'h	cdb4;
36807	:douta	=	16'h	de34;
36808	:douta	=	16'h	ddd4;
36809	:douta	=	16'h	cd94;
36810	:douta	=	16'h	ad14;
36811	:douta	=	16'h	7c13;
36812	:douta	=	16'h	530f;
36813	:douta	=	16'h	6b90;
36814	:douta	=	16'h	5b50;
36815	:douta	=	16'h	4aef;
36816	:douta	=	16'h	42cf;
36817	:douta	=	16'h	428e;
36818	:douta	=	16'h	322d;
36819	:douta	=	16'h	29ca;
36820	:douta	=	16'h	3a4d;
36821	:douta	=	16'h	2126;
36822	:douta	=	16'h	29a8;
36823	:douta	=	16'h	2988;
36824	:douta	=	16'h	2147;
36825	:douta	=	16'h	1906;
36826	:douta	=	16'h	5371;
36827	:douta	=	16'h	9d59;
36828	:douta	=	16'h	a5da;
36829	:douta	=	16'h	7cd8;
36830	:douta	=	16'h	1020;
36831	:douta	=	16'h	2904;
36832	:douta	=	16'h	59a4;
36833	:douta	=	16'h	8264;
36834	:douta	=	16'h	7a44;
36835	:douta	=	16'h	7a44;
36836	:douta	=	16'h	7a65;
36837	:douta	=	16'h	7a45;
36838	:douta	=	16'h	7244;
36839	:douta	=	16'h	7245;
36840	:douta	=	16'h	7224;
36841	:douta	=	16'h	6a25;
36842	:douta	=	16'h	6a24;
36843	:douta	=	16'h	6a24;
36844	:douta	=	16'h	6a04;
36845	:douta	=	16'h	6a05;
36846	:douta	=	16'h	6205;
36847	:douta	=	16'h	6205;
36848	:douta	=	16'h	6205;
36849	:douta	=	16'h	61e5;
36850	:douta	=	16'h	59e5;
36851	:douta	=	16'h	61e5;
36852	:douta	=	16'h	59e5;
36853	:douta	=	16'h	59e5;
36854	:douta	=	16'h	59c5;
36855	:douta	=	16'h	51c6;
36856	:douta	=	16'h	4964;
36857	:douta	=	16'h	4144;
36858	:douta	=	16'h	7b4e;
36859	:douta	=	16'h	5208;
36860	:douta	=	16'h	41a7;
36861	:douta	=	16'h	49e7;
36862	:douta	=	16'h	49e8;
36863	:douta	=	16'h	41c8;
36864	:douta	=	16'h	edae;
36865	:douta	=	16'h	e58e;
36866	:douta	=	16'h	e58d;
36867	:douta	=	16'h	e56c;
36868	:douta	=	16'h	dd6c;
36869	:douta	=	16'h	f5ed;
36870	:douta	=	16'h	6a26;
36871	:douta	=	16'h	8ae8;
36872	:douta	=	16'h	9bae;
36873	:douta	=	16'h	bcf2;
36874	:douta	=	16'h	b492;
36875	:douta	=	16'h	ac91;
36876	:douta	=	16'h	b4b1;
36877	:douta	=	16'h	e5b3;
36878	:douta	=	16'h	ee56;
36879	:douta	=	16'h	ee97;
36880	:douta	=	16'h	b514;
36881	:douta	=	16'h	a4f5;
36882	:douta	=	16'h	63b2;
36883	:douta	=	16'h	7c76;
36884	:douta	=	16'h	84b7;
36885	:douta	=	16'h	6c14;
36886	:douta	=	16'h	1106;
36887	:douta	=	16'h	2168;
36888	:douta	=	16'h	2188;
36889	:douta	=	16'h	29a9;
36890	:douta	=	16'h	2a2b;
36891	:douta	=	16'h	322d;
36892	:douta	=	16'h	324d;
36893	:douta	=	16'h	3a8e;
36894	:douta	=	16'h	3a8e;
36895	:douta	=	16'h	3a8e;
36896	:douta	=	16'h	3a8d;
36897	:douta	=	16'h	3a8d;
36898	:douta	=	16'h	3a8d;
36899	:douta	=	16'h	324c;
36900	:douta	=	16'h	29ca;
36901	:douta	=	16'h	29ca;
36902	:douta	=	16'h	320b;
36903	:douta	=	16'h	320b;
36904	:douta	=	16'h	3a4c;
36905	:douta	=	16'h	3a4c;
36906	:douta	=	16'h	42ad;
36907	:douta	=	16'h	428d;
36908	:douta	=	16'h	428d;
36909	:douta	=	16'h	42ad;
36910	:douta	=	16'h	42ad;
36911	:douta	=	16'h	4ace;
36912	:douta	=	16'h	42ad;
36913	:douta	=	16'h	4aad;
36914	:douta	=	16'h	4aad;
36915	:douta	=	16'h	4aac;
36916	:douta	=	16'h	4aac;
36917	:douta	=	16'h	4acc;
36918	:douta	=	16'h	4acd;
36919	:douta	=	16'h	4aed;
36920	:douta	=	16'h	534f;
36921	:douta	=	16'h	5b6f;
36922	:douta	=	16'h	536f;
36923	:douta	=	16'h	534f;
36924	:douta	=	16'h	532f;
36925	:douta	=	16'h	530e;
36926	:douta	=	16'h	532e;
36927	:douta	=	16'h	532e;
36928	:douta	=	16'h	5b4f;
36929	:douta	=	16'h	5b4f;
36930	:douta	=	16'h	532f;
36931	:douta	=	16'h	5b4f;
36932	:douta	=	16'h	534f;
36933	:douta	=	16'h	63b1;
36934	:douta	=	16'h	5b4f;
36935	:douta	=	16'h	5b6e;
36936	:douta	=	16'h	5b6f;
36937	:douta	=	16'h	638f;
36938	:douta	=	16'h	636f;
36939	:douta	=	16'h	638f;
36940	:douta	=	16'h	636f;
36941	:douta	=	16'h	636f;
36942	:douta	=	16'h	634f;
36943	:douta	=	16'h	638f;
36944	:douta	=	16'h	638f;
36945	:douta	=	16'h	63b0;
36946	:douta	=	16'h	638f;
36947	:douta	=	16'h	6bd0;
36948	:douta	=	16'h	6b6e;
36949	:douta	=	16'h	6b6d;
36950	:douta	=	16'h	7bae;
36951	:douta	=	16'h	738e;
36952	:douta	=	16'h	8bce;
36953	:douta	=	16'h	b4b2;
36954	:douta	=	16'h	eed7;
36955	:douta	=	16'h	e676;
36956	:douta	=	16'h	e6b7;
36957	:douta	=	16'h	a4d4;
36958	:douta	=	16'h	c5b6;
36959	:douta	=	16'h	bd75;
36960	:douta	=	16'h	b556;
36961	:douta	=	16'h	b556;
36962	:douta	=	16'h	b596;
36963	:douta	=	16'h	94f6;
36964	:douta	=	16'h	8c54;
36965	:douta	=	16'h	9495;
36966	:douta	=	16'h	8433;
36967	:douta	=	16'h	6b6f;
36968	:douta	=	16'h	6b6f;
36969	:douta	=	16'h	7390;
36970	:douta	=	16'h	734f;
36971	:douta	=	16'h	7b90;
36972	:douta	=	16'h	8412;
36973	:douta	=	16'h	83d0;
36974	:douta	=	16'h	632f;
36975	:douta	=	16'h	8b4c;
36976	:douta	=	16'h	dd92;
36977	:douta	=	16'h	d593;
36978	:douta	=	16'h	ddf3;
36979	:douta	=	16'h	c553;
36980	:douta	=	16'h	8c74;
36981	:douta	=	16'h	9c94;
36982	:douta	=	16'h	8c74;
36983	:douta	=	16'h	8c74;
36984	:douta	=	16'h	8454;
36985	:douta	=	16'h	7bf2;
36986	:douta	=	16'h	7c12;
36987	:douta	=	16'h	73b0;
36988	:douta	=	16'h	6b6f;
36989	:douta	=	16'h	6b0d;
36990	:douta	=	16'h	62cb;
36991	:douta	=	16'h	62ab;
36992	:douta	=	16'h	62ab;
36993	:douta	=	16'h	5a8b;
36994	:douta	=	16'h	7b2c;
36995	:douta	=	16'h	b4f4;
36996	:douta	=	16'h	8c53;
36997	:douta	=	16'h	73f2;
36998	:douta	=	16'h	73b1;
36999	:douta	=	16'h	52ad;
37000	:douta	=	16'h	31eb;
37001	:douta	=	16'h	3a2b;
37002	:douta	=	16'h	732d;
37003	:douta	=	16'h	7b6d;
37004	:douta	=	16'h	6aec;
37005	:douta	=	16'h	6acb;
37006	:douta	=	16'h	6aab;
37007	:douta	=	16'h	72ec;
37008	:douta	=	16'h	5a6a;
37009	:douta	=	16'h	5aac;
37010	:douta	=	16'h	e5f4;
37011	:douta	=	16'h	e5d4;
37012	:douta	=	16'h	bd54;
37013	:douta	=	16'h	acf4;
37014	:douta	=	16'h	9cd5;
37015	:douta	=	16'h	8454;
37016	:douta	=	16'h	6b72;
37017	:douta	=	16'h	6b70;
37018	:douta	=	16'h	8c32;
37019	:douta	=	16'h	7bf1;
37020	:douta	=	16'h	632f;
37021	:douta	=	16'h	7390;
37022	:douta	=	16'h	83f2;
37023	:douta	=	16'h	6b4f;
37024	:douta	=	16'h	31ec;
37025	:douta	=	16'h	424d;
37026	:douta	=	16'h	426d;
37027	:douta	=	16'h	4a8c;
37028	:douta	=	16'h	6b2d;
37029	:douta	=	16'h	cd72;
37030	:douta	=	16'h	de35;
37031	:douta	=	16'h	bd33;
37032	:douta	=	16'h	de35;
37033	:douta	=	16'h	d616;
37034	:douta	=	16'h	c5b5;
37035	:douta	=	16'h	c595;
37036	:douta	=	16'h	bd76;
37037	:douta	=	16'h	b535;
37038	:douta	=	16'h	ad36;
37039	:douta	=	16'h	a515;
37040	:douta	=	16'h	9cd4;
37041	:douta	=	16'h	8c32;
37042	:douta	=	16'h	9452;
37043	:douta	=	16'h	8c31;
37044	:douta	=	16'h	9cb3;
37045	:douta	=	16'h	9cb4;
37046	:douta	=	16'h	9cd4;
37047	:douta	=	16'h	9494;
37048	:douta	=	16'h	8c73;
37049	:douta	=	16'h	7bf1;
37050	:douta	=	16'h	7bd1;
37051	:douta	=	16'h	7bf2;
37052	:douta	=	16'h	7bd1;
37053	:douta	=	16'h	73b0;
37054	:douta	=	16'h	73d1;
37055	:douta	=	16'h	7bb1;
37056	:douta	=	16'h	5acc;
37057	:douta	=	16'h	5a49;
37058	:douta	=	16'h	6aeb;
37059	:douta	=	16'h	c531;
37060	:douta	=	16'h	d5d3;
37061	:douta	=	16'h	eeb6;
37062	:douta	=	16'h	e676;
37063	:douta	=	16'h	d5f4;
37064	:douta	=	16'h	c554;
37065	:douta	=	16'h	b534;
37066	:douta	=	16'h	9cd5;
37067	:douta	=	16'h	8c95;
37068	:douta	=	16'h	7c54;
37069	:douta	=	16'h	6bb1;
37070	:douta	=	16'h	5b50;
37071	:douta	=	16'h	5351;
37072	:douta	=	16'h	4b10;
37073	:douta	=	16'h	4aaf;
37074	:douta	=	16'h	3a6e;
37075	:douta	=	16'h	324d;
37076	:douta	=	16'h	21a9;
37077	:douta	=	16'h	1926;
37078	:douta	=	16'h	31a9;
37079	:douta	=	16'h	2167;
37080	:douta	=	16'h	1927;
37081	:douta	=	16'h	2127;
37082	:douta	=	16'h	08a4;
37083	:douta	=	16'h	08a4;
37084	:douta	=	16'h	8cf7;
37085	:douta	=	16'h	6c56;
37086	:douta	=	16'h	1021;
37087	:douta	=	16'h	51a4;
37088	:douta	=	16'h	7a63;
37089	:douta	=	16'h	7a65;
37090	:douta	=	16'h	7a65;
37091	:douta	=	16'h	7a65;
37092	:douta	=	16'h	7a44;
37093	:douta	=	16'h	7245;
37094	:douta	=	16'h	7244;
37095	:douta	=	16'h	7224;
37096	:douta	=	16'h	7224;
37097	:douta	=	16'h	6a24;
37098	:douta	=	16'h	6a04;
37099	:douta	=	16'h	6204;
37100	:douta	=	16'h	6205;
37101	:douta	=	16'h	6205;
37102	:douta	=	16'h	61e4;
37103	:douta	=	16'h	6205;
37104	:douta	=	16'h	61e5;
37105	:douta	=	16'h	6205;
37106	:douta	=	16'h	61e5;
37107	:douta	=	16'h	59e5;
37108	:douta	=	16'h	59c5;
37109	:douta	=	16'h	59e5;
37110	:douta	=	16'h	59c5;
37111	:douta	=	16'h	51c5;
37112	:douta	=	16'h	51a5;
37113	:douta	=	16'h	4964;
37114	:douta	=	16'h	49a5;
37115	:douta	=	16'h	4986;
37116	:douta	=	16'h	49e8;
37117	:douta	=	16'h	41a7;
37118	:douta	=	16'h	3965;
37119	:douta	=	16'h	3966;
37120	:douta	=	16'h	ed8e;
37121	:douta	=	16'h	e58d;
37122	:douta	=	16'h	e58d;
37123	:douta	=	16'h	e56c;
37124	:douta	=	16'h	e56e;
37125	:douta	=	16'h	edad;
37126	:douta	=	16'h	8b08;
37127	:douta	=	16'h	7a66;
37128	:douta	=	16'h	e5d5;
37129	:douta	=	16'h	c512;
37130	:douta	=	16'h	c4f3;
37131	:douta	=	16'h	bcb1;
37132	:douta	=	16'h	b470;
37133	:douta	=	16'h	ff18;
37134	:douta	=	16'h	f6f8;
37135	:douta	=	16'h	e697;
37136	:douta	=	16'h	bd35;
37137	:douta	=	16'h	8434;
37138	:douta	=	16'h	7c55;
37139	:douta	=	16'h	8496;
37140	:douta	=	16'h	8cd7;
37141	:douta	=	16'h	2147;
37142	:douta	=	16'h	0882;
37143	:douta	=	16'h	10e5;
37144	:douta	=	16'h	29a9;
37145	:douta	=	16'h	29ca;
37146	:douta	=	16'h	2a2b;
37147	:douta	=	16'h	2a0c;
37148	:douta	=	16'h	322d;
37149	:douta	=	16'h	324d;
37150	:douta	=	16'h	3a8e;
37151	:douta	=	16'h	3a6d;
37152	:douta	=	16'h	326d;
37153	:douta	=	16'h	3a8d;
37154	:douta	=	16'h	3a8d;
37155	:douta	=	16'h	3a6d;
37156	:douta	=	16'h	21ca;
37157	:douta	=	16'h	29ea;
37158	:douta	=	16'h	3a4c;
37159	:douta	=	16'h	2a0b;
37160	:douta	=	16'h	2a0b;
37161	:douta	=	16'h	324c;
37162	:douta	=	16'h	324b;
37163	:douta	=	16'h	3a8d;
37164	:douta	=	16'h	42ad;
37165	:douta	=	16'h	3a6c;
37166	:douta	=	16'h	2167;
37167	:douta	=	16'h	2125;
37168	:douta	=	16'h	2125;
37169	:douta	=	16'h	2125;
37170	:douta	=	16'h	2926;
37171	:douta	=	16'h	31a7;
37172	:douta	=	16'h	39c8;
37173	:douta	=	16'h	31c8;
37174	:douta	=	16'h	31a7;
37175	:douta	=	16'h	2987;
37176	:douta	=	16'h	2967;
37177	:douta	=	16'h	2146;
37178	:douta	=	16'h	2125;
37179	:douta	=	16'h	2967;
37180	:douta	=	16'h	29c8;
37181	:douta	=	16'h	42ac;
37182	:douta	=	16'h	42ee;
37183	:douta	=	16'h	5350;
37184	:douta	=	16'h	42ce;
37185	:douta	=	16'h	42cd;
37186	:douta	=	16'h	4b0e;
37187	:douta	=	16'h	530e;
37188	:douta	=	16'h	5b4f;
37189	:douta	=	16'h	5b4f;
37190	:douta	=	16'h	532e;
37191	:douta	=	16'h	5b4e;
37192	:douta	=	16'h	5b4f;
37193	:douta	=	16'h	5b4f;
37194	:douta	=	16'h	636f;
37195	:douta	=	16'h	5b4e;
37196	:douta	=	16'h	636f;
37197	:douta	=	16'h	6b90;
37198	:douta	=	16'h	638f;
37199	:douta	=	16'h	638f;
37200	:douta	=	16'h	638f;
37201	:douta	=	16'h	638f;
37202	:douta	=	16'h	638f;
37203	:douta	=	16'h	6b8f;
37204	:douta	=	16'h	638f;
37205	:douta	=	16'h	6b90;
37206	:douta	=	16'h	638f;
37207	:douta	=	16'h	6b90;
37208	:douta	=	16'h	5b4e;
37209	:douta	=	16'h	532e;
37210	:douta	=	16'h	8c10;
37211	:douta	=	16'h	cdb6;
37212	:douta	=	16'h	c595;
37213	:douta	=	16'h	b556;
37214	:douta	=	16'h	b556;
37215	:douta	=	16'h	bd96;
37216	:douta	=	16'h	a516;
37217	:douta	=	16'h	a4f5;
37218	:douta	=	16'h	9cf5;
37219	:douta	=	16'h	9cd6;
37220	:douta	=	16'h	7bd1;
37221	:douta	=	16'h	7390;
37222	:douta	=	16'h	7bf1;
37223	:douta	=	16'h	7bd1;
37224	:douta	=	16'h	7390;
37225	:douta	=	16'h	7bd0;
37226	:douta	=	16'h	736f;
37227	:douta	=	16'h	732e;
37228	:douta	=	16'h	5acd;
37229	:douta	=	16'h	5a8c;
37230	:douta	=	16'h	cd31;
37231	:douta	=	16'h	f6b4;
37232	:douta	=	16'h	d593;
37233	:douta	=	16'h	acf4;
37234	:douta	=	16'h	b515;
37235	:douta	=	16'h	9cd6;
37236	:douta	=	16'h	8c74;
37237	:douta	=	16'h	8453;
37238	:douta	=	16'h	94b5;
37239	:douta	=	16'h	8413;
37240	:douta	=	16'h	7390;
37241	:douta	=	16'h	6b70;
37242	:douta	=	16'h	6b0e;
37243	:douta	=	16'h	62cc;
37244	:douta	=	16'h	6acc;
37245	:douta	=	16'h	62ec;
37246	:douta	=	16'h	62cc;
37247	:douta	=	16'h	5a49;
37248	:douta	=	16'h	5a6b;
37249	:douta	=	16'h	62cd;
37250	:douta	=	16'h	93f0;
37251	:douta	=	16'h	8c94;
37252	:douta	=	16'h	7433;
37253	:douta	=	16'h	6b4f;
37254	:douta	=	16'h	630e;
37255	:douta	=	16'h	62cd;
37256	:douta	=	16'h	62ac;
37257	:douta	=	16'h	424b;
37258	:douta	=	16'h	2988;
37259	:douta	=	16'h	29a8;
37260	:douta	=	16'h	31c8;
37261	:douta	=	16'h	524a;
37262	:douta	=	16'h	5a4b;
37263	:douta	=	16'h	730c;
37264	:douta	=	16'h	c4f0;
37265	:douta	=	16'h	94b4;
37266	:douta	=	16'h	7c12;
37267	:douta	=	16'h	94b5;
37268	:douta	=	16'h	94d5;
37269	:douta	=	16'h	94b5;
37270	:douta	=	16'h	8473;
37271	:douta	=	16'h	7c13;
37272	:douta	=	16'h	8433;
37273	:douta	=	16'h	52ef;
37274	:douta	=	16'h	3a4c;
37275	:douta	=	16'h	52ce;
37276	:douta	=	16'h	7bd0;
37277	:douta	=	16'h	83b0;
37278	:douta	=	16'h	6b4f;
37279	:douta	=	16'h	632e;
37280	:douta	=	16'h	630f;
37281	:douta	=	16'h	8bef;
37282	:douta	=	16'h	acb0;
37283	:douta	=	16'h	e656;
37284	:douta	=	16'h	f6d8;
37285	:douta	=	16'h	d616;
37286	:douta	=	16'h	de57;
37287	:douta	=	16'h	bd74;
37288	:douta	=	16'h	bd95;
37289	:douta	=	16'h	c5b6;
37290	:douta	=	16'h	bd96;
37291	:douta	=	16'h	ad15;
37292	:douta	=	16'h	ad35;
37293	:douta	=	16'h	a515;
37294	:douta	=	16'h	9cf5;
37295	:douta	=	16'h	a4f5;
37296	:douta	=	16'h	9cd4;
37297	:douta	=	16'h	9cd3;
37298	:douta	=	16'h	8c32;
37299	:douta	=	16'h	8c52;
37300	:douta	=	16'h	8411;
37301	:douta	=	16'h	8411;
37302	:douta	=	16'h	7bf1;
37303	:douta	=	16'h	7bf1;
37304	:douta	=	16'h	8432;
37305	:douta	=	16'h	8412;
37306	:douta	=	16'h	8412;
37307	:douta	=	16'h	7bf2;
37308	:douta	=	16'h	738f;
37309	:douta	=	16'h	62cc;
37310	:douta	=	16'h	3144;
37311	:douta	=	16'h	1061;
37312	:douta	=	16'h	a42e;
37313	:douta	=	16'h	cdb2;
37314	:douta	=	16'h	d5d3;
37315	:douta	=	16'h	d5f5;
37316	:douta	=	16'h	d5d4;
37317	:douta	=	16'h	cdb5;
37318	:douta	=	16'h	bd54;
37319	:douta	=	16'h	b535;
37320	:douta	=	16'h	9cf5;
37321	:douta	=	16'h	a515;
37322	:douta	=	16'h	9cf6;
37323	:douta	=	16'h	7c34;
37324	:douta	=	16'h	7434;
37325	:douta	=	16'h	7c55;
37326	:douta	=	16'h	7c55;
37327	:douta	=	16'h	5b31;
37328	:douta	=	16'h	42cf;
37329	:douta	=	16'h	42cf;
37330	:douta	=	16'h	42af;
37331	:douta	=	16'h	3a4d;
37332	:douta	=	16'h	2147;
37333	:douta	=	16'h	4aae;
37334	:douta	=	16'h	5b2f;
37335	:douta	=	16'h	29a8;
37336	:douta	=	16'h	1105;
37337	:douta	=	16'h	0884;
37338	:douta	=	16'h	18e5;
37339	:douta	=	16'h	2968;
37340	:douta	=	16'h	5393;
37341	:douta	=	16'h	42ae;
37342	:douta	=	16'h	3945;
37343	:douta	=	16'h	8284;
37344	:douta	=	16'h	8284;
37345	:douta	=	16'h	7a64;
37346	:douta	=	16'h	7a84;
37347	:douta	=	16'h	7a44;
37348	:douta	=	16'h	7a44;
37349	:douta	=	16'h	7245;
37350	:douta	=	16'h	7244;
37351	:douta	=	16'h	7224;
37352	:douta	=	16'h	6a24;
37353	:douta	=	16'h	6a24;
37354	:douta	=	16'h	6a04;
37355	:douta	=	16'h	6204;
37356	:douta	=	16'h	6204;
37357	:douta	=	16'h	61e4;
37358	:douta	=	16'h	61e4;
37359	:douta	=	16'h	61e5;
37360	:douta	=	16'h	6205;
37361	:douta	=	16'h	61e5;
37362	:douta	=	16'h	59e5;
37363	:douta	=	16'h	61e5;
37364	:douta	=	16'h	59c5;
37365	:douta	=	16'h	59c5;
37366	:douta	=	16'h	59e5;
37367	:douta	=	16'h	51a5;
37368	:douta	=	16'h	4985;
37369	:douta	=	16'h	4964;
37370	:douta	=	16'h	4123;
37371	:douta	=	16'h	4123;
37372	:douta	=	16'h	3923;
37373	:douta	=	16'h	4165;
37374	:douta	=	16'h	49e7;
37375	:douta	=	16'h	630c;
37376	:douta	=	16'h	e5ad;
37377	:douta	=	16'h	e58d;
37378	:douta	=	16'h	e58c;
37379	:douta	=	16'h	e54c;
37380	:douta	=	16'h	e54c;
37381	:douta	=	16'h	e56c;
37382	:douta	=	16'h	a3e8;
37383	:douta	=	16'h	7204;
37384	:douta	=	16'h	f698;
37385	:douta	=	16'h	cd12;
37386	:douta	=	16'h	cd12;
37387	:douta	=	16'h	c4f1;
37388	:douta	=	16'h	c4af;
37389	:douta	=	16'h	ff9b;
37390	:douta	=	16'h	f718;
37391	:douta	=	16'h	eed9;
37392	:douta	=	16'h	acf5;
37393	:douta	=	16'h	7413;
37394	:douta	=	16'h	8496;
37395	:douta	=	16'h	8496;
37396	:douta	=	16'h	8d19;
37397	:douta	=	16'h	29a8;
37398	:douta	=	16'h	6370;
37399	:douta	=	16'h	6bd3;
37400	:douta	=	16'h	428e;
37401	:douta	=	16'h	21aa;
37402	:douta	=	16'h	2a0b;
37403	:douta	=	16'h	2a0b;
37404	:douta	=	16'h	2a0c;
37405	:douta	=	16'h	326d;
37406	:douta	=	16'h	326d;
37407	:douta	=	16'h	3a8e;
37408	:douta	=	16'h	3a8d;
37409	:douta	=	16'h	324d;
37410	:douta	=	16'h	3a8d;
37411	:douta	=	16'h	3aad;
37412	:douta	=	16'h	2189;
37413	:douta	=	16'h	29c9;
37414	:douta	=	16'h	2a0b;
37415	:douta	=	16'h	31eb;
37416	:douta	=	16'h	320b;
37417	:douta	=	16'h	2a0b;
37418	:douta	=	16'h	322b;
37419	:douta	=	16'h	322b;
37420	:douta	=	16'h	29a7;
37421	:douta	=	16'h	2125;
37422	:douta	=	16'h	18c4;
37423	:douta	=	16'h	18e4;
37424	:douta	=	16'h	2125;
37425	:douta	=	16'h	2946;
37426	:douta	=	16'h	2966;
37427	:douta	=	16'h	3187;
37428	:douta	=	16'h	2967;
37429	:douta	=	16'h	31a7;
37430	:douta	=	16'h	2986;
37431	:douta	=	16'h	2966;
37432	:douta	=	16'h	2967;
37433	:douta	=	16'h	2146;
37434	:douta	=	16'h	2126;
37435	:douta	=	16'h	1905;
37436	:douta	=	16'h	18e5;
37437	:douta	=	16'h	1905;
37438	:douta	=	16'h	2147;
37439	:douta	=	16'h	3a6b;
37440	:douta	=	16'h	4b0e;
37441	:douta	=	16'h	532f;
37442	:douta	=	16'h	4aee;
37443	:douta	=	16'h	4aee;
37444	:douta	=	16'h	5b6f;
37445	:douta	=	16'h	534f;
37446	:douta	=	16'h	532e;
37447	:douta	=	16'h	5b4e;
37448	:douta	=	16'h	5b4f;
37449	:douta	=	16'h	5b4e;
37450	:douta	=	16'h	5b4e;
37451	:douta	=	16'h	530e;
37452	:douta	=	16'h	5b2e;
37453	:douta	=	16'h	5b4e;
37454	:douta	=	16'h	638f;
37455	:douta	=	16'h	636e;
37456	:douta	=	16'h	636f;
37457	:douta	=	16'h	638f;
37458	:douta	=	16'h	638f;
37459	:douta	=	16'h	6bb0;
37460	:douta	=	16'h	6b90;
37461	:douta	=	16'h	638f;
37462	:douta	=	16'h	6bb0;
37463	:douta	=	16'h	6bd0;
37464	:douta	=	16'h	6baf;
37465	:douta	=	16'h	636e;
37466	:douta	=	16'h	530d;
37467	:douta	=	16'h	9471;
37468	:douta	=	16'h	bd34;
37469	:douta	=	16'h	ad15;
37470	:douta	=	16'h	ad36;
37471	:douta	=	16'h	ad35;
37472	:douta	=	16'h	ad35;
37473	:douta	=	16'h	9cb5;
37474	:douta	=	16'h	9c94;
37475	:douta	=	16'h	94d5;
37476	:douta	=	16'h	8c73;
37477	:douta	=	16'h	7bd1;
37478	:douta	=	16'h	8432;
37479	:douta	=	16'h	7bd1;
37480	:douta	=	16'h	7bd1;
37481	:douta	=	16'h	6b6f;
37482	:douta	=	16'h	6b2e;
37483	:douta	=	16'h	630d;
37484	:douta	=	16'h	6acc;
37485	:douta	=	16'h	ac0e;
37486	:douta	=	16'h	d5b3;
37487	:douta	=	16'h	cd94;
37488	:douta	=	16'h	9c94;
37489	:douta	=	16'h	9475;
37490	:douta	=	16'h	acf5;
37491	:douta	=	16'h	9cd5;
37492	:douta	=	16'h	8453;
37493	:douta	=	16'h	8433;
37494	:douta	=	16'h	8433;
37495	:douta	=	16'h	7c12;
37496	:douta	=	16'h	632f;
37497	:douta	=	16'h	6b4f;
37498	:douta	=	16'h	632e;
37499	:douta	=	16'h	62ac;
37500	:douta	=	16'h	62cc;
37501	:douta	=	16'h	62ac;
37502	:douta	=	16'h	5229;
37503	:douta	=	16'h	72cb;
37504	:douta	=	16'h	52ef;
37505	:douta	=	16'h	5aac;
37506	:douta	=	16'h	9c31;
37507	:douta	=	16'h	8414;
37508	:douta	=	16'h	6b50;
37509	:douta	=	16'h	62cd;
37510	:douta	=	16'h	6b0d;
37511	:douta	=	16'h	5acc;
37512	:douta	=	16'h	62ac;
37513	:douta	=	16'h	5a8b;
37514	:douta	=	16'h	524b;
37515	:douta	=	16'h	4a2a;
37516	:douta	=	16'h	41e8;
37517	:douta	=	16'h	20e7;
37518	:douta	=	16'h	5249;
37519	:douta	=	16'h	ddf4;
37520	:douta	=	16'h	ee55;
37521	:douta	=	16'h	94d5;
37522	:douta	=	16'h	6bb2;
37523	:douta	=	16'h	8c53;
37524	:douta	=	16'h	9495;
37525	:douta	=	16'h	8c53;
37526	:douta	=	16'h	7c32;
37527	:douta	=	16'h	73f2;
37528	:douta	=	16'h	73b1;
37529	:douta	=	16'h	7350;
37530	:douta	=	16'h	632f;
37531	:douta	=	16'h	322c;
37532	:douta	=	16'h	424d;
37533	:douta	=	16'h	52ae;
37534	:douta	=	16'h	5aee;
37535	:douta	=	16'h	52ad;
37536	:douta	=	16'h	8bef;
37537	:douta	=	16'h	de15;
37538	:douta	=	16'h	ee97;
37539	:douta	=	16'h	eed8;
37540	:douta	=	16'h	eeb7;
37541	:douta	=	16'h	d616;
37542	:douta	=	16'h	de37;
37543	:douta	=	16'h	cdf6;
37544	:douta	=	16'h	b555;
37545	:douta	=	16'h	bd76;
37546	:douta	=	16'h	bd96;
37547	:douta	=	16'h	ad15;
37548	:douta	=	16'h	9494;
37549	:douta	=	16'h	a4b4;
37550	:douta	=	16'h	a515;
37551	:douta	=	16'h	9493;
37552	:douta	=	16'h	9473;
37553	:douta	=	16'h	9c93;
37554	:douta	=	16'h	8411;
37555	:douta	=	16'h	8412;
37556	:douta	=	16'h	7bf1;
37557	:douta	=	16'h	7c11;
37558	:douta	=	16'h	7c11;
37559	:douta	=	16'h	73b0;
37560	:douta	=	16'h	6b4f;
37561	:douta	=	16'h	7370;
37562	:douta	=	16'h	73b1;
37563	:douta	=	16'h	630d;
37564	:douta	=	16'h	5249;
37565	:douta	=	16'h	5a49;
37566	:douta	=	16'h	5a8a;
37567	:douta	=	16'h	5a69;
37568	:douta	=	16'h	5a28;
37569	:douta	=	16'h	ac8d;
37570	:douta	=	16'h	cd71;
37571	:douta	=	16'h	e655;
37572	:douta	=	16'h	d5d3;
37573	:douta	=	16'h	bd54;
37574	:douta	=	16'h	ad34;
37575	:douta	=	16'h	ad14;
37576	:douta	=	16'h	9d15;
37577	:douta	=	16'h	9cf5;
37578	:douta	=	16'h	94d5;
37579	:douta	=	16'h	7c54;
37580	:douta	=	16'h	7c54;
37581	:douta	=	16'h	7434;
37582	:douta	=	16'h	7435;
37583	:douta	=	16'h	6392;
37584	:douta	=	16'h	4b10;
37585	:douta	=	16'h	4b10;
37586	:douta	=	16'h	42af;
37587	:douta	=	16'h	3a8e;
37588	:douta	=	16'h	29a9;
37589	:douta	=	16'h	2988;
37590	:douta	=	16'h	6b91;
37591	:douta	=	16'h	31a8;
37592	:douta	=	16'h	0883;
37593	:douta	=	16'h	10c4;
37594	:douta	=	16'h	0884;
37595	:douta	=	16'h	10c5;
37596	:douta	=	16'h	29a9;
37597	:douta	=	16'h	2168;
37598	:douta	=	16'h	6a24;
37599	:douta	=	16'h	8285;
37600	:douta	=	16'h	8285;
37601	:douta	=	16'h	7a64;
37602	:douta	=	16'h	7a84;
37603	:douta	=	16'h	7a65;
37604	:douta	=	16'h	7a44;
37605	:douta	=	16'h	7224;
37606	:douta	=	16'h	7224;
37607	:douta	=	16'h	7224;
37608	:douta	=	16'h	7225;
37609	:douta	=	16'h	6a25;
37610	:douta	=	16'h	6a24;
37611	:douta	=	16'h	6204;
37612	:douta	=	16'h	6205;
37613	:douta	=	16'h	61e4;
37614	:douta	=	16'h	61e4;
37615	:douta	=	16'h	61e5;
37616	:douta	=	16'h	61e5;
37617	:douta	=	16'h	61e5;
37618	:douta	=	16'h	59e4;
37619	:douta	=	16'h	59c5;
37620	:douta	=	16'h	51a5;
37621	:douta	=	16'h	5164;
37622	:douta	=	16'h	5144;
37623	:douta	=	16'h	4943;
37624	:douta	=	16'h	51a5;
37625	:douta	=	16'h	59e6;
37626	:douta	=	16'h	628a;
37627	:douta	=	16'h	62cb;
37628	:douta	=	16'h	736d;
37629	:douta	=	16'h	7bae;
37630	:douta	=	16'h	83f0;
37631	:douta	=	16'h	7c10;
37632	:douta	=	16'h	ed8c;
37633	:douta	=	16'h	ed6b;
37634	:douta	=	16'h	e54b;
37635	:douta	=	16'h	e54b;
37636	:douta	=	16'h	dd29;
37637	:douta	=	16'h	dd09;
37638	:douta	=	16'h	bc45;
37639	:douta	=	16'h	92c8;
37640	:douta	=	16'h	e656;
37641	:douta	=	16'h	d573;
37642	:douta	=	16'h	cd73;
37643	:douta	=	16'h	cd92;
37644	:douta	=	16'h	ddd4;
37645	:douta	=	16'h	f77a;
37646	:douta	=	16'h	e677;
37647	:douta	=	16'h	ddf6;
37648	:douta	=	16'h	8433;
37649	:douta	=	16'h	6bd3;
37650	:douta	=	16'h	7c55;
37651	:douta	=	16'h	84b7;
37652	:douta	=	16'h	8475;
37653	:douta	=	16'h	73b2;
37654	:douta	=	16'h	8496;
37655	:douta	=	16'h	8496;
37656	:douta	=	16'h	9d39;
37657	:douta	=	16'h	9579;
37658	:douta	=	16'h	29eb;
37659	:douta	=	16'h	326d;
37660	:douta	=	16'h	3a8e;
37661	:douta	=	16'h	3aae;
37662	:douta	=	16'h	328e;
37663	:douta	=	16'h	3aae;
37664	:douta	=	16'h	3a8e;
37665	:douta	=	16'h	3a8e;
37666	:douta	=	16'h	3aae;
37667	:douta	=	16'h	3a8d;
37668	:douta	=	16'h	21ca;
37669	:douta	=	16'h	21a9;
37670	:douta	=	16'h	29ea;
37671	:douta	=	16'h	29ea;
37672	:douta	=	16'h	29c9;
37673	:douta	=	16'h	2167;
37674	:douta	=	16'h	18e4;
37675	:douta	=	16'h	10a3;
37676	:douta	=	16'h	18c4;
37677	:douta	=	16'h	1905;
37678	:douta	=	16'h	2145;
37679	:douta	=	16'h	2967;
37680	:douta	=	16'h	31c9;
37681	:douta	=	16'h	39ea;
37682	:douta	=	16'h	422a;
37683	:douta	=	16'h	422a;
37684	:douta	=	16'h	4a4b;
37685	:douta	=	16'h	422a;
37686	:douta	=	16'h	422a;
37687	:douta	=	16'h	39ea;
37688	:douta	=	16'h	31c9;
37689	:douta	=	16'h	31a9;
37690	:douta	=	16'h	29a8;
37691	:douta	=	16'h	2146;
37692	:douta	=	16'h	1905;
37693	:douta	=	16'h	10e5;
37694	:douta	=	16'h	10e6;
37695	:douta	=	16'h	10e5;
37696	:douta	=	16'h	0883;
37697	:douta	=	16'h	10a4;
37698	:douta	=	16'h	3a4c;
37699	:douta	=	16'h	42ee;
37700	:douta	=	16'h	4aed;
37701	:douta	=	16'h	4b0d;
37702	:douta	=	16'h	532f;
37703	:douta	=	16'h	52ed;
37704	:douta	=	16'h	530d;
37705	:douta	=	16'h	5b4e;
37706	:douta	=	16'h	5b2e;
37707	:douta	=	16'h	5b0e;
37708	:douta	=	16'h	636f;
37709	:douta	=	16'h	6b90;
37710	:douta	=	16'h	636f;
37711	:douta	=	16'h	638f;
37712	:douta	=	16'h	6bb0;
37713	:douta	=	16'h	6bd0;
37714	:douta	=	16'h	6bd0;
37715	:douta	=	16'h	6bb0;
37716	:douta	=	16'h	636f;
37717	:douta	=	16'h	634e;
37718	:douta	=	16'h	6b8f;
37719	:douta	=	16'h	6bb0;
37720	:douta	=	16'h	636f;
37721	:douta	=	16'h	636e;
37722	:douta	=	16'h	5b4e;
37723	:douta	=	16'h	638f;
37724	:douta	=	16'h	636e;
37725	:douta	=	16'h	73af;
37726	:douta	=	16'h	8410;
37727	:douta	=	16'h	9cb3;
37728	:douta	=	16'h	9cb3;
37729	:douta	=	16'h	ad14;
37730	:douta	=	16'h	9493;
37731	:douta	=	16'h	9493;
37732	:douta	=	16'h	8c32;
37733	:douta	=	16'h	8412;
37734	:douta	=	16'h	83f1;
37735	:douta	=	16'h	7bf1;
37736	:douta	=	16'h	736f;
37737	:douta	=	16'h	526b;
37738	:douta	=	16'h	730d;
37739	:douta	=	16'h	93ee;
37740	:douta	=	16'h	f6d6;
37741	:douta	=	16'h	e655;
37742	:douta	=	16'h	ad15;
37743	:douta	=	16'h	acf5;
37744	:douta	=	16'h	94b6;
37745	:douta	=	16'h	8c95;
37746	:douta	=	16'h	8c74;
37747	:douta	=	16'h	8c95;
37748	:douta	=	16'h	7390;
37749	:douta	=	16'h	736f;
37750	:douta	=	16'h	7390;
37751	:douta	=	16'h	7b90;
37752	:douta	=	16'h	6b0d;
37753	:douta	=	16'h	5aab;
37754	:douta	=	16'h	628b;
37755	:douta	=	16'h	62cc;
37756	:douta	=	16'h	5a6b;
37757	:douta	=	16'h	62cb;
37758	:douta	=	16'h	b4d3;
37759	:douta	=	16'h	acd3;
37760	:douta	=	16'h	428d;
37761	:douta	=	16'h	4a2a;
37762	:douta	=	16'h	83d1;
37763	:douta	=	16'h	6b4f;
37764	:douta	=	16'h	6b2e;
37765	:douta	=	16'h	524a;
37766	:douta	=	16'h	41c8;
37767	:douta	=	16'h	2988;
37768	:douta	=	16'h	39e8;
37769	:douta	=	16'h	41e8;
37770	:douta	=	16'h	420a;
37771	:douta	=	16'h	2968;
37772	:douta	=	16'h	732d;
37773	:douta	=	16'h	d5b2;
37774	:douta	=	16'h	c574;
37775	:douta	=	16'h	bd13;
37776	:douta	=	16'h	acf5;
37777	:douta	=	16'h	7c13;
37778	:douta	=	16'h	6391;
37779	:douta	=	16'h	6370;
37780	:douta	=	16'h	8c74;
37781	:douta	=	16'h	83f2;
37782	:douta	=	16'h	6b70;
37783	:douta	=	16'h	6b2f;
37784	:douta	=	16'h	6b2e;
37785	:douta	=	16'h	62ed;
37786	:douta	=	16'h	6b0e;
37787	:douta	=	16'h	736f;
37788	:douta	=	16'h	6b4f;
37789	:douta	=	16'h	7bb0;
37790	:douta	=	16'h	a470;
37791	:douta	=	16'h	d5f4;
37792	:douta	=	16'h	eeb7;
37793	:douta	=	16'h	de77;
37794	:douta	=	16'h	e677;
37795	:douta	=	16'h	cdf7;
37796	:douta	=	16'h	b577;
37797	:douta	=	16'h	c5d7;
37798	:douta	=	16'h	c5d7;
37799	:douta	=	16'h	c5b6;
37800	:douta	=	16'h	bd96;
37801	:douta	=	16'h	ad56;
37802	:douta	=	16'h	b556;
37803	:douta	=	16'h	a515;
37804	:douta	=	16'h	8c74;
37805	:douta	=	16'h	7c34;
37806	:douta	=	16'h	8453;
37807	:douta	=	16'h	9472;
37808	:douta	=	16'h	9473;
37809	:douta	=	16'h	9473;
37810	:douta	=	16'h	8c73;
37811	:douta	=	16'h	8432;
37812	:douta	=	16'h	73b0;
37813	:douta	=	16'h	83f1;
37814	:douta	=	16'h	7c12;
37815	:douta	=	16'h	62ee;
37816	:douta	=	16'h	630d;
37817	:douta	=	16'h	6aeb;
37818	:douta	=	16'h	730b;
37819	:douta	=	16'h	a46f;
37820	:douta	=	16'h	d5d3;
37821	:douta	=	16'h	de13;
37822	:douta	=	16'h	de55;
37823	:douta	=	16'h	e634;
37824	:douta	=	16'h	e655;
37825	:douta	=	16'h	e655;
37826	:douta	=	16'h	de15;
37827	:douta	=	16'h	de34;
37828	:douta	=	16'h	de15;
37829	:douta	=	16'h	bd33;
37830	:douta	=	16'h	ad14;
37831	:douta	=	16'h	ad14;
37832	:douta	=	16'h	a4f5;
37833	:douta	=	16'h	9cf6;
37834	:douta	=	16'h	8cb5;
37835	:douta	=	16'h	7c34;
37836	:douta	=	16'h	7414;
37837	:douta	=	16'h	7455;
37838	:douta	=	16'h	7c75;
37839	:douta	=	16'h	63f4;
37840	:douta	=	16'h	5351;
37841	:douta	=	16'h	4b10;
37842	:douta	=	16'h	42cf;
37843	:douta	=	16'h	42ae;
37844	:douta	=	16'h	29aa;
37845	:douta	=	16'h	2989;
37846	:douta	=	16'h	0064;
37847	:douta	=	16'h	7c54;
37848	:douta	=	16'h	1927;
37849	:douta	=	16'h	1907;
37850	:douta	=	16'h	1906;
37851	:douta	=	16'h	18e5;
37852	:douta	=	16'h	1927;
37853	:douta	=	16'h	1949;
37854	:douta	=	16'h	8ac5;
37855	:douta	=	16'h	7aa5;
37856	:douta	=	16'h	8285;
37857	:douta	=	16'h	7a85;
37858	:douta	=	16'h	7a84;
37859	:douta	=	16'h	7a65;
37860	:douta	=	16'h	7a64;
37861	:douta	=	16'h	7a65;
37862	:douta	=	16'h	7224;
37863	:douta	=	16'h	7224;
37864	:douta	=	16'h	6a25;
37865	:douta	=	16'h	61e4;
37866	:douta	=	16'h	6a04;
37867	:douta	=	16'h	61c4;
37868	:douta	=	16'h	61a4;
37869	:douta	=	16'h	59a4;
37870	:douta	=	16'h	59a4;
37871	:douta	=	16'h	59e5;
37872	:douta	=	16'h	6a88;
37873	:douta	=	16'h	72ea;
37874	:douta	=	16'h	7b8c;
37875	:douta	=	16'h	8c51;
37876	:douta	=	16'h	9492;
37877	:douta	=	16'h	9d13;
37878	:douta	=	16'h	a534;
37879	:douta	=	16'h	9d13;
37880	:douta	=	16'h	94b1;
37881	:douta	=	16'h	8c50;
37882	:douta	=	16'h	83ee;
37883	:douta	=	16'h	7b8d;
37884	:douta	=	16'h	6aea;
37885	:douta	=	16'h	5a69;
37886	:douta	=	16'h	5a69;
37887	:douta	=	16'h	4a27;
37888	:douta	=	16'h	ed6b;
37889	:douta	=	16'h	e52a;
37890	:douta	=	16'h	e54a;
37891	:douta	=	16'h	e52a;
37892	:douta	=	16'h	dd2a;
37893	:douta	=	16'h	e52a;
37894	:douta	=	16'h	cc44;
37895	:douta	=	16'h	cd11;
37896	:douta	=	16'h	ddf4;
37897	:douta	=	16'h	d594;
37898	:douta	=	16'h	d594;
37899	:douta	=	16'h	ddb3;
37900	:douta	=	16'h	ee76;
37901	:douta	=	16'h	ff5b;
37902	:douta	=	16'h	de57;
37903	:douta	=	16'h	d5f6;
37904	:douta	=	16'h	73f2;
37905	:douta	=	16'h	7413;
37906	:douta	=	16'h	7c75;
37907	:douta	=	16'h	8496;
37908	:douta	=	16'h	73d2;
37909	:douta	=	16'h	8433;
37910	:douta	=	16'h	8cb6;
37911	:douta	=	16'h	8cd7;
37912	:douta	=	16'h	94f8;
37913	:douta	=	16'h	8496;
37914	:douta	=	16'h	29eb;
37915	:douta	=	16'h	322d;
37916	:douta	=	16'h	322c;
37917	:douta	=	16'h	3a8e;
37918	:douta	=	16'h	3aae;
37919	:douta	=	16'h	3a8e;
37920	:douta	=	16'h	3a8e;
37921	:douta	=	16'h	3a6d;
37922	:douta	=	16'h	3a4e;
37923	:douta	=	16'h	324d;
37924	:douta	=	16'h	2a0b;
37925	:douta	=	16'h	29ca;
37926	:douta	=	16'h	2168;
37927	:douta	=	16'h	29ea;
37928	:douta	=	16'h	29ca;
37929	:douta	=	16'h	10e5;
37930	:douta	=	16'h	18e5;
37931	:douta	=	16'h	10c3;
37932	:douta	=	16'h	18e5;
37933	:douta	=	16'h	2126;
37934	:douta	=	16'h	31c9;
37935	:douta	=	16'h	39ea;
37936	:douta	=	16'h	39e9;
37937	:douta	=	16'h	4a6c;
37938	:douta	=	16'h	52ac;
37939	:douta	=	16'h	62cd;
37940	:douta	=	16'h	62ed;
37941	:douta	=	16'h	6b0e;
37942	:douta	=	16'h	52ac;
37943	:douta	=	16'h	528c;
37944	:douta	=	16'h	4a8d;
37945	:douta	=	16'h	426d;
37946	:douta	=	16'h	3a2c;
37947	:douta	=	16'h	31ea;
37948	:douta	=	16'h	29a9;
37949	:douta	=	16'h	2168;
37950	:douta	=	16'h	1106;
37951	:douta	=	16'h	10c5;
37952	:douta	=	16'h	10e4;
37953	:douta	=	16'h	10a4;
37954	:douta	=	16'h	10a4;
37955	:douta	=	16'h	1946;
37956	:douta	=	16'h	3a8c;
37957	:douta	=	16'h	3a4c;
37958	:douta	=	16'h	4aad;
37959	:douta	=	16'h	426b;
37960	:douta	=	16'h	4aac;
37961	:douta	=	16'h	530d;
37962	:douta	=	16'h	5b2e;
37963	:douta	=	16'h	4acd;
37964	:douta	=	16'h	636f;
37965	:douta	=	16'h	636f;
37966	:douta	=	16'h	6b90;
37967	:douta	=	16'h	638f;
37968	:douta	=	16'h	638f;
37969	:douta	=	16'h	6bb0;
37970	:douta	=	16'h	6bd0;
37971	:douta	=	16'h	636f;
37972	:douta	=	16'h	6bb0;
37973	:douta	=	16'h	6b8f;
37974	:douta	=	16'h	6bb0;
37975	:douta	=	16'h	6bb0;
37976	:douta	=	16'h	6b8f;
37977	:douta	=	16'h	6bb0;
37978	:douta	=	16'h	638f;
37979	:douta	=	16'h	6baf;
37980	:douta	=	16'h	6baf;
37981	:douta	=	16'h	6b6e;
37982	:douta	=	16'h	6b6e;
37983	:douta	=	16'h	73cf;
37984	:douta	=	16'h	9452;
37985	:douta	=	16'h	9c73;
37986	:douta	=	16'h	a4d4;
37987	:douta	=	16'h	a4d4;
37988	:douta	=	16'h	9473;
37989	:douta	=	16'h	83f1;
37990	:douta	=	16'h	7bf1;
37991	:douta	=	16'h	736e;
37992	:douta	=	16'h	6b2d;
37993	:douta	=	16'h	62cd;
37994	:douta	=	16'h	d593;
37995	:douta	=	16'h	cd72;
37996	:douta	=	16'h	e655;
37997	:douta	=	16'h	c595;
37998	:douta	=	16'h	a4f5;
37999	:douta	=	16'h	ad36;
38000	:douta	=	16'h	94b6;
38001	:douta	=	16'h	94d6;
38002	:douta	=	16'h	9496;
38003	:douta	=	16'h	8c74;
38004	:douta	=	16'h	7bf1;
38005	:douta	=	16'h	7bd1;
38006	:douta	=	16'h	736f;
38007	:douta	=	16'h	738f;
38008	:douta	=	16'h	6b0e;
38009	:douta	=	16'h	62cc;
38010	:douta	=	16'h	6acc;
38011	:douta	=	16'h	524a;
38012	:douta	=	16'h	5a6b;
38013	:douta	=	16'h	a493;
38014	:douta	=	16'h	9c73;
38015	:douta	=	16'h	9453;
38016	:douta	=	16'h	4a8c;
38017	:douta	=	16'h	422b;
38018	:douta	=	16'h	83d0;
38019	:douta	=	16'h	62ed;
38020	:douta	=	16'h	62cc;
38021	:douta	=	16'h	62ab;
38022	:douta	=	16'h	5a6a;
38023	:douta	=	16'h	41c8;
38024	:douta	=	16'h	2147;
38025	:douta	=	16'h	2127;
38026	:douta	=	16'h	2966;
38027	:douta	=	16'h	422a;
38028	:douta	=	16'h	b4f4;
38029	:douta	=	16'h	bd74;
38030	:douta	=	16'h	94b4;
38031	:douta	=	16'h	ad15;
38032	:douta	=	16'h	a4f5;
38033	:douta	=	16'h	5b2f;
38034	:douta	=	16'h	7bf3;
38035	:douta	=	16'h	5b30;
38036	:douta	=	16'h	8412;
38037	:douta	=	16'h	7bf1;
38038	:douta	=	16'h	6b2f;
38039	:douta	=	16'h	6b2e;
38040	:douta	=	16'h	6b0e;
38041	:douta	=	16'h	5a8c;
38042	:douta	=	16'h	630e;
38043	:douta	=	16'h	5aee;
38044	:douta	=	16'h	acd2;
38045	:douta	=	16'h	acd1;
38046	:douta	=	16'h	e697;
38047	:douta	=	16'h	eed9;
38048	:douta	=	16'h	e698;
38049	:douta	=	16'h	de57;
38050	:douta	=	16'h	d616;
38051	:douta	=	16'h	c5f7;
38052	:douta	=	16'h	b577;
38053	:douta	=	16'h	b576;
38054	:douta	=	16'h	b597;
38055	:douta	=	16'h	b577;
38056	:douta	=	16'h	b577;
38057	:douta	=	16'h	ad36;
38058	:douta	=	16'h	bdb7;
38059	:douta	=	16'h	b597;
38060	:douta	=	16'h	94d5;
38061	:douta	=	16'h	7c33;
38062	:douta	=	16'h	7bf3;
38063	:douta	=	16'h	7c33;
38064	:douta	=	16'h	8c52;
38065	:douta	=	16'h	8c53;
38066	:douta	=	16'h	8432;
38067	:douta	=	16'h	8432;
38068	:douta	=	16'h	7bf2;
38069	:douta	=	16'h	7bb2;
38070	:douta	=	16'h	5acc;
38071	:douta	=	16'h	a46f;
38072	:douta	=	16'h	c511;
38073	:douta	=	16'h	c552;
38074	:douta	=	16'h	cd93;
38075	:douta	=	16'h	d5d2;
38076	:douta	=	16'h	e635;
38077	:douta	=	16'h	de35;
38078	:douta	=	16'h	de35;
38079	:douta	=	16'h	e676;
38080	:douta	=	16'h	e676;
38081	:douta	=	16'h	e636;
38082	:douta	=	16'h	de15;
38083	:douta	=	16'h	c594;
38084	:douta	=	16'h	c574;
38085	:douta	=	16'h	a514;
38086	:douta	=	16'h	a4f5;
38087	:douta	=	16'h	a515;
38088	:douta	=	16'h	a516;
38089	:douta	=	16'h	94f5;
38090	:douta	=	16'h	8c95;
38091	:douta	=	16'h	7c34;
38092	:douta	=	16'h	7434;
38093	:douta	=	16'h	7413;
38094	:douta	=	16'h	7c55;
38095	:douta	=	16'h	7414;
38096	:douta	=	16'h	63b3;
38097	:douta	=	16'h	4b10;
38098	:douta	=	16'h	5310;
38099	:douta	=	16'h	42cf;
38100	:douta	=	16'h	31ca;
38101	:douta	=	16'h	31ea;
38102	:douta	=	16'h	2988;
38103	:douta	=	16'h	5351;
38104	:douta	=	16'h	5b71;
38105	:douta	=	16'h	29a8;
38106	:douta	=	16'h	1906;
38107	:douta	=	16'h	1906;
38108	:douta	=	16'h	2167;
38109	:douta	=	16'h	1947;
38110	:douta	=	16'h	7a66;
38111	:douta	=	16'h	8285;
38112	:douta	=	16'h	8285;
38113	:douta	=	16'h	7a64;
38114	:douta	=	16'h	7a64;
38115	:douta	=	16'h	7a44;
38116	:douta	=	16'h	7244;
38117	:douta	=	16'h	7245;
38118	:douta	=	16'h	6a04;
38119	:douta	=	16'h	69e4;
38120	:douta	=	16'h	61c4;
38121	:douta	=	16'h	61c4;
38122	:douta	=	16'h	6205;
38123	:douta	=	16'h	6a66;
38124	:douta	=	16'h	72c8;
38125	:douta	=	16'h	836a;
38126	:douta	=	16'h	8c0e;
38127	:douta	=	16'h	944f;
38128	:douta	=	16'h	a513;
38129	:douta	=	16'h	ad54;
38130	:douta	=	16'h	ad53;
38131	:douta	=	16'h	a513;
38132	:douta	=	16'h	a4d2;
38133	:douta	=	16'h	8c2f;
38134	:douta	=	16'h	83ee;
38135	:douta	=	16'h	734b;
38136	:douta	=	16'h	62c9;
38137	:douta	=	16'h	6288;
38138	:douta	=	16'h	5207;
38139	:douta	=	16'h	4985;
38140	:douta	=	16'h	4164;
38141	:douta	=	16'h	4144;
38142	:douta	=	16'h	4124;
38143	:douta	=	16'h	3944;
38144	:douta	=	16'h	e528;
38145	:douta	=	16'h	e507;
38146	:douta	=	16'h	e507;
38147	:douta	=	16'h	e4e7;
38148	:douta	=	16'h	dd07;
38149	:douta	=	16'h	dcc6;
38150	:douta	=	16'h	ff1a;
38151	:douta	=	16'h	f73b;
38152	:douta	=	16'h	fed8;
38153	:douta	=	16'h	ee96;
38154	:douta	=	16'h	e635;
38155	:douta	=	16'h	ee56;
38156	:douta	=	16'h	ff5b;
38157	:douta	=	16'h	f6f8;
38158	:douta	=	16'h	e636;
38159	:douta	=	16'h	bd95;
38160	:douta	=	16'h	7bf3;
38161	:douta	=	16'h	8454;
38162	:douta	=	16'h	8c75;
38163	:douta	=	16'h	7c54;
38164	:douta	=	16'h	5b0e;
38165	:douta	=	16'h	8c75;
38166	:douta	=	16'h	8cd7;
38167	:douta	=	16'h	94f8;
38168	:douta	=	16'h	9518;
38169	:douta	=	16'h	3a8d;
38170	:douta	=	16'h	29ca;
38171	:douta	=	16'h	2a0c;
38172	:douta	=	16'h	326d;
38173	:douta	=	16'h	326d;
38174	:douta	=	16'h	324d;
38175	:douta	=	16'h	42af;
38176	:douta	=	16'h	3a8e;
38177	:douta	=	16'h	3a8e;
38178	:douta	=	16'h	328e;
38179	:douta	=	16'h	326d;
38180	:douta	=	16'h	1127;
38181	:douta	=	16'h	1967;
38182	:douta	=	16'h	1926;
38183	:douta	=	16'h	2147;
38184	:douta	=	16'h	29ca;
38185	:douta	=	16'h	18e5;
38186	:douta	=	16'h	29a9;
38187	:douta	=	16'h	2146;
38188	:douta	=	16'h	29a9;
38189	:douta	=	16'h	31ea;
38190	:douta	=	16'h	31e9;
38191	:douta	=	16'h	31c9;
38192	:douta	=	16'h	31c9;
38193	:douta	=	16'h	39ea;
38194	:douta	=	16'h	3a0a;
38195	:douta	=	16'h	424b;
38196	:douta	=	16'h	4a6c;
38197	:douta	=	16'h	4a8c;
38198	:douta	=	16'h	424b;
38199	:douta	=	16'h	424c;
38200	:douta	=	16'h	422c;
38201	:douta	=	16'h	426d;
38202	:douta	=	16'h	428e;
38203	:douta	=	16'h	4acf;
38204	:douta	=	16'h	4aae;
38205	:douta	=	16'h	3a4c;
38206	:douta	=	16'h	3a4c;
38207	:douta	=	16'h	420b;
38208	:douta	=	16'h	1906;
38209	:douta	=	16'h	10e5;
38210	:douta	=	16'h	10c4;
38211	:douta	=	16'h	10c5;
38212	:douta	=	16'h	0884;
38213	:douta	=	16'h	29c9;
38214	:douta	=	16'h	3a6b;
38215	:douta	=	16'h	4acd;
38216	:douta	=	16'h	530e;
38217	:douta	=	16'h	530d;
38218	:douta	=	16'h	52cd;
38219	:douta	=	16'h	530d;
38220	:douta	=	16'h	5b2e;
38221	:douta	=	16'h	5b4e;
38222	:douta	=	16'h	5b4e;
38223	:douta	=	16'h	5b4f;
38224	:douta	=	16'h	636f;
38225	:douta	=	16'h	636f;
38226	:douta	=	16'h	6b8f;
38227	:douta	=	16'h	6b8f;
38228	:douta	=	16'h	636f;
38229	:douta	=	16'h	634f;
38230	:douta	=	16'h	6b90;
38231	:douta	=	16'h	6bb0;
38232	:douta	=	16'h	6bb0;
38233	:douta	=	16'h	6bb0;
38234	:douta	=	16'h	6b8f;
38235	:douta	=	16'h	73d0;
38236	:douta	=	16'h	73d0;
38237	:douta	=	16'h	73cf;
38238	:douta	=	16'h	73d0;
38239	:douta	=	16'h	6b8f;
38240	:douta	=	16'h	73cf;
38241	:douta	=	16'h	73cf;
38242	:douta	=	16'h	6b6e;
38243	:douta	=	16'h	6b6d;
38244	:douta	=	16'h	6b8e;
38245	:douta	=	16'h	7bef;
38246	:douta	=	16'h	83ef;
38247	:douta	=	16'h	738e;
38248	:douta	=	16'h	8bcf;
38249	:douta	=	16'h	cd33;
38250	:douta	=	16'h	a4f5;
38251	:douta	=	16'h	94d5;
38252	:douta	=	16'h	ad35;
38253	:douta	=	16'h	a4f6;
38254	:douta	=	16'h	94b5;
38255	:douta	=	16'h	8c53;
38256	:douta	=	16'h	7c11;
38257	:douta	=	16'h	73b0;
38258	:douta	=	16'h	736f;
38259	:douta	=	16'h	7b90;
38260	:douta	=	16'h	736e;
38261	:douta	=	16'h	732e;
38262	:douta	=	16'h	736e;
38263	:douta	=	16'h	736e;
38264	:douta	=	16'h	736d;
38265	:douta	=	16'h	62ab;
38266	:douta	=	16'h	5a6b;
38267	:douta	=	16'h	acb2;
38268	:douta	=	16'h	b4f2;
38269	:douta	=	16'h	73f2;
38270	:douta	=	16'h	8c53;
38271	:douta	=	16'h	8433;
38272	:douta	=	16'h	52ed;
38273	:douta	=	16'h	3a0a;
38274	:douta	=	16'h	73b0;
38275	:douta	=	16'h	62ac;
38276	:douta	=	16'h	6acb;
38277	:douta	=	16'h	62ab;
38278	:douta	=	16'h	5a8a;
38279	:douta	=	16'h	6289;
38280	:douta	=	16'h	51e8;
38281	:douta	=	16'h	6aab;
38282	:douta	=	16'h	6bd3;
38283	:douta	=	16'h	7c34;
38284	:douta	=	16'h	9c94;
38285	:douta	=	16'h	a515;
38286	:douta	=	16'h	a4f5;
38287	:douta	=	16'h	8474;
38288	:douta	=	16'h	8454;
38289	:douta	=	16'h	632f;
38290	:douta	=	16'h	426d;
38291	:douta	=	16'h	52ae;
38292	:douta	=	16'h	6b6f;
38293	:douta	=	16'h	736f;
38294	:douta	=	16'h	736e;
38295	:douta	=	16'h	62ed;
38296	:douta	=	16'h	5a8d;
38297	:douta	=	16'h	4a6c;
38298	:douta	=	16'h	5a6b;
38299	:douta	=	16'h	de35;
38300	:douta	=	16'h	c574;
38301	:douta	=	16'h	de56;
38302	:douta	=	16'h	e677;
38303	:douta	=	16'h	de56;
38304	:douta	=	16'h	d5f6;
38305	:douta	=	16'h	c5b6;
38306	:douta	=	16'h	bd96;
38307	:douta	=	16'h	b577;
38308	:douta	=	16'h	ad57;
38309	:douta	=	16'h	8c94;
38310	:douta	=	16'h	a516;
38311	:douta	=	16'h	9d16;
38312	:douta	=	16'h	a556;
38313	:douta	=	16'h	a557;
38314	:douta	=	16'h	9d16;
38315	:douta	=	16'h	9494;
38316	:douta	=	16'h	9474;
38317	:douta	=	16'h	8432;
38318	:douta	=	16'h	7c12;
38319	:douta	=	16'h	6b90;
38320	:douta	=	16'h	6b90;
38321	:douta	=	16'h	6b70;
38322	:douta	=	16'h	5aed;
38323	:douta	=	16'h	524a;
38324	:douta	=	16'h	5228;
38325	:douta	=	16'h	62c9;
38326	:douta	=	16'h	7b4c;
38327	:douta	=	16'h	49e7;
38328	:douta	=	16'h	5208;
38329	:douta	=	16'h	ac90;
38330	:douta	=	16'h	bd13;
38331	:douta	=	16'h	bd12;
38332	:douta	=	16'h	ee95;
38333	:douta	=	16'h	e676;
38334	:douta	=	16'h	d5d4;
38335	:douta	=	16'h	c574;
38336	:douta	=	16'h	acf3;
38337	:douta	=	16'h	bd34;
38338	:douta	=	16'h	ad14;
38339	:douta	=	16'h	a4d5;
38340	:douta	=	16'h	9cd5;
38341	:douta	=	16'h	9cd5;
38342	:douta	=	16'h	94d5;
38343	:douta	=	16'h	94d5;
38344	:douta	=	16'h	8c74;
38345	:douta	=	16'h	8c75;
38346	:douta	=	16'h	8454;
38347	:douta	=	16'h	7433;
38348	:douta	=	16'h	7413;
38349	:douta	=	16'h	73f3;
38350	:douta	=	16'h	6bd3;
38351	:douta	=	16'h	7434;
38352	:douta	=	16'h	63d3;
38353	:douta	=	16'h	4b10;
38354	:douta	=	16'h	4acf;
38355	:douta	=	16'h	29eb;
38356	:douta	=	16'h	636f;
38357	:douta	=	16'h	5b0f;
38358	:douta	=	16'h	324c;
38359	:douta	=	16'h	4b0f;
38360	:douta	=	16'h	42ad;
38361	:douta	=	16'h	31ea;
38362	:douta	=	16'h	2126;
38363	:douta	=	16'h	2127;
38364	:douta	=	16'h	2106;
38365	:douta	=	16'h	10e5;
38366	:douta	=	16'h	6289;
38367	:douta	=	16'h	7a24;
38368	:douta	=	16'h	7244;
38369	:douta	=	16'h	7a86;
38370	:douta	=	16'h	82c7;
38371	:douta	=	16'h	936a;
38372	:douta	=	16'h	9c0c;
38373	:douta	=	16'h	a44d;
38374	:douta	=	16'h	b510;
38375	:douta	=	16'h	bd51;
38376	:douta	=	16'h	c5b2;
38377	:douta	=	16'h	c592;
38378	:douta	=	16'h	bd51;
38379	:douta	=	16'h	ad0f;
38380	:douta	=	16'h	a4cf;
38381	:douta	=	16'h	942d;
38382	:douta	=	16'h	838c;
38383	:douta	=	16'h	7b4a;
38384	:douta	=	16'h	6aa8;
38385	:douta	=	16'h	6267;
38386	:douta	=	16'h	5a05;
38387	:douta	=	16'h	5184;
38388	:douta	=	16'h	4964;
38389	:douta	=	16'h	5164;
38390	:douta	=	16'h	4964;
38391	:douta	=	16'h	51a5;
38392	:douta	=	16'h	4965;
38393	:douta	=	16'h	5185;
38394	:douta	=	16'h	4985;
38395	:douta	=	16'h	4985;
38396	:douta	=	16'h	4985;
38397	:douta	=	16'h	49a5;
38398	:douta	=	16'h	49a5;
38399	:douta	=	16'h	4185;
38400	:douta	=	16'h	e506;
38401	:douta	=	16'h	e4e6;
38402	:douta	=	16'h	dd06;
38403	:douta	=	16'h	e4e6;
38404	:douta	=	16'h	dce6;
38405	:douta	=	16'h	d461;
38406	:douta	=	16'h	ff7d;
38407	:douta	=	16'h	f6f8;
38408	:douta	=	16'h	ff39;
38409	:douta	=	16'h	eeb7;
38410	:douta	=	16'h	e676;
38411	:douta	=	16'h	eeb8;
38412	:douta	=	16'h	ff7c;
38413	:douta	=	16'h	eeb7;
38414	:douta	=	16'h	de36;
38415	:douta	=	16'h	ad15;
38416	:douta	=	16'h	73f3;
38417	:douta	=	16'h	8455;
38418	:douta	=	16'h	8c76;
38419	:douta	=	16'h	73f2;
38420	:douta	=	16'h	5aee;
38421	:douta	=	16'h	8cb6;
38422	:douta	=	16'h	9539;
38423	:douta	=	16'h	8cb7;
38424	:douta	=	16'h	84b6;
38425	:douta	=	16'h	29eb;
38426	:douta	=	16'h	29eb;
38427	:douta	=	16'h	322c;
38428	:douta	=	16'h	324d;
38429	:douta	=	16'h	324d;
38430	:douta	=	16'h	326e;
38431	:douta	=	16'h	3a8e;
38432	:douta	=	16'h	3aaf;
38433	:douta	=	16'h	324d;
38434	:douta	=	16'h	326d;
38435	:douta	=	16'h	3a6e;
38436	:douta	=	16'h	1927;
38437	:douta	=	16'h	2168;
38438	:douta	=	16'h	1926;
38439	:douta	=	16'h	1947;
38440	:douta	=	16'h	2189;
38441	:douta	=	16'h	2127;
38442	:douta	=	16'h	29a9;
38443	:douta	=	16'h	2168;
38444	:douta	=	16'h	31ca;
38445	:douta	=	16'h	320a;
38446	:douta	=	16'h	31c9;
38447	:douta	=	16'h	31a8;
38448	:douta	=	16'h	29a8;
38449	:douta	=	16'h	39e9;
38450	:douta	=	16'h	3a0a;
38451	:douta	=	16'h	422a;
38452	:douta	=	16'h	424b;
38453	:douta	=	16'h	422b;
38454	:douta	=	16'h	3a0a;
38455	:douta	=	16'h	3a0a;
38456	:douta	=	16'h	3a2b;
38457	:douta	=	16'h	424c;
38458	:douta	=	16'h	424c;
38459	:douta	=	16'h	39eb;
38460	:douta	=	16'h	31eb;
38461	:douta	=	16'h	3a2b;
38462	:douta	=	16'h	3a2b;
38463	:douta	=	16'h	3a2b;
38464	:douta	=	16'h	3a0a;
38465	:douta	=	16'h	2988;
38466	:douta	=	16'h	18e5;
38467	:douta	=	16'h	1084;
38468	:douta	=	16'h	10a4;
38469	:douta	=	16'h	18e5;
38470	:douta	=	16'h	31c9;
38471	:douta	=	16'h	4aac;
38472	:douta	=	16'h	4aac;
38473	:douta	=	16'h	530d;
38474	:douta	=	16'h	4acd;
38475	:douta	=	16'h	52ed;
38476	:douta	=	16'h	530d;
38477	:douta	=	16'h	530d;
38478	:douta	=	16'h	5b2e;
38479	:douta	=	16'h	5b4e;
38480	:douta	=	16'h	5b2e;
38481	:douta	=	16'h	5b4e;
38482	:douta	=	16'h	636f;
38483	:douta	=	16'h	5b4e;
38484	:douta	=	16'h	5b4e;
38485	:douta	=	16'h	636f;
38486	:douta	=	16'h	636f;
38487	:douta	=	16'h	636f;
38488	:douta	=	16'h	6b90;
38489	:douta	=	16'h	6b90;
38490	:douta	=	16'h	6bb0;
38491	:douta	=	16'h	73d0;
38492	:douta	=	16'h	6baf;
38493	:douta	=	16'h	738f;
38494	:douta	=	16'h	73af;
38495	:douta	=	16'h	73cf;
38496	:douta	=	16'h	6b8f;
38497	:douta	=	16'h	73af;
38498	:douta	=	16'h	6b8f;
38499	:douta	=	16'h	6b8e;
38500	:douta	=	16'h	7baf;
38501	:douta	=	16'h	738f;
38502	:douta	=	16'h	7bcf;
38503	:douta	=	16'h	6b4d;
38504	:douta	=	16'h	5aeb;
38505	:douta	=	16'h	83ae;
38506	:douta	=	16'h	9c92;
38507	:douta	=	16'h	a4b4;
38508	:douta	=	16'h	a4f5;
38509	:douta	=	16'h	9cb4;
38510	:douta	=	16'h	9453;
38511	:douta	=	16'h	8412;
38512	:douta	=	16'h	83f1;
38513	:douta	=	16'h	7bd1;
38514	:douta	=	16'h	7b8f;
38515	:douta	=	16'h	734e;
38516	:douta	=	16'h	7b6e;
38517	:douta	=	16'h	734d;
38518	:douta	=	16'h	734d;
38519	:douta	=	16'h	732d;
38520	:douta	=	16'h	6acb;
38521	:douta	=	16'h	7b2b;
38522	:douta	=	16'h	a451;
38523	:douta	=	16'h	bd13;
38524	:douta	=	16'h	acd3;
38525	:douta	=	16'h	7bf2;
38526	:douta	=	16'h	8433;
38527	:douta	=	16'h	73b1;
38528	:douta	=	16'h	62ed;
38529	:douta	=	16'h	4a2b;
38530	:douta	=	16'h	7bf1;
38531	:douta	=	16'h	62cc;
38532	:douta	=	16'h	62aa;
38533	:douta	=	16'h	5a8a;
38534	:douta	=	16'h	628a;
38535	:douta	=	16'h	49c7;
38536	:douta	=	16'h	838e;
38537	:douta	=	16'h	9495;
38538	:douta	=	16'h	6b71;
38539	:douta	=	16'h	8c74;
38540	:douta	=	16'h	acf5;
38541	:douta	=	16'h	9d15;
38542	:douta	=	16'h	9cd5;
38543	:douta	=	16'h	8412;
38544	:douta	=	16'h	7bf2;
38545	:douta	=	16'h	7390;
38546	:douta	=	16'h	4aad;
38547	:douta	=	16'h	424c;
38548	:douta	=	16'h	3a4c;
38549	:douta	=	16'h	4a8d;
38550	:douta	=	16'h	62ed;
38551	:douta	=	16'h	4a6b;
38552	:douta	=	16'h	5aad;
38553	:douta	=	16'h	5aac;
38554	:douta	=	16'h	b4b2;
38555	:douta	=	16'h	f6d8;
38556	:douta	=	16'h	cdb5;
38557	:douta	=	16'h	cdf5;
38558	:douta	=	16'h	de56;
38559	:douta	=	16'h	cdf6;
38560	:douta	=	16'h	c5b6;
38561	:douta	=	16'h	b576;
38562	:douta	=	16'h	ad36;
38563	:douta	=	16'h	a4f5;
38564	:douta	=	16'h	9cf5;
38565	:douta	=	16'h	8c95;
38566	:douta	=	16'h	9494;
38567	:douta	=	16'h	9cf5;
38568	:douta	=	16'h	9cd6;
38569	:douta	=	16'h	94b5;
38570	:douta	=	16'h	9cf6;
38571	:douta	=	16'h	94b5;
38572	:douta	=	16'h	8453;
38573	:douta	=	16'h	7c11;
38574	:douta	=	16'h	7bf2;
38575	:douta	=	16'h	6b90;
38576	:douta	=	16'h	6b90;
38577	:douta	=	16'h	52ac;
38578	:douta	=	16'h	62aa;
38579	:douta	=	16'h	836c;
38580	:douta	=	16'h	a44e;
38581	:douta	=	16'h	bd30;
38582	:douta	=	16'h	c551;
38583	:douta	=	16'h	b4d0;
38584	:douta	=	16'h	834c;
38585	:douta	=	16'h	72ca;
38586	:douta	=	16'h	ac50;
38587	:douta	=	16'h	acf1;
38588	:douta	=	16'h	cd93;
38589	:douta	=	16'h	e655;
38590	:douta	=	16'h	de34;
38591	:douta	=	16'h	e655;
38592	:douta	=	16'h	b513;
38593	:douta	=	16'h	9c93;
38594	:douta	=	16'h	9cb3;
38595	:douta	=	16'h	a4f5;
38596	:douta	=	16'h	a515;
38597	:douta	=	16'h	94b5;
38598	:douta	=	16'h	8c94;
38599	:douta	=	16'h	8c95;
38600	:douta	=	16'h	8474;
38601	:douta	=	16'h	8454;
38602	:douta	=	16'h	7c13;
38603	:douta	=	16'h	7c34;
38604	:douta	=	16'h	7413;
38605	:douta	=	16'h	73f3;
38606	:douta	=	16'h	6bb3;
38607	:douta	=	16'h	63b2;
38608	:douta	=	16'h	63b3;
38609	:douta	=	16'h	63b3;
38610	:douta	=	16'h	5331;
38611	:douta	=	16'h	4aaf;
38612	:douta	=	16'h	428d;
38613	:douta	=	16'h	7bf1;
38614	:douta	=	16'h	320b;
38615	:douta	=	16'h	6c13;
38616	:douta	=	16'h	428d;
38617	:douta	=	16'h	6371;
38618	:douta	=	16'h	1906;
38619	:douta	=	16'h	1906;
38620	:douta	=	16'h	2127;
38621	:douta	=	16'h	2147;
38622	:douta	=	16'h	1927;
38623	:douta	=	16'h	9beb;
38624	:douta	=	16'h	9c0b;
38625	:douta	=	16'h	bd30;
38626	:douta	=	16'h	c572;
38627	:douta	=	16'h	ce13;
38628	:douta	=	16'h	d612;
38629	:douta	=	16'h	ce12;
38630	:douta	=	16'h	c5b1;
38631	:douta	=	16'h	bd70;
38632	:douta	=	16'h	a4ad;
38633	:douta	=	16'h	940c;
38634	:douta	=	16'h	8bab;
38635	:douta	=	16'h	7b09;
38636	:douta	=	16'h	72c8;
38637	:douta	=	16'h	6246;
38638	:douta	=	16'h	59c5;
38639	:douta	=	16'h	51a4;
38640	:douta	=	16'h	59a5;
38641	:douta	=	16'h	5184;
38642	:douta	=	16'h	51a5;
38643	:douta	=	16'h	59c5;
38644	:douta	=	16'h	51c5;
38645	:douta	=	16'h	51c5;
38646	:douta	=	16'h	51c5;
38647	:douta	=	16'h	51c5;
38648	:douta	=	16'h	4985;
38649	:douta	=	16'h	4965;
38650	:douta	=	16'h	4985;
38651	:douta	=	16'h	4985;
38652	:douta	=	16'h	4985;
38653	:douta	=	16'h	49a5;
38654	:douta	=	16'h	4986;
38655	:douta	=	16'h	4985;
38656	:douta	=	16'h	dca3;
38657	:douta	=	16'h	d484;
38658	:douta	=	16'h	d4a3;
38659	:douta	=	16'h	d484;
38660	:douta	=	16'h	cc20;
38661	:douta	=	16'h	ee55;
38662	:douta	=	16'h	f6f8;
38663	:douta	=	16'h	ff3a;
38664	:douta	=	16'h	ff3a;
38665	:douta	=	16'h	eeb8;
38666	:douta	=	16'h	eeb8;
38667	:douta	=	16'h	ff3a;
38668	:douta	=	16'h	ff9c;
38669	:douta	=	16'h	ee98;
38670	:douta	=	16'h	b555;
38671	:douta	=	16'h	8433;
38672	:douta	=	16'h	8455;
38673	:douta	=	16'h	8c75;
38674	:douta	=	16'h	8c95;
38675	:douta	=	16'h	6b2f;
38676	:douta	=	16'h	7b91;
38677	:douta	=	16'h	8496;
38678	:douta	=	16'h	8c76;
38679	:douta	=	16'h	9518;
38680	:douta	=	16'h	5330;
38681	:douta	=	16'h	08e6;
38682	:douta	=	16'h	21a9;
38683	:douta	=	16'h	21ca;
38684	:douta	=	16'h	2a2c;
38685	:douta	=	16'h	324d;
38686	:douta	=	16'h	324c;
38687	:douta	=	16'h	3a6d;
38688	:douta	=	16'h	322c;
38689	:douta	=	16'h	324d;
38690	:douta	=	16'h	3a4d;
38691	:douta	=	16'h	42af;
38692	:douta	=	16'h	1127;
38693	:douta	=	16'h	1948;
38694	:douta	=	16'h	1968;
38695	:douta	=	16'h	1947;
38696	:douta	=	16'h	2147;
38697	:douta	=	16'h	18e5;
38698	:douta	=	16'h	1926;
38699	:douta	=	16'h	1927;
38700	:douta	=	16'h	31c9;
38701	:douta	=	16'h	29a8;
38702	:douta	=	16'h	2988;
38703	:douta	=	16'h	31c9;
38704	:douta	=	16'h	39ea;
38705	:douta	=	16'h	422c;
38706	:douta	=	16'h	424c;
38707	:douta	=	16'h	426c;
38708	:douta	=	16'h	424c;
38709	:douta	=	16'h	424c;
38710	:douta	=	16'h	426c;
38711	:douta	=	16'h	4a8c;
38712	:douta	=	16'h	4a8d;
38713	:douta	=	16'h	426c;
38714	:douta	=	16'h	3a2b;
38715	:douta	=	16'h	424c;
38716	:douta	=	16'h	3a2b;
38717	:douta	=	16'h	39eb;
38718	:douta	=	16'h	31ca;
38719	:douta	=	16'h	31c9;
38720	:douta	=	16'h	3189;
38721	:douta	=	16'h	31a9;
38722	:douta	=	16'h	422a;
38723	:douta	=	16'h	29a8;
38724	:douta	=	16'h	1084;
38725	:douta	=	16'h	10a4;
38726	:douta	=	16'h	1906;
38727	:douta	=	16'h	320a;
38728	:douta	=	16'h	3a2b;
38729	:douta	=	16'h	52cd;
38730	:douta	=	16'h	4acc;
38731	:douta	=	16'h	52cd;
38732	:douta	=	16'h	4acd;
38733	:douta	=	16'h	4acd;
38734	:douta	=	16'h	52ed;
38735	:douta	=	16'h	5b2e;
38736	:douta	=	16'h	5b2e;
38737	:douta	=	16'h	530e;
38738	:douta	=	16'h	5b4e;
38739	:douta	=	16'h	5b2e;
38740	:douta	=	16'h	634f;
38741	:douta	=	16'h	634e;
38742	:douta	=	16'h	5b4e;
38743	:douta	=	16'h	636f;
38744	:douta	=	16'h	6baf;
38745	:douta	=	16'h	6b8f;
38746	:douta	=	16'h	6baf;
38747	:douta	=	16'h	73f0;
38748	:douta	=	16'h	73af;
38749	:douta	=	16'h	6b6e;
38750	:douta	=	16'h	634d;
38751	:douta	=	16'h	634d;
38752	:douta	=	16'h	632d;
38753	:douta	=	16'h	632d;
38754	:douta	=	16'h	634e;
38755	:douta	=	16'h	6b6e;
38756	:douta	=	16'h	6b8e;
38757	:douta	=	16'h	738f;
38758	:douta	=	16'h	6b6e;
38759	:douta	=	16'h	7baf;
38760	:douta	=	16'h	7bae;
38761	:douta	=	16'h	7baf;
38762	:douta	=	16'h	736d;
38763	:douta	=	16'h	736d;
38764	:douta	=	16'h	83ef;
38765	:douta	=	16'h	8bef;
38766	:douta	=	16'h	8c0f;
38767	:douta	=	16'h	8bcf;
38768	:douta	=	16'h	8bf0;
38769	:douta	=	16'h	83af;
38770	:douta	=	16'h	838f;
38771	:douta	=	16'h	736d;
38772	:douta	=	16'h	732c;
38773	:douta	=	16'h	732c;
38774	:douta	=	16'h	730b;
38775	:douta	=	16'h	836d;
38776	:douta	=	16'h	a4b3;
38777	:douta	=	16'h	9c92;
38778	:douta	=	16'h	8412;
38779	:douta	=	16'h	8c32;
38780	:douta	=	16'h	7bf1;
38781	:douta	=	16'h	734e;
38782	:douta	=	16'h	734d;
38783	:douta	=	16'h	732d;
38784	:douta	=	16'h	6b2c;
38785	:douta	=	16'h	6aeb;
38786	:douta	=	16'h	6aab;
38787	:douta	=	16'h	6acb;
38788	:douta	=	16'h	62ab;
38789	:douta	=	16'h	6269;
38790	:douta	=	16'h	730b;
38791	:douta	=	16'h	c574;
38792	:douta	=	16'h	8413;
38793	:douta	=	16'h	7bf1;
38794	:douta	=	16'h	6b50;
38795	:douta	=	16'h	9495;
38796	:douta	=	16'h	a516;
38797	:douta	=	16'h	94b5;
38798	:douta	=	16'h	8453;
38799	:douta	=	16'h	7bf1;
38800	:douta	=	16'h	7bd1;
38801	:douta	=	16'h	7390;
38802	:douta	=	16'h	7390;
38803	:douta	=	16'h	734f;
38804	:douta	=	16'h	62cd;
38805	:douta	=	16'h	52ad;
38806	:douta	=	16'h	422b;
38807	:douta	=	16'h	b535;
38808	:douta	=	16'h	a493;
38809	:douta	=	16'h	de77;
38810	:douta	=	16'h	f6f8;
38811	:douta	=	16'h	d5f6;
38812	:douta	=	16'h	bd96;
38813	:douta	=	16'h	9cd5;
38814	:douta	=	16'h	a515;
38815	:douta	=	16'h	ad56;
38816	:douta	=	16'h	a516;
38817	:douta	=	16'h	94b5;
38818	:douta	=	16'h	8c74;
38819	:douta	=	16'h	7bf1;
38820	:douta	=	16'h	7bd1;
38821	:douta	=	16'h	8412;
38822	:douta	=	16'h	8c94;
38823	:douta	=	16'h	7bf2;
38824	:douta	=	16'h	8c94;
38825	:douta	=	16'h	94d5;
38826	:douta	=	16'h	7c33;
38827	:douta	=	16'h	7c12;
38828	:douta	=	16'h	8433;
38829	:douta	=	16'h	6b91;
38830	:douta	=	16'h	5aad;
38831	:douta	=	16'h	524a;
38832	:douta	=	16'h	5a69;
38833	:douta	=	16'h	cdb4;
38834	:douta	=	16'h	cd92;
38835	:douta	=	16'h	ddf4;
38836	:douta	=	16'h	de14;
38837	:douta	=	16'h	e656;
38838	:douta	=	16'h	e655;
38839	:douta	=	16'h	de35;
38840	:douta	=	16'h	e675;
38841	:douta	=	16'h	f6b7;
38842	:douta	=	16'h	d5f4;
38843	:douta	=	16'h	acd1;
38844	:douta	=	16'h	acb2;
38845	:douta	=	16'h	a451;
38846	:douta	=	16'h	acd4;
38847	:douta	=	16'h	acb4;
38848	:douta	=	16'h	b514;
38849	:douta	=	16'h	bd54;
38850	:douta	=	16'h	ad14;
38851	:douta	=	16'h	9cb4;
38852	:douta	=	16'h	9cb4;
38853	:douta	=	16'h	94b4;
38854	:douta	=	16'h	8c54;
38855	:douta	=	16'h	8453;
38856	:douta	=	16'h	73f1;
38857	:douta	=	16'h	73f2;
38858	:douta	=	16'h	73d2;
38859	:douta	=	16'h	73b2;
38860	:douta	=	16'h	6bb1;
38861	:douta	=	16'h	5b50;
38862	:douta	=	16'h	6371;
38863	:douta	=	16'h	5b51;
38864	:douta	=	16'h	6371;
38865	:douta	=	16'h	4aee;
38866	:douta	=	16'h	3a4c;
38867	:douta	=	16'h	6b2d;
38868	:douta	=	16'h	94b4;
38869	:douta	=	16'h	3a4c;
38870	:douta	=	16'h	5aed;
38871	:douta	=	16'h	52cc;
38872	:douta	=	16'h	3a4c;
38873	:douta	=	16'h	29ca;
38874	:douta	=	16'h	10a4;
38875	:douta	=	16'h	1926;
38876	:douta	=	16'h	1905;
38877	:douta	=	16'h	18e5;
38878	:douta	=	16'h	18c4;
38879	:douta	=	16'h	83cc;
38880	:douta	=	16'h	bced;
38881	:douta	=	16'h	9bca;
38882	:douta	=	16'h	936a;
38883	:douta	=	16'h	82c7;
38884	:douta	=	16'h	7265;
38885	:douta	=	16'h	7225;
38886	:douta	=	16'h	69e4;
38887	:douta	=	16'h	61c4;
38888	:douta	=	16'h	69e4;
38889	:douta	=	16'h	61e5;
38890	:douta	=	16'h	61e5;
38891	:douta	=	16'h	61e5;
38892	:douta	=	16'h	61e5;
38893	:douta	=	16'h	61e4;
38894	:douta	=	16'h	59e4;
38895	:douta	=	16'h	59e5;
38896	:douta	=	16'h	59c5;
38897	:douta	=	16'h	59e5;
38898	:douta	=	16'h	51c5;
38899	:douta	=	16'h	51a5;
38900	:douta	=	16'h	59c5;
38901	:douta	=	16'h	51a5;
38902	:douta	=	16'h	51a5;
38903	:douta	=	16'h	4985;
38904	:douta	=	16'h	49a5;
38905	:douta	=	16'h	4985;
38906	:douta	=	16'h	4985;
38907	:douta	=	16'h	49a5;
38908	:douta	=	16'h	4985;
38909	:douta	=	16'h	4985;
38910	:douta	=	16'h	4986;
38911	:douta	=	16'h	4186;
38912	:douta	=	16'h	cc01;
38913	:douta	=	16'h	cc21;
38914	:douta	=	16'h	d443;
38915	:douta	=	16'h	d462;
38916	:douta	=	16'h	dccb;
38917	:douta	=	16'h	ff7c;
38918	:douta	=	16'h	f6f9;
38919	:douta	=	16'h	ff5b;
38920	:douta	=	16'h	ff3a;
38921	:douta	=	16'h	f6d8;
38922	:douta	=	16'h	f6b8;
38923	:douta	=	16'h	ff7b;
38924	:douta	=	16'h	ff7b;
38925	:douta	=	16'h	ee98;
38926	:douta	=	16'h	9493;
38927	:douta	=	16'h	7c13;
38928	:douta	=	16'h	8475;
38929	:douta	=	16'h	94d5;
38930	:douta	=	16'h	8cb6;
38931	:douta	=	16'h	6b2e;
38932	:douta	=	16'h	8412;
38933	:douta	=	16'h	8c75;
38934	:douta	=	16'h	8cb6;
38935	:douta	=	16'h	94d7;
38936	:douta	=	16'h	322b;
38937	:douta	=	16'h	0884;
38938	:douta	=	16'h	2168;
38939	:douta	=	16'h	2189;
38940	:douta	=	16'h	2189;
38941	:douta	=	16'h	29eb;
38942	:douta	=	16'h	322c;
38943	:douta	=	16'h	3a8e;
38944	:douta	=	16'h	324d;
38945	:douta	=	16'h	2a0c;
38946	:douta	=	16'h	3a4e;
38947	:douta	=	16'h	328e;
38948	:douta	=	16'h	1968;
38949	:douta	=	16'h	1947;
38950	:douta	=	16'h	1947;
38951	:douta	=	16'h	2147;
38952	:douta	=	16'h	2147;
38953	:douta	=	16'h	1905;
38954	:douta	=	16'h	1905;
38955	:douta	=	16'h	10a5;
38956	:douta	=	16'h	31ca;
38957	:douta	=	16'h	31ea;
38958	:douta	=	16'h	2987;
38959	:douta	=	16'h	39e9;
38960	:douta	=	16'h	424b;
38961	:douta	=	16'h	426d;
38962	:douta	=	16'h	424c;
38963	:douta	=	16'h	426c;
38964	:douta	=	16'h	3a4c;
38965	:douta	=	16'h	3a2b;
38966	:douta	=	16'h	3a2c;
38967	:douta	=	16'h	3a2c;
38968	:douta	=	16'h	426c;
38969	:douta	=	16'h	4a8d;
38970	:douta	=	16'h	4ace;
38971	:douta	=	16'h	426c;
38972	:douta	=	16'h	426d;
38973	:douta	=	16'h	3a2b;
38974	:douta	=	16'h	426c;
38975	:douta	=	16'h	3a0a;
38976	:douta	=	16'h	3188;
38977	:douta	=	16'h	2967;
38978	:douta	=	16'h	39ea;
38979	:douta	=	16'h	422b;
38980	:douta	=	16'h	18e5;
38981	:douta	=	16'h	18e5;
38982	:douta	=	16'h	0883;
38983	:douta	=	16'h	31ca;
38984	:douta	=	16'h	3a2b;
38985	:douta	=	16'h	4aac;
38986	:douta	=	16'h	4acd;
38987	:douta	=	16'h	52ed;
38988	:douta	=	16'h	52ed;
38989	:douta	=	16'h	530d;
38990	:douta	=	16'h	530d;
38991	:douta	=	16'h	530e;
38992	:douta	=	16'h	530d;
38993	:douta	=	16'h	5b2e;
38994	:douta	=	16'h	5b2e;
38995	:douta	=	16'h	5b2e;
38996	:douta	=	16'h	5b4e;
38997	:douta	=	16'h	634e;
38998	:douta	=	16'h	5b0d;
38999	:douta	=	16'h	5b4e;
39000	:douta	=	16'h	73d0;
39001	:douta	=	16'h	6b8f;
39002	:douta	=	16'h	6b90;
39003	:douta	=	16'h	6b8f;
39004	:douta	=	16'h	6b4e;
39005	:douta	=	16'h	5b0c;
39006	:douta	=	16'h	634d;
39007	:douta	=	16'h	634d;
39008	:douta	=	16'h	634e;
39009	:douta	=	16'h	6b6e;
39010	:douta	=	16'h	73af;
39011	:douta	=	16'h	73cf;
39012	:douta	=	16'h	73cf;
39013	:douta	=	16'h	6b8e;
39014	:douta	=	16'h	6b8e;
39015	:douta	=	16'h	738e;
39016	:douta	=	16'h	6b4d;
39017	:douta	=	16'h	738d;
39018	:douta	=	16'h	7bae;
39019	:douta	=	16'h	7bae;
39020	:douta	=	16'h	736d;
39021	:douta	=	16'h	7b6e;
39022	:douta	=	16'h	8c10;
39023	:douta	=	16'h	8bf0;
39024	:douta	=	16'h	83cf;
39025	:douta	=	16'h	8bef;
39026	:douta	=	16'h	8bef;
39027	:douta	=	16'h	8bcf;
39028	:douta	=	16'h	838e;
39029	:douta	=	16'h	838d;
39030	:douta	=	16'h	7b6d;
39031	:douta	=	16'h	8bef;
39032	:douta	=	16'h	a4b4;
39033	:douta	=	16'h	83f0;
39034	:douta	=	16'h	7baf;
39035	:douta	=	16'h	838f;
39036	:douta	=	16'h	7b6e;
39037	:douta	=	16'h	730c;
39038	:douta	=	16'h	6b0c;
39039	:douta	=	16'h	730c;
39040	:douta	=	16'h	6acc;
39041	:douta	=	16'h	6aca;
39042	:douta	=	16'h	6aaa;
39043	:douta	=	16'h	6aab;
39044	:douta	=	16'h	6a8a;
39045	:douta	=	16'h	bcd0;
39046	:douta	=	16'h	cd71;
39047	:douta	=	16'h	8412;
39048	:douta	=	16'h	7bb0;
39049	:douta	=	16'h	736f;
39050	:douta	=	16'h	62cd;
39051	:douta	=	16'h	7bb0;
39052	:douta	=	16'h	8411;
39053	:douta	=	16'h	83f1;
39054	:douta	=	16'h	83d1;
39055	:douta	=	16'h	7bf1;
39056	:douta	=	16'h	73b0;
39057	:douta	=	16'h	7390;
39058	:douta	=	16'h	734f;
39059	:douta	=	16'h	6b2e;
39060	:douta	=	16'h	62ed;
39061	:douta	=	16'h	5a8c;
39062	:douta	=	16'h	9c70;
39063	:douta	=	16'h	8c73;
39064	:douta	=	16'h	acb1;
39065	:douta	=	16'h	f6f9;
39066	:douta	=	16'h	de36;
39067	:douta	=	16'h	cdd6;
39068	:douta	=	16'h	c596;
39069	:douta	=	16'h	9cf6;
39070	:douta	=	16'h	a4f5;
39071	:douta	=	16'h	9cd5;
39072	:douta	=	16'h	9cd5;
39073	:douta	=	16'h	8c53;
39074	:douta	=	16'h	9494;
39075	:douta	=	16'h	7bf0;
39076	:douta	=	16'h	7bb0;
39077	:douta	=	16'h	7390;
39078	:douta	=	16'h	8c53;
39079	:douta	=	16'h	8433;
39080	:douta	=	16'h	73d1;
39081	:douta	=	16'h	8413;
39082	:douta	=	16'h	8453;
39083	:douta	=	16'h	7c12;
39084	:douta	=	16'h	6b4f;
39085	:douta	=	16'h	4a69;
39086	:douta	=	16'h	6aeb;
39087	:douta	=	16'h	bd73;
39088	:douta	=	16'h	c572;
39089	:douta	=	16'h	e656;
39090	:douta	=	16'h	e656;
39091	:douta	=	16'h	e676;
39092	:douta	=	16'h	d5f4;
39093	:douta	=	16'h	e676;
39094	:douta	=	16'h	cd93;
39095	:douta	=	16'h	d5d4;
39096	:douta	=	16'h	cd93;
39097	:douta	=	16'h	cd94;
39098	:douta	=	16'h	d5f4;
39099	:douta	=	16'h	e655;
39100	:douta	=	16'h	bd32;
39101	:douta	=	16'h	acd1;
39102	:douta	=	16'h	9c72;
39103	:douta	=	16'h	9c93;
39104	:douta	=	16'h	83f1;
39105	:douta	=	16'h	9473;
39106	:douta	=	16'h	9cb3;
39107	:douta	=	16'h	9c94;
39108	:douta	=	16'h	8c73;
39109	:douta	=	16'h	8432;
39110	:douta	=	16'h	8453;
39111	:douta	=	16'h	8454;
39112	:douta	=	16'h	7c12;
39113	:douta	=	16'h	73d2;
39114	:douta	=	16'h	6350;
39115	:douta	=	16'h	6b91;
39116	:douta	=	16'h	6b91;
39117	:douta	=	16'h	5b30;
39118	:douta	=	16'h	6371;
39119	:douta	=	16'h	6330;
39120	:douta	=	16'h	41e7;
39121	:douta	=	16'h	4a28;
39122	:douta	=	16'h	9c4e;
39123	:douta	=	16'h	bd72;
39124	:douta	=	16'h	4aae;
39125	:douta	=	16'h	632e;
39126	:douta	=	16'h	52cd;
39127	:douta	=	16'h	52cc;
39128	:douta	=	16'h	3a4c;
39129	:douta	=	16'h	18e5;
39130	:douta	=	16'h	10c4;
39131	:douta	=	16'h	0863;
39132	:douta	=	16'h	1083;
39133	:douta	=	16'h	10a4;
39134	:douta	=	16'h	1906;
39135	:douta	=	16'h	2127;
39136	:douta	=	16'h	7aa7;
39137	:douta	=	16'h	7204;
39138	:douta	=	16'h	7224;
39139	:douta	=	16'h	7224;
39140	:douta	=	16'h	7225;
39141	:douta	=	16'h	7225;
39142	:douta	=	16'h	7225;
39143	:douta	=	16'h	7225;
39144	:douta	=	16'h	6a25;
39145	:douta	=	16'h	6a25;
39146	:douta	=	16'h	6204;
39147	:douta	=	16'h	6205;
39148	:douta	=	16'h	61e5;
39149	:douta	=	16'h	61e5;
39150	:douta	=	16'h	61e5;
39151	:douta	=	16'h	59c5;
39152	:douta	=	16'h	59e5;
39153	:douta	=	16'h	59c5;
39154	:douta	=	16'h	59c5;
39155	:douta	=	16'h	51c5;
39156	:douta	=	16'h	51c5;
39157	:douta	=	16'h	51c5;
39158	:douta	=	16'h	51a5;
39159	:douta	=	16'h	51a5;
39160	:douta	=	16'h	49a5;
39161	:douta	=	16'h	49a6;
39162	:douta	=	16'h	4985;
39163	:douta	=	16'h	4985;
39164	:douta	=	16'h	4986;
39165	:douta	=	16'h	4986;
39166	:douta	=	16'h	41a5;
39167	:douta	=	16'h	4165;
39168	:douta	=	16'h	d56e;
39169	:douta	=	16'h	cd4c;
39170	:douta	=	16'h	9b22;
39171	:douta	=	16'h	aae0;
39172	:douta	=	16'h	ffbc;
39173	:douta	=	16'h	ff1a;
39174	:douta	=	16'h	ff3a;
39175	:douta	=	16'h	ff3b;
39176	:douta	=	16'h	ff3b;
39177	:douta	=	16'h	f6d8;
39178	:douta	=	16'h	f6d8;
39179	:douta	=	16'h	ff9c;
39180	:douta	=	16'h	f6f8;
39181	:douta	=	16'h	de17;
39182	:douta	=	16'h	8c74;
39183	:douta	=	16'h	8c34;
39184	:douta	=	16'h	8c95;
39185	:douta	=	16'h	8c95;
39186	:douta	=	16'h	8434;
39187	:douta	=	16'h	7bd2;
39188	:douta	=	16'h	8c54;
39189	:douta	=	16'h	94d6;
39190	:douta	=	16'h	8cb5;
39191	:douta	=	16'h	9d18;
39192	:douta	=	16'h	08c5;
39193	:douta	=	16'h	2147;
39194	:douta	=	16'h	1968;
39195	:douta	=	16'h	2189;
39196	:douta	=	16'h	21aa;
39197	:douta	=	16'h	29ca;
39198	:douta	=	16'h	21a9;
39199	:douta	=	16'h	21ca;
39200	:douta	=	16'h	322c;
39201	:douta	=	16'h	29ea;
39202	:douta	=	16'h	29ea;
39203	:douta	=	16'h	29ca;
39204	:douta	=	16'h	2189;
39205	:douta	=	16'h	2168;
39206	:douta	=	16'h	1947;
39207	:douta	=	16'h	1106;
39208	:douta	=	16'h	1947;
39209	:douta	=	16'h	2168;
39210	:douta	=	16'h	1105;
39211	:douta	=	16'h	2168;
39212	:douta	=	16'h	10e5;
39213	:douta	=	16'h	2147;
39214	:douta	=	16'h	2988;
39215	:douta	=	16'h	31a9;
39216	:douta	=	16'h	4a8c;
39217	:douta	=	16'h	428d;
39218	:douta	=	16'h	4a8d;
39219	:douta	=	16'h	3a0b;
39220	:douta	=	16'h	320a;
39221	:douta	=	16'h	4a6c;
39222	:douta	=	16'h	52ad;
39223	:douta	=	16'h	426c;
39224	:douta	=	16'h	3a2b;
39225	:douta	=	16'h	3a2b;
39226	:douta	=	16'h	3a2b;
39227	:douta	=	16'h	424c;
39228	:douta	=	16'h	424c;
39229	:douta	=	16'h	4a8d;
39230	:douta	=	16'h	424c;
39231	:douta	=	16'h	31c9;
39232	:douta	=	16'h	3a0a;
39233	:douta	=	16'h	31a8;
39234	:douta	=	16'h	31a8;
39235	:douta	=	16'h	2967;
39236	:douta	=	16'h	422b;
39237	:douta	=	16'h	2126;
39238	:douta	=	16'h	31c8;
39239	:douta	=	16'h	2167;
39240	:douta	=	16'h	3a4c;
39241	:douta	=	16'h	4aad;
39242	:douta	=	16'h	4aad;
39243	:douta	=	16'h	4aed;
39244	:douta	=	16'h	4aad;
39245	:douta	=	16'h	4aac;
39246	:douta	=	16'h	530d;
39247	:douta	=	16'h	530d;
39248	:douta	=	16'h	5b0e;
39249	:douta	=	16'h	530d;
39250	:douta	=	16'h	530d;
39251	:douta	=	16'h	4aac;
39252	:douta	=	16'h	4aab;
39253	:douta	=	16'h	4aac;
39254	:douta	=	16'h	5aed;
39255	:douta	=	16'h	5aed;
39256	:douta	=	16'h	4aac;
39257	:douta	=	16'h	634e;
39258	:douta	=	16'h	634e;
39259	:douta	=	16'h	6b8f;
39260	:douta	=	16'h	7bf1;
39261	:douta	=	16'h	73d0;
39262	:douta	=	16'h	73d0;
39263	:douta	=	16'h	6b8f;
39264	:douta	=	16'h	634d;
39265	:douta	=	16'h	632d;
39266	:douta	=	16'h	5acc;
39267	:douta	=	16'h	5acb;
39268	:douta	=	16'h	632d;
39269	:douta	=	16'h	6b2d;
39270	:douta	=	16'h	6b4d;
39271	:douta	=	16'h	6b6d;
39272	:douta	=	16'h	6b4d;
39273	:douta	=	16'h	6b4d;
39274	:douta	=	16'h	62eb;
39275	:douta	=	16'h	6aeb;
39276	:douta	=	16'h	736e;
39277	:douta	=	16'h	738e;
39278	:douta	=	16'h	736d;
39279	:douta	=	16'h	736e;
39280	:douta	=	16'h	738e;
39281	:douta	=	16'h	732d;
39282	:douta	=	16'h	732d;
39283	:douta	=	16'h	734d;
39284	:douta	=	16'h	7b6e;
39285	:douta	=	16'h	7b6e;
39286	:douta	=	16'h	83ae;
39287	:douta	=	16'h	7b4d;
39288	:douta	=	16'h	732d;
39289	:douta	=	16'h	7b8e;
39290	:douta	=	16'h	83ae;
39291	:douta	=	16'h	8bcf;
39292	:douta	=	16'h	8bcf;
39293	:douta	=	16'h	834d;
39294	:douta	=	16'h	7b2c;
39295	:douta	=	16'h	7b0b;
39296	:douta	=	16'h	832b;
39297	:douta	=	16'h	834b;
39298	:douta	=	16'h	8bae;
39299	:douta	=	16'h	9471;
39300	:douta	=	16'h	9451;
39301	:douta	=	16'h	836f;
39302	:douta	=	16'h	7b8f;
39303	:douta	=	16'h	734e;
39304	:douta	=	16'h	7bb0;
39305	:douta	=	16'h	7bb0;
39306	:douta	=	16'h	630d;
39307	:douta	=	16'h	630e;
39308	:douta	=	16'h	8c11;
39309	:douta	=	16'h	736f;
39310	:douta	=	16'h	734e;
39311	:douta	=	16'h	732d;
39312	:douta	=	16'h	732d;
39313	:douta	=	16'h	6aed;
39314	:douta	=	16'h	5a8b;
39315	:douta	=	16'h	734e;
39316	:douta	=	16'h	940e;
39317	:douta	=	16'h	d5d4;
39318	:douta	=	16'h	cdf8;
39319	:douta	=	16'h	b535;
39320	:douta	=	16'h	de56;
39321	:douta	=	16'h	c5b6;
39322	:douta	=	16'h	bd76;
39323	:douta	=	16'h	b557;
39324	:douta	=	16'h	9cf6;
39325	:douta	=	16'h	9cd6;
39326	:douta	=	16'h	7c13;
39327	:douta	=	16'h	8453;
39328	:douta	=	16'h	9493;
39329	:douta	=	16'h	7bf2;
39330	:douta	=	16'h	6b2f;
39331	:douta	=	16'h	6b70;
39332	:douta	=	16'h	7370;
39333	:douta	=	16'h	6b6f;
39334	:douta	=	16'h	6b2e;
39335	:douta	=	16'h	7370;
39336	:douta	=	16'h	734f;
39337	:douta	=	16'h	734f;
39338	:douta	=	16'h	4a28;
39339	:douta	=	16'h	49e8;
39340	:douta	=	16'h	9c6f;
39341	:douta	=	16'h	e615;
39342	:douta	=	16'h	e676;
39343	:douta	=	16'h	bd13;
39344	:douta	=	16'h	b4d3;
39345	:douta	=	16'h	e676;
39346	:douta	=	16'h	de36;
39347	:douta	=	16'h	de35;
39348	:douta	=	16'h	de15;
39349	:douta	=	16'h	cd93;
39350	:douta	=	16'h	acd3;
39351	:douta	=	16'h	acf4;
39352	:douta	=	16'h	acd3;
39353	:douta	=	16'h	8c52;
39354	:douta	=	16'h	8c32;
39355	:douta	=	16'h	8c12;
39356	:douta	=	16'h	9c72;
39357	:douta	=	16'h	a4b3;
39358	:douta	=	16'h	a4d4;
39359	:douta	=	16'h	9cb3;
39360	:douta	=	16'h	9453;
39361	:douta	=	16'h	8c73;
39362	:douta	=	16'h	8c52;
39363	:douta	=	16'h	83f1;
39364	:douta	=	16'h	73b0;
39365	:douta	=	16'h	7390;
39366	:douta	=	16'h	73b0;
39367	:douta	=	16'h	7390;
39368	:douta	=	16'h	7391;
39369	:douta	=	16'h	6b70;
39370	:douta	=	16'h	6b71;
39371	:douta	=	16'h	6bb2;
39372	:douta	=	16'h	6bb1;
39373	:douta	=	16'h	4a49;
39374	:douta	=	16'h	41c7;
39375	:douta	=	16'h	5a88;
39376	:douta	=	16'h	a48f;
39377	:douta	=	16'h	bd11;
39378	:douta	=	16'h	de14;
39379	:douta	=	16'h	9451;
39380	:douta	=	16'h	3a0a;
39381	:douta	=	16'h	630d;
39382	:douta	=	16'h	632d;
39383	:douta	=	16'h	5b4f;
39384	:douta	=	16'h	3a0a;
39385	:douta	=	16'h	29a8;
39386	:douta	=	16'h	18e5;
39387	:douta	=	16'h	52ad;
39388	:douta	=	16'h	1906;
39389	:douta	=	16'h	2147;
39390	:douta	=	16'h	2127;
39391	:douta	=	16'h	10c5;
39392	:douta	=	16'h	1926;
39393	:douta	=	16'h	8286;
39394	:douta	=	16'h	8286;
39395	:douta	=	16'h	7a45;
39396	:douta	=	16'h	7a45;
39397	:douta	=	16'h	7225;
39398	:douta	=	16'h	7225;
39399	:douta	=	16'h	7225;
39400	:douta	=	16'h	6a25;
39401	:douta	=	16'h	6a05;
39402	:douta	=	16'h	6a05;
39403	:douta	=	16'h	6205;
39404	:douta	=	16'h	61e4;
39405	:douta	=	16'h	61e5;
39406	:douta	=	16'h	59e5;
39407	:douta	=	16'h	59e5;
39408	:douta	=	16'h	59c5;
39409	:douta	=	16'h	59c5;
39410	:douta	=	16'h	51c5;
39411	:douta	=	16'h	51c5;
39412	:douta	=	16'h	51a5;
39413	:douta	=	16'h	51a5;
39414	:douta	=	16'h	51a5;
39415	:douta	=	16'h	51a5;
39416	:douta	=	16'h	49a5;
39417	:douta	=	16'h	49a6;
39418	:douta	=	16'h	4986;
39419	:douta	=	16'h	49a5;
39420	:douta	=	16'h	4165;
39421	:douta	=	16'h	4185;
39422	:douta	=	16'h	4185;
39423	:douta	=	16'h	4165;
39424	:douta	=	16'h	f718;
39425	:douta	=	16'h	ac8a;
39426	:douta	=	16'h	71a1;
39427	:douta	=	16'h	89e1;
39428	:douta	=	16'h	ffbd;
39429	:douta	=	16'h	f6f9;
39430	:douta	=	16'h	ff3b;
39431	:douta	=	16'h	ff3a;
39432	:douta	=	16'h	ff3a;
39433	:douta	=	16'h	f6d8;
39434	:douta	=	16'h	f6f8;
39435	:douta	=	16'h	ff9c;
39436	:douta	=	16'h	eeb7;
39437	:douta	=	16'h	c596;
39438	:douta	=	16'h	9494;
39439	:douta	=	16'h	8c53;
39440	:douta	=	16'h	8cb5;
39441	:douta	=	16'h	8cb5;
39442	:douta	=	16'h	8433;
39443	:douta	=	16'h	8c53;
39444	:douta	=	16'h	8c74;
39445	:douta	=	16'h	94b6;
39446	:douta	=	16'h	8cb5;
39447	:douta	=	16'h	8475;
39448	:douta	=	16'h	10e5;
39449	:douta	=	16'h	1926;
39450	:douta	=	16'h	2189;
39451	:douta	=	16'h	21aa;
39452	:douta	=	16'h	21a9;
39453	:douta	=	16'h	2168;
39454	:douta	=	16'h	1967;
39455	:douta	=	16'h	1126;
39456	:douta	=	16'h	1948;
39457	:douta	=	16'h	1127;
39458	:douta	=	16'h	1947;
39459	:douta	=	16'h	1968;
39460	:douta	=	16'h	2168;
39461	:douta	=	16'h	1948;
39462	:douta	=	16'h	1106;
39463	:douta	=	16'h	1948;
39464	:douta	=	16'h	2168;
39465	:douta	=	16'h	2189;
39466	:douta	=	16'h	1967;
39467	:douta	=	16'h	29a9;
39468	:douta	=	16'h	18e6;
39469	:douta	=	16'h	18e5;
39470	:douta	=	16'h	2168;
39471	:douta	=	16'h	29a9;
39472	:douta	=	16'h	31c9;
39473	:douta	=	16'h	4a6e;
39474	:douta	=	16'h	426d;
39475	:douta	=	16'h	31ea;
39476	:douta	=	16'h	31ea;
39477	:douta	=	16'h	422b;
39478	:douta	=	16'h	4a6c;
39479	:douta	=	16'h	424c;
39480	:douta	=	16'h	424c;
39481	:douta	=	16'h	422c;
39482	:douta	=	16'h	320b;
39483	:douta	=	16'h	3a0b;
39484	:douta	=	16'h	3a0b;
39485	:douta	=	16'h	3a4c;
39486	:douta	=	16'h	3a2c;
39487	:douta	=	16'h	39ea;
39488	:douta	=	16'h	420a;
39489	:douta	=	16'h	39ea;
39490	:douta	=	16'h	424a;
39491	:douta	=	16'h	2968;
39492	:douta	=	16'h	39e9;
39493	:douta	=	16'h	2147;
39494	:douta	=	16'h	2967;
39495	:douta	=	16'h	31ca;
39496	:douta	=	16'h	3a2b;
39497	:douta	=	16'h	4aad;
39498	:douta	=	16'h	4aad;
39499	:douta	=	16'h	4aed;
39500	:douta	=	16'h	4aad;
39501	:douta	=	16'h	4acd;
39502	:douta	=	16'h	4acd;
39503	:douta	=	16'h	530d;
39504	:douta	=	16'h	4aac;
39505	:douta	=	16'h	4acc;
39506	:douta	=	16'h	4aac;
39507	:douta	=	16'h	4aac;
39508	:douta	=	16'h	4aab;
39509	:douta	=	16'h	4aac;
39510	:douta	=	16'h	5b0d;
39511	:douta	=	16'h	632e;
39512	:douta	=	16'h	636e;
39513	:douta	=	16'h	6b8f;
39514	:douta	=	16'h	6b8f;
39515	:douta	=	16'h	6b6f;
39516	:douta	=	16'h	6b8f;
39517	:douta	=	16'h	634e;
39518	:douta	=	16'h	632e;
39519	:douta	=	16'h	634d;
39520	:douta	=	16'h	5acb;
39521	:douta	=	16'h	528a;
39522	:douta	=	16'h	62cb;
39523	:douta	=	16'h	62cb;
39524	:douta	=	16'h	62cb;
39525	:douta	=	16'h	630c;
39526	:douta	=	16'h	6b0c;
39527	:douta	=	16'h	62cb;
39528	:douta	=	16'h	630c;
39529	:douta	=	16'h	62ec;
39530	:douta	=	16'h	6aeb;
39531	:douta	=	16'h	62cb;
39532	:douta	=	16'h	6b0c;
39533	:douta	=	16'h	6b0c;
39534	:douta	=	16'h	630c;
39535	:douta	=	16'h	6b0c;
39536	:douta	=	16'h	6b2c;
39537	:douta	=	16'h	732d;
39538	:douta	=	16'h	6b0c;
39539	:douta	=	16'h	62cb;
39540	:douta	=	16'h	6b0b;
39541	:douta	=	16'h	6aeb;
39542	:douta	=	16'h	734c;
39543	:douta	=	16'h	6b0b;
39544	:douta	=	16'h	732c;
39545	:douta	=	16'h	734d;
39546	:douta	=	16'h	732d;
39547	:douta	=	16'h	83ef;
39548	:douta	=	16'h	9431;
39549	:douta	=	16'h	8bee;
39550	:douta	=	16'h	8bef;
39551	:douta	=	16'h	9430;
39552	:douta	=	16'h	9491;
39553	:douta	=	16'h	9492;
39554	:douta	=	16'h	8c50;
39555	:douta	=	16'h	b597;
39556	:douta	=	16'h	b5b6;
39557	:douta	=	16'h	8bf0;
39558	:douta	=	16'h	7baf;
39559	:douta	=	16'h	7b90;
39560	:douta	=	16'h	736f;
39561	:douta	=	16'h	734f;
39562	:douta	=	16'h	632e;
39563	:douta	=	16'h	6b2e;
39564	:douta	=	16'h	7b8e;
39565	:douta	=	16'h	7b6f;
39566	:douta	=	16'h	7baf;
39567	:douta	=	16'h	732e;
39568	:douta	=	16'h	732e;
39569	:douta	=	16'h	528c;
39570	:douta	=	16'h	b4b0;
39571	:douta	=	16'h	c571;
39572	:douta	=	16'h	e697;
39573	:douta	=	16'h	f6d8;
39574	:douta	=	16'h	9cf5;
39575	:douta	=	16'h	bd55;
39576	:douta	=	16'h	d616;
39577	:douta	=	16'h	bd96;
39578	:douta	=	16'h	ad57;
39579	:douta	=	16'h	9d16;
39580	:douta	=	16'h	8c94;
39581	:douta	=	16'h	8c53;
39582	:douta	=	16'h	8454;
39583	:douta	=	16'h	73f2;
39584	:douta	=	16'h	8432;
39585	:douta	=	16'h	8432;
39586	:douta	=	16'h	73b0;
39587	:douta	=	16'h	52cd;
39588	:douta	=	16'h	5aef;
39589	:douta	=	16'h	5acd;
39590	:douta	=	16'h	52ac;
39591	:douta	=	16'h	5aad;
39592	:douta	=	16'h	526a;
39593	:douta	=	16'h	4a29;
39594	:douta	=	16'h	730b;
39595	:douta	=	16'h	8bee;
39596	:douta	=	16'h	de13;
39597	:douta	=	16'h	e677;
39598	:douta	=	16'h	e697;
39599	:douta	=	16'h	bd54;
39600	:douta	=	16'h	bd34;
39601	:douta	=	16'h	c574;
39602	:douta	=	16'h	ddf5;
39603	:douta	=	16'h	cdb6;
39604	:douta	=	16'h	cdd4;
39605	:douta	=	16'h	c573;
39606	:douta	=	16'h	a4b4;
39607	:douta	=	16'h	9473;
39608	:douta	=	16'h	9452;
39609	:douta	=	16'h	9473;
39610	:douta	=	16'h	9432;
39611	:douta	=	16'h	7bd1;
39612	:douta	=	16'h	73b0;
39613	:douta	=	16'h	6b90;
39614	:douta	=	16'h	8411;
39615	:douta	=	16'h	8c53;
39616	:douta	=	16'h	8412;
39617	:douta	=	16'h	8c32;
39618	:douta	=	16'h	8c33;
39619	:douta	=	16'h	8c32;
39620	:douta	=	16'h	7bf1;
39621	:douta	=	16'h	7390;
39622	:douta	=	16'h	7390;
39623	:douta	=	16'h	7390;
39624	:douta	=	16'h	6b4f;
39625	:douta	=	16'h	630e;
39626	:douta	=	16'h	630e;
39627	:douta	=	16'h	526a;
39628	:douta	=	16'h	41c8;
39629	:douta	=	16'h	4a27;
39630	:douta	=	16'h	732b;
39631	:douta	=	16'h	ac6f;
39632	:douta	=	16'h	cdd2;
39633	:douta	=	16'h	de55;
39634	:douta	=	16'h	c573;
39635	:douta	=	16'h	9c52;
39636	:douta	=	16'h	6390;
39637	:douta	=	16'h	6b90;
39638	:douta	=	16'h	6b90;
39639	:douta	=	16'h	5b2f;
39640	:douta	=	16'h	29a9;
39641	:douta	=	16'h	31c9;
39642	:douta	=	16'h	18e5;
39643	:douta	=	16'h	1926;
39644	:douta	=	16'h	29a9;
39645	:douta	=	16'h	10e5;
39646	:douta	=	16'h	10e5;
39647	:douta	=	16'h	18e4;
39648	:douta	=	16'h	10e5;
39649	:douta	=	16'h	2104;
39650	:douta	=	16'h	8286;
39651	:douta	=	16'h	7a65;
39652	:douta	=	16'h	7a65;
39653	:douta	=	16'h	7245;
39654	:douta	=	16'h	7225;
39655	:douta	=	16'h	7245;
39656	:douta	=	16'h	6a04;
39657	:douta	=	16'h	6a05;
39658	:douta	=	16'h	61e5;
39659	:douta	=	16'h	6205;
39660	:douta	=	16'h	61e5;
39661	:douta	=	16'h	61e5;
39662	:douta	=	16'h	59c5;
39663	:douta	=	16'h	59e5;
39664	:douta	=	16'h	59c5;
39665	:douta	=	16'h	51a5;
39666	:douta	=	16'h	51c5;
39667	:douta	=	16'h	51a5;
39668	:douta	=	16'h	51c5;
39669	:douta	=	16'h	49a5;
39670	:douta	=	16'h	51a5;
39671	:douta	=	16'h	49a5;
39672	:douta	=	16'h	49a5;
39673	:douta	=	16'h	49a6;
39674	:douta	=	16'h	49a5;
39675	:douta	=	16'h	4185;
39676	:douta	=	16'h	4985;
39677	:douta	=	16'h	4185;
39678	:douta	=	16'h	4185;
39679	:douta	=	16'h	4165;
39680	:douta	=	16'h	e653;
39681	:douta	=	16'h	cd2b;
39682	:douta	=	16'h	cd6c;
39683	:douta	=	16'h	f6b7;
39684	:douta	=	16'h	f6f8;
39685	:douta	=	16'h	f6d8;
39686	:douta	=	16'h	ff5b;
39687	:douta	=	16'h	ff3a;
39688	:douta	=	16'h	f719;
39689	:douta	=	16'h	f6f9;
39690	:douta	=	16'h	ff5b;
39691	:douta	=	16'h	f718;
39692	:douta	=	16'h	e697;
39693	:douta	=	16'h	9cb4;
39694	:douta	=	16'h	8c53;
39695	:douta	=	16'h	8c94;
39696	:douta	=	16'h	94b6;
39697	:douta	=	16'h	8cb6;
39698	:douta	=	16'h	7bf2;
39699	:douta	=	16'h	8c74;
39700	:douta	=	16'h	94b6;
39701	:douta	=	16'h	94d6;
39702	:douta	=	16'h	94f7;
39703	:douta	=	16'h	31e9;
39704	:douta	=	16'h	10c3;
39705	:douta	=	16'h	18e4;
39706	:douta	=	16'h	18e4;
39707	:douta	=	16'h	18e5;
39708	:douta	=	16'h	2168;
39709	:douta	=	16'h	2168;
39710	:douta	=	16'h	1947;
39711	:douta	=	16'h	1926;
39712	:douta	=	16'h	1105;
39713	:douta	=	16'h	1906;
39714	:douta	=	16'h	1927;
39715	:douta	=	16'h	1967;
39716	:douta	=	16'h	1947;
39717	:douta	=	16'h	1947;
39718	:douta	=	16'h	1968;
39719	:douta	=	16'h	1148;
39720	:douta	=	16'h	1947;
39721	:douta	=	16'h	2189;
39722	:douta	=	16'h	2168;
39723	:douta	=	16'h	1906;
39724	:douta	=	16'h	29ca;
39725	:douta	=	16'h	29ca;
39726	:douta	=	16'h	1926;
39727	:douta	=	16'h	18e5;
39728	:douta	=	16'h	1927;
39729	:douta	=	16'h	31ea;
39730	:douta	=	16'h	3a0b;
39731	:douta	=	16'h	2148;
39732	:douta	=	16'h	2188;
39733	:douta	=	16'h	3a0a;
39734	:douta	=	16'h	6b2e;
39735	:douta	=	16'h	5b30;
39736	:douta	=	16'h	42f0;
39737	:douta	=	16'h	322c;
39738	:douta	=	16'h	31c9;
39739	:douta	=	16'h	2988;
39740	:douta	=	16'h	29a9;
39741	:douta	=	16'h	3a2b;
39742	:douta	=	16'h	3a0b;
39743	:douta	=	16'h	31a9;
39744	:douta	=	16'h	39a9;
39745	:douta	=	16'h	41ea;
39746	:douta	=	16'h	2967;
39747	:douta	=	16'h	31c9;
39748	:douta	=	16'h	31c9;
39749	:douta	=	16'h	31c8;
39750	:douta	=	16'h	2147;
39751	:douta	=	16'h	29ea;
39752	:douta	=	16'h	320a;
39753	:douta	=	16'h	3a6b;
39754	:douta	=	16'h	428c;
39755	:douta	=	16'h	4aad;
39756	:douta	=	16'h	4acd;
39757	:douta	=	16'h	52cd;
39758	:douta	=	16'h	530d;
39759	:douta	=	16'h	52ed;
39760	:douta	=	16'h	530d;
39761	:douta	=	16'h	530d;
39762	:douta	=	16'h	52cc;
39763	:douta	=	16'h	634e;
39764	:douta	=	16'h	5b2e;
39765	:douta	=	16'h	5b0d;
39766	:douta	=	16'h	634e;
39767	:douta	=	16'h	5b2d;
39768	:douta	=	16'h	5b0d;
39769	:douta	=	16'h	632d;
39770	:douta	=	16'h	5b2d;
39771	:douta	=	16'h	52ab;
39772	:douta	=	16'h	524a;
39773	:douta	=	16'h	5aab;
39774	:douta	=	16'h	5aec;
39775	:douta	=	16'h	528a;
39776	:douta	=	16'h	528b;
39777	:douta	=	16'h	632d;
39778	:douta	=	16'h	632d;
39779	:douta	=	16'h	5acb;
39780	:douta	=	16'h	62ec;
39781	:douta	=	16'h	62cb;
39782	:douta	=	16'h	5acb;
39783	:douta	=	16'h	630c;
39784	:douta	=	16'h	62ec;
39785	:douta	=	16'h	62cb;
39786	:douta	=	16'h	62cb;
39787	:douta	=	16'h	62cb;
39788	:douta	=	16'h	6b0c;
39789	:douta	=	16'h	6b0c;
39790	:douta	=	16'h	6b2c;
39791	:douta	=	16'h	734d;
39792	:douta	=	16'h	734d;
39793	:douta	=	16'h	7b8e;
39794	:douta	=	16'h	7bcf;
39795	:douta	=	16'h	7baf;
39796	:douta	=	16'h	83ef;
39797	:douta	=	16'h	8c51;
39798	:douta	=	16'h	7b6d;
39799	:douta	=	16'h	83cf;
39800	:douta	=	16'h	736d;
39801	:douta	=	16'h	83cf;
39802	:douta	=	16'h	83d0;
39803	:douta	=	16'h	8431;
39804	:douta	=	16'h	83cf;
39805	:douta	=	16'h	a557;
39806	:douta	=	16'h	a534;
39807	:douta	=	16'h	b533;
39808	:douta	=	16'h	b552;
39809	:douta	=	16'h	cdb3;
39810	:douta	=	16'h	c4ad;
39811	:douta	=	16'h	ccaa;
39812	:douta	=	16'h	d4aa;
39813	:douta	=	16'h	dca7;
39814	:douta	=	16'h	dcc4;
39815	:douta	=	16'h	c468;
39816	:douta	=	16'h	a42c;
39817	:douta	=	16'h	940e;
39818	:douta	=	16'h	7b8f;
39819	:douta	=	16'h	7b6f;
39820	:douta	=	16'h	734f;
39821	:douta	=	16'h	6b2e;
39822	:douta	=	16'h	736d;
39823	:douta	=	16'h	7b4d;
39824	:douta	=	16'h	93ef;
39825	:douta	=	16'h	ee97;
39826	:douta	=	16'h	de76;
39827	:douta	=	16'h	e697;
39828	:douta	=	16'h	d637;
39829	:douta	=	16'h	cdf6;
39830	:douta	=	16'h	7c33;
39831	:douta	=	16'h	bd96;
39832	:douta	=	16'h	c595;
39833	:douta	=	16'h	a517;
39834	:douta	=	16'h	94d5;
39835	:douta	=	16'h	94d5;
39836	:douta	=	16'h	7bf1;
39837	:douta	=	16'h	8412;
39838	:douta	=	16'h	7bd1;
39839	:douta	=	16'h	736f;
39840	:douta	=	16'h	6b70;
39841	:douta	=	16'h	736f;
39842	:douta	=	16'h	6b4f;
39843	:douta	=	16'h	6b2e;
39844	:douta	=	16'h	630e;
39845	:douta	=	16'h	5acd;
39846	:douta	=	16'h	4a4a;
39847	:douta	=	16'h	8bee;
39848	:douta	=	16'h	ac6e;
39849	:douta	=	16'h	cd91;
39850	:douta	=	16'h	de14;
39851	:douta	=	16'h	e656;
39852	:douta	=	16'h	e677;
39853	:douta	=	16'h	de35;
39854	:douta	=	16'h	e656;
39855	:douta	=	16'h	ddf5;
39856	:douta	=	16'h	bd33;
39857	:douta	=	16'h	ad14;
39858	:douta	=	16'h	b555;
39859	:douta	=	16'h	bd95;
39860	:douta	=	16'h	ad55;
39861	:douta	=	16'h	a4f5;
39862	:douta	=	16'h	8c53;
39863	:douta	=	16'h	8c74;
39864	:douta	=	16'h	7bd1;
39865	:douta	=	16'h	73b0;
39866	:douta	=	16'h	7bd0;
39867	:douta	=	16'h	7bd1;
39868	:douta	=	16'h	6b8f;
39869	:douta	=	16'h	7390;
39870	:douta	=	16'h	7390;
39871	:douta	=	16'h	6b4f;
39872	:douta	=	16'h	734f;
39873	:douta	=	16'h	6b2d;
39874	:douta	=	16'h	6b0d;
39875	:douta	=	16'h	5acc;
39876	:douta	=	16'h	5aed;
39877	:douta	=	16'h	632e;
39878	:douta	=	16'h	524a;
39879	:douta	=	16'h	5a8a;
39880	:douta	=	16'h	730c;
39881	:douta	=	16'h	62cb;
39882	:douta	=	16'h	7b6c;
39883	:douta	=	16'h	942e;
39884	:douta	=	16'h	9c4f;
39885	:douta	=	16'h	accf;
39886	:douta	=	16'h	b510;
39887	:douta	=	16'h	d5d3;
39888	:douta	=	16'h	de35;
39889	:douta	=	16'h	de14;
39890	:douta	=	16'h	bd33;
39891	:douta	=	16'h	acf4;
39892	:douta	=	16'h	8c73;
39893	:douta	=	16'h	7c12;
39894	:douta	=	16'h	7c12;
39895	:douta	=	16'h	5b30;
39896	:douta	=	16'h	42ae;
39897	:douta	=	16'h	3a4c;
39898	:douta	=	16'h	31eb;
39899	:douta	=	16'h	31ea;
39900	:douta	=	16'h	426d;
39901	:douta	=	16'h	3a2b;
39902	:douta	=	16'h	1905;
39903	:douta	=	16'h	1906;
39904	:douta	=	16'h	2147;
39905	:douta	=	16'h	1106;
39906	:douta	=	16'h	2105;
39907	:douta	=	16'h	8286;
39908	:douta	=	16'h	6a44;
39909	:douta	=	16'h	7225;
39910	:douta	=	16'h	6a25;
39911	:douta	=	16'h	6a04;
39912	:douta	=	16'h	6a25;
39913	:douta	=	16'h	61e5;
39914	:douta	=	16'h	6205;
39915	:douta	=	16'h	61e4;
39916	:douta	=	16'h	61e5;
39917	:douta	=	16'h	59e5;
39918	:douta	=	16'h	59e5;
39919	:douta	=	16'h	59c5;
39920	:douta	=	16'h	51a5;
39921	:douta	=	16'h	59c5;
39922	:douta	=	16'h	59c5;
39923	:douta	=	16'h	51c5;
39924	:douta	=	16'h	51c5;
39925	:douta	=	16'h	51c6;
39926	:douta	=	16'h	51c5;
39927	:douta	=	16'h	51c5;
39928	:douta	=	16'h	49a6;
39929	:douta	=	16'h	49a6;
39930	:douta	=	16'h	4986;
39931	:douta	=	16'h	49a6;
39932	:douta	=	16'h	4986;
39933	:douta	=	16'h	4185;
39934	:douta	=	16'h	4165;
39935	:douta	=	16'h	41a6;
39936	:douta	=	16'h	de32;
39937	:douta	=	16'h	ddcf;
39938	:douta	=	16'h	d58e;
39939	:douta	=	16'h	ff5b;
39940	:douta	=	16'h	f6f8;
39941	:douta	=	16'h	f719;
39942	:douta	=	16'h	ff3a;
39943	:douta	=	16'h	ff3a;
39944	:douta	=	16'h	f719;
39945	:douta	=	16'h	f719;
39946	:douta	=	16'h	ff7c;
39947	:douta	=	16'h	eeb7;
39948	:douta	=	16'h	de16;
39949	:douta	=	16'h	a4d5;
39950	:douta	=	16'h	8c54;
39951	:douta	=	16'h	94b5;
39952	:douta	=	16'h	8c74;
39953	:douta	=	16'h	94b5;
39954	:douta	=	16'h	8412;
39955	:douta	=	16'h	8c74;
39956	:douta	=	16'h	94b6;
39957	:douta	=	16'h	8cb5;
39958	:douta	=	16'h	9d17;
39959	:douta	=	16'h	1105;
39960	:douta	=	16'h	0842;
39961	:douta	=	16'h	0841;
39962	:douta	=	16'h	0882;
39963	:douta	=	16'h	10c4;
39964	:douta	=	16'h	1905;
39965	:douta	=	16'h	2147;
39966	:douta	=	16'h	1927;
39967	:douta	=	16'h	1905;
39968	:douta	=	16'h	10e5;
39969	:douta	=	16'h	10e5;
39970	:douta	=	16'h	1927;
39971	:douta	=	16'h	1948;
39972	:douta	=	16'h	1947;
39973	:douta	=	16'h	1127;
39974	:douta	=	16'h	1968;
39975	:douta	=	16'h	2168;
39976	:douta	=	16'h	2168;
39977	:douta	=	16'h	2189;
39978	:douta	=	16'h	2189;
39979	:douta	=	16'h	1927;
39980	:douta	=	16'h	2188;
39981	:douta	=	16'h	2168;
39982	:douta	=	16'h	2988;
39983	:douta	=	16'h	2147;
39984	:douta	=	16'h	10e5;
39985	:douta	=	16'h	1926;
39986	:douta	=	16'h	2988;
39987	:douta	=	16'h	31ca;
39988	:douta	=	16'h	31c9;
39989	:douta	=	16'h	31ea;
39990	:douta	=	16'h	9c31;
39991	:douta	=	16'h	73d2;
39992	:douta	=	16'h	4332;
39993	:douta	=	16'h	3a4d;
39994	:douta	=	16'h	2988;
39995	:douta	=	16'h	31ca;
39996	:douta	=	16'h	2988;
39997	:douta	=	16'h	3a2b;
39998	:douta	=	16'h	31ca;
39999	:douta	=	16'h	2988;
40000	:douta	=	16'h	39e9;
40001	:douta	=	16'h	39c9;
40002	:douta	=	16'h	2988;
40003	:douta	=	16'h	31c9;
40004	:douta	=	16'h	2988;
40005	:douta	=	16'h	2147;
40006	:douta	=	16'h	29a9;
40007	:douta	=	16'h	3a2b;
40008	:douta	=	16'h	3a4b;
40009	:douta	=	16'h	428c;
40010	:douta	=	16'h	4aad;
40011	:douta	=	16'h	4aad;
40012	:douta	=	16'h	4aac;
40013	:douta	=	16'h	4aad;
40014	:douta	=	16'h	52cd;
40015	:douta	=	16'h	52ed;
40016	:douta	=	16'h	52ed;
40017	:douta	=	16'h	52ed;
40018	:douta	=	16'h	52cc;
40019	:douta	=	16'h	52ed;
40020	:douta	=	16'h	5b0d;
40021	:douta	=	16'h	52cd;
40022	:douta	=	16'h	5b2d;
40023	:douta	=	16'h	5b2d;
40024	:douta	=	16'h	52cc;
40025	:douta	=	16'h	52ab;
40026	:douta	=	16'h	5b0d;
40027	:douta	=	16'h	62ed;
40028	:douta	=	16'h	528b;
40029	:douta	=	16'h	5aab;
40030	:douta	=	16'h	5aab;
40031	:douta	=	16'h	5acb;
40032	:douta	=	16'h	634d;
40033	:douta	=	16'h	6b6e;
40034	:douta	=	16'h	73af;
40035	:douta	=	16'h	62ec;
40036	:douta	=	16'h	62eb;
40037	:douta	=	16'h	5aaa;
40038	:douta	=	16'h	630c;
40039	:douta	=	16'h	62ec;
40040	:douta	=	16'h	62cb;
40041	:douta	=	16'h	62cb;
40042	:douta	=	16'h	732c;
40043	:douta	=	16'h	6b0c;
40044	:douta	=	16'h	6b0c;
40045	:douta	=	16'h	6b2c;
40046	:douta	=	16'h	738d;
40047	:douta	=	16'h	736e;
40048	:douta	=	16'h	7b8e;
40049	:douta	=	16'h	83cf;
40050	:douta	=	16'h	8c31;
40051	:douta	=	16'h	8410;
40052	:douta	=	16'h	7bcf;
40053	:douta	=	16'h	83ef;
40054	:douta	=	16'h	83f0;
40055	:douta	=	16'h	7bef;
40056	:douta	=	16'h	8c51;
40057	:douta	=	16'h	a4f3;
40058	:douta	=	16'h	ad55;
40059	:douta	=	16'h	c638;
40060	:douta	=	16'h	ce38;
40061	:douta	=	16'h	e6b7;
40062	:douta	=	16'h	cd0c;
40063	:douta	=	16'h	d4ea;
40064	:douta	=	16'h	d4a7;
40065	:douta	=	16'h	d466;
40066	:douta	=	16'h	dc85;
40067	:douta	=	16'h	cc23;
40068	:douta	=	16'h	cc44;
40069	:douta	=	16'h	d446;
40070	:douta	=	16'h	cc46;
40071	:douta	=	16'h	dc84;
40072	:douta	=	16'h	dc84;
40073	:douta	=	16'h	d467;
40074	:douta	=	16'h	bc4b;
40075	:douta	=	16'h	b42a;
40076	:douta	=	16'h	b42c;
40077	:douta	=	16'h	ac2c;
40078	:douta	=	16'h	cdd5;
40079	:douta	=	16'h	d5d4;
40080	:douta	=	16'h	e677;
40081	:douta	=	16'h	d5f6;
40082	:douta	=	16'h	de16;
40083	:douta	=	16'h	d5f6;
40084	:douta	=	16'h	c5d7;
40085	:douta	=	16'h	b597;
40086	:douta	=	16'h	7c33;
40087	:douta	=	16'h	bd96;
40088	:douta	=	16'h	c5b6;
40089	:douta	=	16'h	94d5;
40090	:douta	=	16'h	9495;
40091	:douta	=	16'h	8c53;
40092	:douta	=	16'h	7bd1;
40093	:douta	=	16'h	7bb0;
40094	:douta	=	16'h	7bb0;
40095	:douta	=	16'h	736f;
40096	:douta	=	16'h	7390;
40097	:douta	=	16'h	62ed;
40098	:douta	=	16'h	62cd;
40099	:douta	=	16'h	52ad;
40100	:douta	=	16'h	52ad;
40101	:douta	=	16'h	4a2a;
40102	:douta	=	16'h	b4d1;
40103	:douta	=	16'h	e634;
40104	:douta	=	16'h	d5f4;
40105	:douta	=	16'h	e656;
40106	:douta	=	16'h	e656;
40107	:douta	=	16'h	e656;
40108	:douta	=	16'h	e656;
40109	:douta	=	16'h	d5d5;
40110	:douta	=	16'h	d5f6;
40111	:douta	=	16'h	d5d5;
40112	:douta	=	16'h	cdb4;
40113	:douta	=	16'h	b514;
40114	:douta	=	16'h	ad14;
40115	:douta	=	16'h	b556;
40116	:douta	=	16'h	b556;
40117	:douta	=	16'h	ad16;
40118	:douta	=	16'h	8452;
40119	:douta	=	16'h	8433;
40120	:douta	=	16'h	8412;
40121	:douta	=	16'h	7bd0;
40122	:douta	=	16'h	7bb0;
40123	:douta	=	16'h	7391;
40124	:douta	=	16'h	73b0;
40125	:douta	=	16'h	6b6f;
40126	:douta	=	16'h	73b0;
40127	:douta	=	16'h	6b4f;
40128	:douta	=	16'h	5acd;
40129	:douta	=	16'h	6b2e;
40130	:douta	=	16'h	736f;
40131	:douta	=	16'h	6b2e;
40132	:douta	=	16'h	6b2d;
40133	:douta	=	16'h	41e7;
40134	:douta	=	16'h	3965;
40135	:douta	=	16'h	5a47;
40136	:douta	=	16'h	9c4e;
40137	:douta	=	16'h	acf0;
40138	:douta	=	16'h	bd51;
40139	:douta	=	16'h	cdb2;
40140	:douta	=	16'h	d5b3;
40141	:douta	=	16'h	cdd2;
40142	:douta	=	16'h	d5f3;
40143	:douta	=	16'h	de34;
40144	:douta	=	16'h	de15;
40145	:douta	=	16'h	d5d3;
40146	:douta	=	16'h	b534;
40147	:douta	=	16'h	acf4;
40148	:douta	=	16'h	8c73;
40149	:douta	=	16'h	7c33;
40150	:douta	=	16'h	7c33;
40151	:douta	=	16'h	5b50;
40152	:douta	=	16'h	5310;
40153	:douta	=	16'h	42ce;
40154	:douta	=	16'h	3a4c;
40155	:douta	=	16'h	320b;
40156	:douta	=	16'h	2168;
40157	:douta	=	16'h	4ace;
40158	:douta	=	16'h	10c5;
40159	:douta	=	16'h	2127;
40160	:douta	=	16'h	1926;
40161	:douta	=	16'h	2146;
40162	:douta	=	16'h	00a5;
40163	:douta	=	16'h	82a5;
40164	:douta	=	16'h	7244;
40165	:douta	=	16'h	7245;
40166	:douta	=	16'h	7225;
40167	:douta	=	16'h	6a24;
40168	:douta	=	16'h	6a04;
40169	:douta	=	16'h	6205;
40170	:douta	=	16'h	6205;
40171	:douta	=	16'h	61e4;
40172	:douta	=	16'h	6205;
40173	:douta	=	16'h	61e5;
40174	:douta	=	16'h	59e5;
40175	:douta	=	16'h	59c5;
40176	:douta	=	16'h	59c5;
40177	:douta	=	16'h	59c5;
40178	:douta	=	16'h	59c5;
40179	:douta	=	16'h	51c5;
40180	:douta	=	16'h	51c6;
40181	:douta	=	16'h	51a5;
40182	:douta	=	16'h	51c5;
40183	:douta	=	16'h	51c6;
40184	:douta	=	16'h	49a6;
40185	:douta	=	16'h	49a6;
40186	:douta	=	16'h	49a6;
40187	:douta	=	16'h	4986;
40188	:douta	=	16'h	49a5;
40189	:douta	=	16'h	4185;
40190	:douta	=	16'h	4165;
40191	:douta	=	16'h	4165;
40192	:douta	=	16'h	ee95;
40193	:douta	=	16'h	e674;
40194	:douta	=	16'h	e675;
40195	:douta	=	16'h	f71a;
40196	:douta	=	16'h	f6f9;
40197	:douta	=	16'h	f71a;
40198	:douta	=	16'h	ff39;
40199	:douta	=	16'h	f739;
40200	:douta	=	16'h	ff19;
40201	:douta	=	16'h	ff3a;
40202	:douta	=	16'h	ff9c;
40203	:douta	=	16'h	de57;
40204	:douta	=	16'h	bd34;
40205	:douta	=	16'h	a4f5;
40206	:douta	=	16'h	9494;
40207	:douta	=	16'h	94b5;
40208	:douta	=	16'h	94d6;
40209	:douta	=	16'h	9494;
40210	:douta	=	16'h	9432;
40211	:douta	=	16'h	94d5;
40212	:douta	=	16'h	94d6;
40213	:douta	=	16'h	94d6;
40214	:douta	=	16'h	8cb5;
40215	:douta	=	16'h	63b3;
40216	:douta	=	16'h	7456;
40217	:douta	=	16'h	7436;
40218	:douta	=	16'h	63d3;
40219	:douta	=	16'h	42ae;
40220	:douta	=	16'h	0000;
40221	:douta	=	16'h	10c4;
40222	:douta	=	16'h	10e5;
40223	:douta	=	16'h	1926;
40224	:douta	=	16'h	1905;
40225	:douta	=	16'h	1927;
40226	:douta	=	16'h	1967;
40227	:douta	=	16'h	1947;
40228	:douta	=	16'h	1968;
40229	:douta	=	16'h	1948;
40230	:douta	=	16'h	1948;
40231	:douta	=	16'h	1948;
40232	:douta	=	16'h	1148;
40233	:douta	=	16'h	2168;
40234	:douta	=	16'h	1968;
40235	:douta	=	16'h	1926;
40236	:douta	=	16'h	18e4;
40237	:douta	=	16'h	10c5;
40238	:douta	=	16'h	1967;
40239	:douta	=	16'h	2188;
40240	:douta	=	16'h	29a9;
40241	:douta	=	16'h	29ca;
40242	:douta	=	16'h	29a9;
40243	:douta	=	16'h	1906;
40244	:douta	=	16'h	1926;
40245	:douta	=	16'h	2967;
40246	:douta	=	16'h	2988;
40247	:douta	=	16'h	2988;
40248	:douta	=	16'h	2967;
40249	:douta	=	16'h	2147;
40250	:douta	=	16'h	2988;
40251	:douta	=	16'h	3189;
40252	:douta	=	16'h	2988;
40253	:douta	=	16'h	2988;
40254	:douta	=	16'h	2988;
40255	:douta	=	16'h	3188;
40256	:douta	=	16'h	2968;
40257	:douta	=	16'h	2988;
40258	:douta	=	16'h	31a9;
40259	:douta	=	16'h	31e9;
40260	:douta	=	16'h	3a0a;
40261	:douta	=	16'h	31e9;
40262	:douta	=	16'h	3a2b;
40263	:douta	=	16'h	322a;
40264	:douta	=	16'h	322a;
40265	:douta	=	16'h	3a4b;
40266	:douta	=	16'h	424b;
40267	:douta	=	16'h	426b;
40268	:douta	=	16'h	426c;
40269	:douta	=	16'h	428c;
40270	:douta	=	16'h	4aac;
40271	:douta	=	16'h	4a8c;
40272	:douta	=	16'h	4aac;
40273	:douta	=	16'h	52cd;
40274	:douta	=	16'h	52ad;
40275	:douta	=	16'h	52ed;
40276	:douta	=	16'h	5b0d;
40277	:douta	=	16'h	5b2e;
40278	:douta	=	16'h	52cc;
40279	:douta	=	16'h	5acc;
40280	:douta	=	16'h	5aec;
40281	:douta	=	16'h	632d;
40282	:douta	=	16'h	5aec;
40283	:douta	=	16'h	5aec;
40284	:douta	=	16'h	630c;
40285	:douta	=	16'h	5aab;
40286	:douta	=	16'h	52aa;
40287	:douta	=	16'h	630c;
40288	:douta	=	16'h	5249;
40289	:douta	=	16'h	4a48;
40290	:douta	=	16'h	5249;
40291	:douta	=	16'h	5a8a;
40292	:douta	=	16'h	5aab;
40293	:douta	=	16'h	734d;
40294	:douta	=	16'h	630c;
40295	:douta	=	16'h	62ec;
40296	:douta	=	16'h	62eb;
40297	:douta	=	16'h	736d;
40298	:douta	=	16'h	83ef;
40299	:douta	=	16'h	83ef;
40300	:douta	=	16'h	83f0;
40301	:douta	=	16'h	8c31;
40302	:douta	=	16'h	7bd0;
40303	:douta	=	16'h	8411;
40304	:douta	=	16'h	9cf4;
40305	:douta	=	16'h	a555;
40306	:douta	=	16'h	adb6;
40307	:douta	=	16'h	ce38;
40308	:douta	=	16'h	d5b1;
40309	:douta	=	16'h	cd6f;
40310	:douta	=	16'h	e5f2;
40311	:douta	=	16'h	e5b0;
40312	:douta	=	16'h	dd2c;
40313	:douta	=	16'h	d467;
40314	:douta	=	16'h	cc02;
40315	:douta	=	16'h	c3e1;
40316	:douta	=	16'h	cbe2;
40317	:douta	=	16'h	cc24;
40318	:douta	=	16'h	cc45;
40319	:douta	=	16'h	cc25;
40320	:douta	=	16'h	cc45;
40321	:douta	=	16'h	cc65;
40322	:douta	=	16'h	cc46;
40323	:douta	=	16'h	cc66;
40324	:douta	=	16'h	cc65;
40325	:douta	=	16'h	d467;
40326	:douta	=	16'h	d466;
40327	:douta	=	16'h	d466;
40328	:douta	=	16'h	d466;
40329	:douta	=	16'h	d466;
40330	:douta	=	16'h	cc66;
40331	:douta	=	16'h	d466;
40332	:douta	=	16'h	d466;
40333	:douta	=	16'h	d465;
40334	:douta	=	16'h	cc23;
40335	:douta	=	16'h	b4d2;
40336	:douta	=	16'h	b514;
40337	:douta	=	16'h	bd97;
40338	:douta	=	16'h	ad36;
40339	:douta	=	16'h	ad16;
40340	:douta	=	16'h	ad77;
40341	:douta	=	16'h	ad57;
40342	:douta	=	16'h	8453;
40343	:douta	=	16'h	b596;
40344	:douta	=	16'h	c596;
40345	:douta	=	16'h	8c53;
40346	:douta	=	16'h	8412;
40347	:douta	=	16'h	7bf2;
40348	:douta	=	16'h	8412;
40349	:douta	=	16'h	8411;
40350	:douta	=	16'h	732e;
40351	:douta	=	16'h	6b2e;
40352	:douta	=	16'h	62cd;
40353	:douta	=	16'h	5acc;
40354	:douta	=	16'h	4a4b;
40355	:douta	=	16'h	acd2;
40356	:douta	=	16'h	a48f;
40357	:douta	=	16'h	a4b0;
40358	:douta	=	16'h	e697;
40359	:douta	=	16'h	cdf4;
40360	:douta	=	16'h	d5b4;
40361	:douta	=	16'h	cd94;
40362	:douta	=	16'h	de55;
40363	:douta	=	16'h	d5f4;
40364	:douta	=	16'h	cdb5;
40365	:douta	=	16'h	c576;
40366	:douta	=	16'h	b555;
40367	:douta	=	16'h	b556;
40368	:douta	=	16'h	b535;
40369	:douta	=	16'h	b535;
40370	:douta	=	16'h	9cb4;
40371	:douta	=	16'h	9cf5;
40372	:douta	=	16'h	a4d5;
40373	:douta	=	16'h	9cb5;
40374	:douta	=	16'h	73d1;
40375	:douta	=	16'h	6b4f;
40376	:douta	=	16'h	6b2f;
40377	:douta	=	16'h	7bd1;
40378	:douta	=	16'h	6b70;
40379	:douta	=	16'h	83f1;
40380	:douta	=	16'h	6b8f;
40381	:douta	=	16'h	632f;
40382	:douta	=	16'h	5b0d;
40383	:douta	=	16'h	630e;
40384	:douta	=	16'h	630e;
40385	:douta	=	16'h	4a29;
40386	:douta	=	16'h	41c7;
40387	:douta	=	16'h	3123;
40388	:douta	=	16'h	28c3;
40389	:douta	=	16'h	5248;
40390	:douta	=	16'h	5a48;
40391	:douta	=	16'h	5a89;
40392	:douta	=	16'h	730b;
40393	:douta	=	16'h	732b;
40394	:douta	=	16'h	a48e;
40395	:douta	=	16'h	cdd3;
40396	:douta	=	16'h	d614;
40397	:douta	=	16'h	e656;
40398	:douta	=	16'h	e656;
40399	:douta	=	16'h	de35;
40400	:douta	=	16'h	d5d4;
40401	:douta	=	16'h	cd73;
40402	:douta	=	16'h	acf4;
40403	:douta	=	16'h	a514;
40404	:douta	=	16'h	94b6;
40405	:douta	=	16'h	8495;
40406	:douta	=	16'h	8475;
40407	:douta	=	16'h	5b50;
40408	:douta	=	16'h	4ace;
40409	:douta	=	16'h	4ace;
40410	:douta	=	16'h	3a6d;
40411	:douta	=	16'h	3a6c;
40412	:douta	=	16'h	31ec;
40413	:douta	=	16'h	2168;
40414	:douta	=	16'h	31c9;
40415	:douta	=	16'h	2988;
40416	:douta	=	16'h	1905;
40417	:douta	=	16'h	10c5;
40418	:douta	=	16'h	1905;
40419	:douta	=	16'h	3965;
40420	:douta	=	16'h	7245;
40421	:douta	=	16'h	7245;
40422	:douta	=	16'h	6a24;
40423	:douta	=	16'h	6a25;
40424	:douta	=	16'h	6a25;
40425	:douta	=	16'h	6205;
40426	:douta	=	16'h	6205;
40427	:douta	=	16'h	61e4;
40428	:douta	=	16'h	61e5;
40429	:douta	=	16'h	59e5;
40430	:douta	=	16'h	59e5;
40431	:douta	=	16'h	59c5;
40432	:douta	=	16'h	59c5;
40433	:douta	=	16'h	51a5;
40434	:douta	=	16'h	59e6;
40435	:douta	=	16'h	59e6;
40436	:douta	=	16'h	51c6;
40437	:douta	=	16'h	51c5;
40438	:douta	=	16'h	51c5;
40439	:douta	=	16'h	51c5;
40440	:douta	=	16'h	49a6;
40441	:douta	=	16'h	49a6;
40442	:douta	=	16'h	49a5;
40443	:douta	=	16'h	49a6;
40444	:douta	=	16'h	4985;
40445	:douta	=	16'h	4185;
40446	:douta	=	16'h	4165;
40447	:douta	=	16'h	4165;
40448	:douta	=	16'h	eeb6;
40449	:douta	=	16'h	e694;
40450	:douta	=	16'h	f6d8;
40451	:douta	=	16'h	f719;
40452	:douta	=	16'h	fef9;
40453	:douta	=	16'h	ff3a;
40454	:douta	=	16'h	ff19;
40455	:douta	=	16'h	f719;
40456	:douta	=	16'h	f719;
40457	:douta	=	16'h	ff5b;
40458	:douta	=	16'h	ff9b;
40459	:douta	=	16'h	d5d6;
40460	:douta	=	16'h	b535;
40461	:douta	=	16'h	9c95;
40462	:douta	=	16'h	9cf6;
40463	:douta	=	16'h	9cd5;
40464	:douta	=	16'h	94d5;
40465	:douta	=	16'h	8c73;
40466	:douta	=	16'h	9c94;
40467	:douta	=	16'h	94d5;
40468	:douta	=	16'h	94d6;
40469	:douta	=	16'h	9cf6;
40470	:douta	=	16'h	8c75;
40471	:douta	=	16'h	5b72;
40472	:douta	=	16'h	7415;
40473	:douta	=	16'h	7456;
40474	:douta	=	16'h	84d8;
40475	:douta	=	16'h	8d3a;
40476	:douta	=	16'h	21a8;
40477	:douta	=	16'h	0882;
40478	:douta	=	16'h	10a3;
40479	:douta	=	16'h	10e5;
40480	:douta	=	16'h	10e4;
40481	:douta	=	16'h	1906;
40482	:douta	=	16'h	1127;
40483	:douta	=	16'h	1927;
40484	:douta	=	16'h	1947;
40485	:douta	=	16'h	1948;
40486	:douta	=	16'h	2169;
40487	:douta	=	16'h	1968;
40488	:douta	=	16'h	2188;
40489	:douta	=	16'h	1927;
40490	:douta	=	16'h	1947;
40491	:douta	=	16'h	1946;
40492	:douta	=	16'h	1947;
40493	:douta	=	16'h	10e4;
40494	:douta	=	16'h	2168;
40495	:douta	=	16'h	29a9;
40496	:douta	=	16'h	2189;
40497	:douta	=	16'h	21a8;
40498	:douta	=	16'h	29a9;
40499	:douta	=	16'h	29a9;
40500	:douta	=	16'h	2187;
40501	:douta	=	16'h	31a9;
40502	:douta	=	16'h	2126;
40503	:douta	=	16'h	1906;
40504	:douta	=	16'h	1906;
40505	:douta	=	16'h	2988;
40506	:douta	=	16'h	2168;
40507	:douta	=	16'h	2167;
40508	:douta	=	16'h	2167;
40509	:douta	=	16'h	2147;
40510	:douta	=	16'h	2126;
40511	:douta	=	16'h	2106;
40512	:douta	=	16'h	1082;
40513	:douta	=	16'h	2127;
40514	:douta	=	16'h	31c9;
40515	:douta	=	16'h	31c9;
40516	:douta	=	16'h	2106;
40517	:douta	=	16'h	3a0a;
40518	:douta	=	16'h	31ea;
40519	:douta	=	16'h	31e9;
40520	:douta	=	16'h	3a0a;
40521	:douta	=	16'h	3a0a;
40522	:douta	=	16'h	424b;
40523	:douta	=	16'h	428c;
40524	:douta	=	16'h	4aad;
40525	:douta	=	16'h	4acd;
40526	:douta	=	16'h	424a;
40527	:douta	=	16'h	4aac;
40528	:douta	=	16'h	4a8c;
40529	:douta	=	16'h	52cc;
40530	:douta	=	16'h	4aac;
40531	:douta	=	16'h	52ac;
40532	:douta	=	16'h	4a8b;
40533	:douta	=	16'h	4a8b;
40534	:douta	=	16'h	4249;
40535	:douta	=	16'h	4249;
40536	:douta	=	16'h	4a4a;
40537	:douta	=	16'h	630d;
40538	:douta	=	16'h	5b0d;
40539	:douta	=	16'h	52cb;
40540	:douta	=	16'h	52cc;
40541	:douta	=	16'h	5aab;
40542	:douta	=	16'h	5269;
40543	:douta	=	16'h	5acb;
40544	:douta	=	16'h	5aaa;
40545	:douta	=	16'h	62eb;
40546	:douta	=	16'h	738f;
40547	:douta	=	16'h	6b8e;
40548	:douta	=	16'h	6b0c;
40549	:douta	=	16'h	6b2c;
40550	:douta	=	16'h	736e;
40551	:douta	=	16'h	62ec;
40552	:douta	=	16'h	6b2d;
40553	:douta	=	16'h	6b6e;
40554	:douta	=	16'h	7bf1;
40555	:douta	=	16'h	73b0;
40556	:douta	=	16'h	83cf;
40557	:douta	=	16'h	8c50;
40558	:douta	=	16'h	b553;
40559	:douta	=	16'h	d615;
40560	:douta	=	16'h	e6b8;
40561	:douta	=	16'h	ddb0;
40562	:douta	=	16'h	e5d0;
40563	:douta	=	16'h	e56d;
40564	:douta	=	16'h	cc24;
40565	:douta	=	16'h	d443;
40566	:douta	=	16'h	c3c2;
40567	:douta	=	16'h	c3c2;
40568	:douta	=	16'h	c3c2;
40569	:douta	=	16'h	c403;
40570	:douta	=	16'h	cc25;
40571	:douta	=	16'h	cc25;
40572	:douta	=	16'h	cc25;
40573	:douta	=	16'h	cc25;
40574	:douta	=	16'h	cc25;
40575	:douta	=	16'h	cc25;
40576	:douta	=	16'h	cc66;
40577	:douta	=	16'h	cc45;
40578	:douta	=	16'h	cc66;
40579	:douta	=	16'h	d466;
40580	:douta	=	16'h	cc45;
40581	:douta	=	16'h	cc66;
40582	:douta	=	16'h	cc66;
40583	:douta	=	16'h	cc66;
40584	:douta	=	16'h	cc66;
40585	:douta	=	16'h	d466;
40586	:douta	=	16'h	d466;
40587	:douta	=	16'h	cc66;
40588	:douta	=	16'h	d466;
40589	:douta	=	16'h	d467;
40590	:douta	=	16'h	d466;
40591	:douta	=	16'h	c447;
40592	:douta	=	16'h	b4b2;
40593	:douta	=	16'h	b535;
40594	:douta	=	16'h	a4f4;
40595	:douta	=	16'h	a4d4;
40596	:douta	=	16'h	a4d5;
40597	:douta	=	16'h	a4f6;
40598	:douta	=	16'h	8c53;
40599	:douta	=	16'h	b576;
40600	:douta	=	16'h	c5d7;
40601	:douta	=	16'h	8c73;
40602	:douta	=	16'h	8453;
40603	:douta	=	16'h	7bd1;
40604	:douta	=	16'h	7bb1;
40605	:douta	=	16'h	7bf1;
40606	:douta	=	16'h	7bb0;
40607	:douta	=	16'h	736f;
40608	:douta	=	16'h	52ac;
40609	:douta	=	16'h	41e9;
40610	:douta	=	16'h	9410;
40611	:douta	=	16'h	d5d4;
40612	:douta	=	16'h	8bee;
40613	:douta	=	16'h	ee97;
40614	:douta	=	16'h	de15;
40615	:douta	=	16'h	ddf5;
40616	:douta	=	16'h	de15;
40617	:douta	=	16'h	c553;
40618	:douta	=	16'h	d5f5;
40619	:douta	=	16'h	cdb4;
40620	:douta	=	16'h	bd56;
40621	:douta	=	16'h	b536;
40622	:douta	=	16'h	a4d6;
40623	:douta	=	16'h	9c95;
40624	:douta	=	16'h	9cd5;
40625	:douta	=	16'h	9cd5;
40626	:douta	=	16'h	a4d5;
40627	:douta	=	16'h	acf5;
40628	:douta	=	16'h	9494;
40629	:douta	=	16'h	9cb5;
40630	:douta	=	16'h	8432;
40631	:douta	=	16'h	6b70;
40632	:douta	=	16'h	62ed;
40633	:douta	=	16'h	73b0;
40634	:douta	=	16'h	6b6f;
40635	:douta	=	16'h	6b4f;
40636	:douta	=	16'h	7bf1;
40637	:douta	=	16'h	7390;
40638	:douta	=	16'h	5b0e;
40639	:douta	=	16'h	630d;
40640	:douta	=	16'h	41e8;
40641	:douta	=	16'h	3186;
40642	:douta	=	16'h	3985;
40643	:douta	=	16'h	62c9;
40644	:douta	=	16'h	732a;
40645	:douta	=	16'h	8bcd;
40646	:douta	=	16'h	942d;
40647	:douta	=	16'h	a4af;
40648	:douta	=	16'h	a4ef;
40649	:douta	=	16'h	a4af;
40650	:douta	=	16'h	9c2e;
40651	:douta	=	16'h	bd4f;
40652	:douta	=	16'h	cdb2;
40653	:douta	=	16'h	de35;
40654	:douta	=	16'h	de15;
40655	:douta	=	16'h	d614;
40656	:douta	=	16'h	c554;
40657	:douta	=	16'h	ad14;
40658	:douta	=	16'h	ad15;
40659	:douta	=	16'h	a4f5;
40660	:douta	=	16'h	94d5;
40661	:douta	=	16'h	8454;
40662	:douta	=	16'h	7c34;
40663	:douta	=	16'h	6bf2;
40664	:douta	=	16'h	5b50;
40665	:douta	=	16'h	4aef;
40666	:douta	=	16'h	4aae;
40667	:douta	=	16'h	428e;
40668	:douta	=	16'h	3a4d;
40669	:douta	=	16'h	29aa;
40670	:douta	=	16'h	532f;
40671	:douta	=	16'h	2147;
40672	:douta	=	16'h	1905;
40673	:douta	=	16'h	10e5;
40674	:douta	=	16'h	18e5;
40675	:douta	=	16'h	00a5;
40676	:douta	=	16'h	8286;
40677	:douta	=	16'h	7a45;
40678	:douta	=	16'h	7225;
40679	:douta	=	16'h	7225;
40680	:douta	=	16'h	6a04;
40681	:douta	=	16'h	6a05;
40682	:douta	=	16'h	6205;
40683	:douta	=	16'h	61e5;
40684	:douta	=	16'h	61e5;
40685	:douta	=	16'h	61e5;
40686	:douta	=	16'h	59e5;
40687	:douta	=	16'h	59c5;
40688	:douta	=	16'h	59c5;
40689	:douta	=	16'h	59c5;
40690	:douta	=	16'h	59e6;
40691	:douta	=	16'h	51e5;
40692	:douta	=	16'h	51c6;
40693	:douta	=	16'h	51c6;
40694	:douta	=	16'h	51c6;
40695	:douta	=	16'h	49c6;
40696	:douta	=	16'h	49a6;
40697	:douta	=	16'h	49a6;
40698	:douta	=	16'h	49a6;
40699	:douta	=	16'h	4985;
40700	:douta	=	16'h	4186;
40701	:douta	=	16'h	4165;
40702	:douta	=	16'h	4185;
40703	:douta	=	16'h	4165;
40704	:douta	=	16'h	f6d7;
40705	:douta	=	16'h	f6f7;
40706	:douta	=	16'h	ff1a;
40707	:douta	=	16'h	f6f9;
40708	:douta	=	16'h	f73a;
40709	:douta	=	16'h	ff3a;
40710	:douta	=	16'h	ff19;
40711	:douta	=	16'h	f6f9;
40712	:douta	=	16'h	ff3a;
40713	:douta	=	16'h	ff9c;
40714	:douta	=	16'h	f6d8;
40715	:douta	=	16'h	c5b6;
40716	:douta	=	16'h	ad16;
40717	:douta	=	16'h	8c53;
40718	:douta	=	16'h	9cf6;
40719	:douta	=	16'h	94b5;
40720	:douta	=	16'h	9cb5;
40721	:douta	=	16'h	9473;
40722	:douta	=	16'h	9c94;
40723	:douta	=	16'h	a517;
40724	:douta	=	16'h	9cf6;
40725	:douta	=	16'h	94b6;
40726	:douta	=	16'h	6c14;
40727	:douta	=	16'h	7435;
40728	:douta	=	16'h	7456;
40729	:douta	=	16'h	6c34;
40730	:douta	=	16'h	7c77;
40731	:douta	=	16'h	8497;
40732	:douta	=	16'h	84b8;
40733	:douta	=	16'h	2a2a;
40734	:douta	=	16'h	0001;
40735	:douta	=	16'h	1105;
40736	:douta	=	16'h	10e5;
40737	:douta	=	16'h	1926;
40738	:douta	=	16'h	1947;
40739	:douta	=	16'h	1947;
40740	:douta	=	16'h	1127;
40741	:douta	=	16'h	1127;
40742	:douta	=	16'h	1967;
40743	:douta	=	16'h	1927;
40744	:douta	=	16'h	1926;
40745	:douta	=	16'h	1947;
40746	:douta	=	16'h	1948;
40747	:douta	=	16'h	1926;
40748	:douta	=	16'h	2167;
40749	:douta	=	16'h	2189;
40750	:douta	=	16'h	18e5;
40751	:douta	=	16'h	1082;
40752	:douta	=	16'h	2188;
40753	:douta	=	16'h	1968;
40754	:douta	=	16'h	2168;
40755	:douta	=	16'h	2168;
40756	:douta	=	16'h	2146;
40757	:douta	=	16'h	1946;
40758	:douta	=	16'h	2126;
40759	:douta	=	16'h	18e4;
40760	:douta	=	16'h	29c9;
40761	:douta	=	16'h	322b;
40762	:douta	=	16'h	3a2b;
40763	:douta	=	16'h	18a1;
40764	:douta	=	16'h	3144;
40765	:douta	=	16'h	0000;
40766	:douta	=	16'h	0800;
40767	:douta	=	16'h	0821;
40768	:douta	=	16'h	0820;
40769	:douta	=	16'h	18e4;
40770	:douta	=	16'h	2126;
40771	:douta	=	16'h	1905;
40772	:douta	=	16'h	29c8;
40773	:douta	=	16'h	31ea;
40774	:douta	=	16'h	31e9;
40775	:douta	=	16'h	3a0a;
40776	:douta	=	16'h	3a2b;
40777	:douta	=	16'h	3a2a;
40778	:douta	=	16'h	31e9;
40779	:douta	=	16'h	31e9;
40780	:douta	=	16'h	31c9;
40781	:douta	=	16'h	31a8;
40782	:douta	=	16'h	39e9;
40783	:douta	=	16'h	39c8;
40784	:douta	=	16'h	4229;
40785	:douta	=	16'h	4a6b;
40786	:douta	=	16'h	4229;
40787	:douta	=	16'h	3a09;
40788	:douta	=	16'h	4a8b;
40789	:douta	=	16'h	4a8b;
40790	:douta	=	16'h	4a4a;
40791	:douta	=	16'h	4a4a;
40792	:douta	=	16'h	526b;
40793	:douta	=	16'h	4a6a;
40794	:douta	=	16'h	5acc;
40795	:douta	=	16'h	638e;
40796	:douta	=	16'h	6baf;
40797	:douta	=	16'h	7390;
40798	:douta	=	16'h	73f1;
40799	:douta	=	16'h	8473;
40800	:douta	=	16'h	73f1;
40801	:douta	=	16'h	6b8f;
40802	:douta	=	16'h	5aed;
40803	:douta	=	16'h	6b8f;
40804	:douta	=	16'h	7b6d;
40805	:douta	=	16'h	93cd;
40806	:douta	=	16'h	ac4e;
40807	:douta	=	16'h	cd70;
40808	:douta	=	16'h	c50e;
40809	:douta	=	16'h	bbc4;
40810	:douta	=	16'h	cc24;
40811	:douta	=	16'h	cbe3;
40812	:douta	=	16'h	c403;
40813	:douta	=	16'h	c3c3;
40814	:douta	=	16'h	bba3;
40815	:douta	=	16'h	c3e2;
40816	:douta	=	16'h	c3e2;
40817	:douta	=	16'h	cc25;
40818	:douta	=	16'h	cc25;
40819	:douta	=	16'h	cc25;
40820	:douta	=	16'h	cc25;
40821	:douta	=	16'h	cc25;
40822	:douta	=	16'h	cc25;
40823	:douta	=	16'h	cc45;
40824	:douta	=	16'h	cc45;
40825	:douta	=	16'h	cc45;
40826	:douta	=	16'h	cc45;
40827	:douta	=	16'h	cc45;
40828	:douta	=	16'h	cc45;
40829	:douta	=	16'h	cc45;
40830	:douta	=	16'h	cc45;
40831	:douta	=	16'h	cc46;
40832	:douta	=	16'h	cc45;
40833	:douta	=	16'h	cc66;
40834	:douta	=	16'h	cc45;
40835	:douta	=	16'h	cc46;
40836	:douta	=	16'h	cc45;
40837	:douta	=	16'h	cc45;
40838	:douta	=	16'h	d465;
40839	:douta	=	16'h	d466;
40840	:douta	=	16'h	cc66;
40841	:douta	=	16'h	d466;
40842	:douta	=	16'h	d466;
40843	:douta	=	16'h	d466;
40844	:douta	=	16'h	cc66;
40845	:douta	=	16'h	d465;
40846	:douta	=	16'h	cc66;
40847	:douta	=	16'h	d486;
40848	:douta	=	16'h	d444;
40849	:douta	=	16'h	bcaf;
40850	:douta	=	16'h	9c53;
40851	:douta	=	16'h	9c51;
40852	:douta	=	16'h	9c72;
40853	:douta	=	16'h	9451;
40854	:douta	=	16'h	9452;
40855	:douta	=	16'h	a4f5;
40856	:douta	=	16'h	a516;
40857	:douta	=	16'h	8c11;
40858	:douta	=	16'h	8412;
40859	:douta	=	16'h	73d0;
40860	:douta	=	16'h	736f;
40861	:douta	=	16'h	6b4f;
40862	:douta	=	16'h	4a6b;
40863	:douta	=	16'h	732e;
40864	:douta	=	16'h	b4b0;
40865	:douta	=	16'h	e677;
40866	:douta	=	16'h	de36;
40867	:douta	=	16'h	bd52;
40868	:douta	=	16'h	de96;
40869	:douta	=	16'h	e6b7;
40870	:douta	=	16'h	d5b4;
40871	:douta	=	16'h	de15;
40872	:douta	=	16'h	de15;
40873	:douta	=	16'h	d5d5;
40874	:douta	=	16'h	bd34;
40875	:douta	=	16'h	b535;
40876	:douta	=	16'h	9c94;
40877	:douta	=	16'h	9494;
40878	:douta	=	16'h	9494;
40879	:douta	=	16'h	8412;
40880	:douta	=	16'h	83f1;
40881	:douta	=	16'h	8c33;
40882	:douta	=	16'h	8453;
40883	:douta	=	16'h	9494;
40884	:douta	=	16'h	a4f6;
40885	:douta	=	16'h	8c74;
40886	:douta	=	16'h	73d1;
40887	:douta	=	16'h	630e;
40888	:douta	=	16'h	5aee;
40889	:douta	=	16'h	632e;
40890	:douta	=	16'h	632f;
40891	:douta	=	16'h	632f;
40892	:douta	=	16'h	524a;
40893	:douta	=	16'h	41e8;
40894	:douta	=	16'h	3985;
40895	:douta	=	16'h	5228;
40896	:douta	=	16'h	93ed;
40897	:douta	=	16'h	cd52;
40898	:douta	=	16'h	c551;
40899	:douta	=	16'h	c550;
40900	:douta	=	16'h	d5b1;
40901	:douta	=	16'h	de14;
40902	:douta	=	16'h	de35;
40903	:douta	=	16'h	e676;
40904	:douta	=	16'h	e656;
40905	:douta	=	16'h	e676;
40906	:douta	=	16'h	e696;
40907	:douta	=	16'h	e656;
40908	:douta	=	16'h	de35;
40909	:douta	=	16'h	de35;
40910	:douta	=	16'h	e655;
40911	:douta	=	16'h	cdb5;
40912	:douta	=	16'h	ad16;
40913	:douta	=	16'h	9cf5;
40914	:douta	=	16'h	9cf5;
40915	:douta	=	16'h	94d5;
40916	:douta	=	16'h	94d6;
40917	:douta	=	16'h	8475;
40918	:douta	=	16'h	7c34;
40919	:douta	=	16'h	6bf3;
40920	:douta	=	16'h	7414;
40921	:douta	=	16'h	6bb2;
40922	:douta	=	16'h	5330;
40923	:douta	=	16'h	4b10;
40924	:douta	=	16'h	5331;
40925	:douta	=	16'h	530f;
40926	:douta	=	16'h	52ef;
40927	:douta	=	16'h	1106;
40928	:douta	=	16'h	2168;
40929	:douta	=	16'h	2168;
40930	:douta	=	16'h	2127;
40931	:douta	=	16'h	10c6;
40932	:douta	=	16'h	8a85;
40933	:douta	=	16'h	7226;
40934	:douta	=	16'h	6a24;
40935	:douta	=	16'h	6a24;
40936	:douta	=	16'h	6a05;
40937	:douta	=	16'h	6a05;
40938	:douta	=	16'h	61e5;
40939	:douta	=	16'h	6205;
40940	:douta	=	16'h	61e5;
40941	:douta	=	16'h	59e5;
40942	:douta	=	16'h	59c5;
40943	:douta	=	16'h	59c5;
40944	:douta	=	16'h	59c5;
40945	:douta	=	16'h	59c5;
40946	:douta	=	16'h	59c6;
40947	:douta	=	16'h	51c6;
40948	:douta	=	16'h	51c6;
40949	:douta	=	16'h	51c5;
40950	:douta	=	16'h	49c6;
40951	:douta	=	16'h	49c6;
40952	:douta	=	16'h	49a5;
40953	:douta	=	16'h	49a6;
40954	:douta	=	16'h	49a6;
40955	:douta	=	16'h	4985;
40956	:douta	=	16'h	4185;
40957	:douta	=	16'h	4186;
40958	:douta	=	16'h	4185;
40959	:douta	=	16'h	4165;
40960	:douta	=	16'h	eed7;
40961	:douta	=	16'h	f6f8;
40962	:douta	=	16'h	f71a;
40963	:douta	=	16'h	f6f9;
40964	:douta	=	16'h	f73a;
40965	:douta	=	16'h	ff3a;
40966	:douta	=	16'h	f6f9;
40967	:douta	=	16'h	ff19;
40968	:douta	=	16'h	ff3a;
40969	:douta	=	16'h	ff7b;
40970	:douta	=	16'h	ee97;
40971	:douta	=	16'h	bd96;
40972	:douta	=	16'h	ad16;
40973	:douta	=	16'h	9473;
40974	:douta	=	16'h	a516;
40975	:douta	=	16'h	94d5;
40976	:douta	=	16'h	9c94;
40977	:douta	=	16'h	9453;
40978	:douta	=	16'h	9cb4;
40979	:douta	=	16'h	9cd6;
40980	:douta	=	16'h	a516;
40981	:douta	=	16'h	8c75;
40982	:douta	=	16'h	7455;
40983	:douta	=	16'h	7c97;
40984	:douta	=	16'h	7cb7;
40985	:douta	=	16'h	7c77;
40986	:douta	=	16'h	7c76;
40987	:douta	=	16'h	7c96;
40988	:douta	=	16'h	7c76;
40989	:douta	=	16'h	84d8;
40990	:douta	=	16'h	3a6c;
40991	:douta	=	16'h	0042;
40992	:douta	=	16'h	1083;
40993	:douta	=	16'h	10e6;
40994	:douta	=	16'h	1947;
40995	:douta	=	16'h	1927;
40996	:douta	=	16'h	1927;
40997	:douta	=	16'h	1947;
40998	:douta	=	16'h	1906;
40999	:douta	=	16'h	1105;
41000	:douta	=	16'h	1105;
41001	:douta	=	16'h	1126;
41002	:douta	=	16'h	1947;
41003	:douta	=	16'h	2189;
41004	:douta	=	16'h	21a9;
41005	:douta	=	16'h	2189;
41006	:douta	=	16'h	2168;
41007	:douta	=	16'h	1927;
41008	:douta	=	16'h	10e4;
41009	:douta	=	16'h	21a8;
41010	:douta	=	16'h	2189;
41011	:douta	=	16'h	2188;
41012	:douta	=	16'h	2168;
41013	:douta	=	16'h	1926;
41014	:douta	=	16'h	2146;
41015	:douta	=	16'h	10c5;
41016	:douta	=	16'h	29a8;
41017	:douta	=	16'h	29a9;
41018	:douta	=	16'h	29ca;
41019	:douta	=	16'h	1061;
41020	:douta	=	16'h	18a2;
41021	:douta	=	16'h	0841;
41022	:douta	=	16'h	0000;
41023	:douta	=	16'h	2924;
41024	:douta	=	16'h	1882;
41025	:douta	=	16'h	1905;
41026	:douta	=	16'h	2967;
41027	:douta	=	16'h	31c9;
41028	:douta	=	16'h	29c9;
41029	:douta	=	16'h	3a0a;
41030	:douta	=	16'h	3a2b;
41031	:douta	=	16'h	31c9;
41032	:douta	=	16'h	3a0a;
41033	:douta	=	16'h	3a2b;
41034	:douta	=	16'h	39c9;
41035	:douta	=	16'h	31a8;
41036	:douta	=	16'h	39e9;
41037	:douta	=	16'h	3a0a;
41038	:douta	=	16'h	39e8;
41039	:douta	=	16'h	39c9;
41040	:douta	=	16'h	39e9;
41041	:douta	=	16'h	424a;
41042	:douta	=	16'h	424a;
41043	:douta	=	16'h	4a6b;
41044	:douta	=	16'h	52ac;
41045	:douta	=	16'h	4a8b;
41046	:douta	=	16'h	4aab;
41047	:douta	=	16'h	52ab;
41048	:douta	=	16'h	528b;
41049	:douta	=	16'h	52ac;
41050	:douta	=	16'h	634e;
41051	:douta	=	16'h	636f;
41052	:douta	=	16'h	6b90;
41053	:douta	=	16'h	6b8f;
41054	:douta	=	16'h	6b4e;
41055	:douta	=	16'h	738f;
41056	:douta	=	16'h	834b;
41057	:douta	=	16'h	7b29;
41058	:douta	=	16'h	8b27;
41059	:douta	=	16'h	9b47;
41060	:douta	=	16'h	b3a5;
41061	:douta	=	16'h	bbc4;
41062	:douta	=	16'h	c3e5;
41063	:douta	=	16'h	c3e3;
41064	:douta	=	16'h	bb83;
41065	:douta	=	16'h	bbc4;
41066	:douta	=	16'h	bbe4;
41067	:douta	=	16'h	bbe5;
41068	:douta	=	16'h	c3e5;
41069	:douta	=	16'h	c406;
41070	:douta	=	16'h	c403;
41071	:douta	=	16'h	c406;
41072	:douta	=	16'h	cc25;
41073	:douta	=	16'h	c406;
41074	:douta	=	16'h	c425;
41075	:douta	=	16'h	cc25;
41076	:douta	=	16'h	cc25;
41077	:douta	=	16'h	cc26;
41078	:douta	=	16'h	c425;
41079	:douta	=	16'h	c425;
41080	:douta	=	16'h	cc45;
41081	:douta	=	16'h	cc45;
41082	:douta	=	16'h	cc45;
41083	:douta	=	16'h	cc45;
41084	:douta	=	16'h	cc25;
41085	:douta	=	16'h	cc45;
41086	:douta	=	16'h	cc45;
41087	:douta	=	16'h	cc66;
41088	:douta	=	16'h	cc45;
41089	:douta	=	16'h	cc65;
41090	:douta	=	16'h	d445;
41091	:douta	=	16'h	cc66;
41092	:douta	=	16'h	cc66;
41093	:douta	=	16'h	cc66;
41094	:douta	=	16'h	cc66;
41095	:douta	=	16'h	d465;
41096	:douta	=	16'h	cc66;
41097	:douta	=	16'h	d467;
41098	:douta	=	16'h	d466;
41099	:douta	=	16'h	cc66;
41100	:douta	=	16'h	d466;
41101	:douta	=	16'h	cc66;
41102	:douta	=	16'h	cc65;
41103	:douta	=	16'h	cc66;
41104	:douta	=	16'h	d466;
41105	:douta	=	16'h	dc44;
41106	:douta	=	16'h	a42d;
41107	:douta	=	16'h	9410;
41108	:douta	=	16'h	9430;
41109	:douta	=	16'h	9411;
41110	:douta	=	16'h	9430;
41111	:douta	=	16'h	9cb3;
41112	:douta	=	16'h	9453;
41113	:douta	=	16'h	8bd0;
41114	:douta	=	16'h	83d0;
41115	:douta	=	16'h	7bb0;
41116	:douta	=	16'h	632f;
41117	:douta	=	16'h	52ac;
41118	:douta	=	16'h	acb0;
41119	:douta	=	16'h	e675;
41120	:douta	=	16'h	93cd;
41121	:douta	=	16'h	e6b8;
41122	:douta	=	16'h	b555;
41123	:douta	=	16'h	c574;
41124	:douta	=	16'h	e677;
41125	:douta	=	16'h	eeb7;
41126	:douta	=	16'h	c554;
41127	:douta	=	16'h	d5d6;
41128	:douta	=	16'h	c595;
41129	:douta	=	16'h	cd95;
41130	:douta	=	16'h	bd34;
41131	:douta	=	16'h	b515;
41132	:douta	=	16'h	9cb4;
41133	:douta	=	16'h	8c53;
41134	:douta	=	16'h	8c73;
41135	:douta	=	16'h	7bf2;
41136	:douta	=	16'h	73b1;
41137	:douta	=	16'h	8412;
41138	:douta	=	16'h	7bf1;
41139	:douta	=	16'h	8432;
41140	:douta	=	16'h	8c73;
41141	:douta	=	16'h	9494;
41142	:douta	=	16'h	7390;
41143	:douta	=	16'h	7370;
41144	:douta	=	16'h	6b50;
41145	:douta	=	16'h	632f;
41146	:douta	=	16'h	632f;
41147	:douta	=	16'h	41e7;
41148	:douta	=	16'h	4a08;
41149	:douta	=	16'h	5249;
41150	:douta	=	16'h	734b;
41151	:douta	=	16'h	83ac;
41152	:douta	=	16'h	93ed;
41153	:douta	=	16'h	ac90;
41154	:douta	=	16'h	cd72;
41155	:douta	=	16'h	de34;
41156	:douta	=	16'h	de14;
41157	:douta	=	16'h	e655;
41158	:douta	=	16'h	e656;
41159	:douta	=	16'h	de55;
41160	:douta	=	16'h	e656;
41161	:douta	=	16'h	de35;
41162	:douta	=	16'h	d5f4;
41163	:douta	=	16'h	d5f4;
41164	:douta	=	16'h	d5f4;
41165	:douta	=	16'h	d5d4;
41166	:douta	=	16'h	cd93;
41167	:douta	=	16'h	b535;
41168	:douta	=	16'h	a516;
41169	:douta	=	16'h	a516;
41170	:douta	=	16'h	94d5;
41171	:douta	=	16'h	94d5;
41172	:douta	=	16'h	8cb5;
41173	:douta	=	16'h	8475;
41174	:douta	=	16'h	7c54;
41175	:douta	=	16'h	7413;
41176	:douta	=	16'h	7413;
41177	:douta	=	16'h	6bd3;
41178	:douta	=	16'h	5330;
41179	:douta	=	16'h	5330;
41180	:douta	=	16'h	5b72;
41181	:douta	=	16'h	5b71;
41182	:douta	=	16'h	324b;
41183	:douta	=	16'h	4a8c;
41184	:douta	=	16'h	2968;
41185	:douta	=	16'h	2988;
41186	:douta	=	16'h	2127;
41187	:douta	=	16'h	1927;
41188	:douta	=	16'h	7a65;
41189	:douta	=	16'h	7245;
41190	:douta	=	16'h	7245;
41191	:douta	=	16'h	6a25;
41192	:douta	=	16'h	6a25;
41193	:douta	=	16'h	6205;
41194	:douta	=	16'h	6205;
41195	:douta	=	16'h	61e5;
41196	:douta	=	16'h	61e5;
41197	:douta	=	16'h	59e5;
41198	:douta	=	16'h	59c5;
41199	:douta	=	16'h	59e5;
41200	:douta	=	16'h	59e5;
41201	:douta	=	16'h	59c5;
41202	:douta	=	16'h	51c5;
41203	:douta	=	16'h	51c6;
41204	:douta	=	16'h	51c5;
41205	:douta	=	16'h	51c5;
41206	:douta	=	16'h	49c6;
41207	:douta	=	16'h	49a5;
41208	:douta	=	16'h	49a6;
41209	:douta	=	16'h	49a5;
41210	:douta	=	16'h	49a6;
41211	:douta	=	16'h	49a6;
41212	:douta	=	16'h	4185;
41213	:douta	=	16'h	4185;
41214	:douta	=	16'h	4185;
41215	:douta	=	16'h	4186;
41216	:douta	=	16'h	eed6;
41217	:douta	=	16'h	ff1a;
41218	:douta	=	16'h	f6f8;
41219	:douta	=	16'h	f6f9;
41220	:douta	=	16'h	ff19;
41221	:douta	=	16'h	f6f9;
41222	:douta	=	16'h	ff19;
41223	:douta	=	16'h	ff19;
41224	:douta	=	16'h	ff5a;
41225	:douta	=	16'h	eeb7;
41226	:douta	=	16'h	de15;
41227	:douta	=	16'h	ad16;
41228	:douta	=	16'h	a4d5;
41229	:douta	=	16'h	a516;
41230	:douta	=	16'h	a516;
41231	:douta	=	16'h	a516;
41232	:douta	=	16'h	9c94;
41233	:douta	=	16'h	a4d5;
41234	:douta	=	16'h	9cd5;
41235	:douta	=	16'h	9cd6;
41236	:douta	=	16'h	a516;
41237	:douta	=	16'h	6bf3;
41238	:douta	=	16'h	6bf3;
41239	:douta	=	16'h	7414;
41240	:douta	=	16'h	7435;
41241	:douta	=	16'h	7c96;
41242	:douta	=	16'h	7c96;
41243	:douta	=	16'h	8497;
41244	:douta	=	16'h	7c56;
41245	:douta	=	16'h	8497;
41246	:douta	=	16'h	8496;
41247	:douta	=	16'h	84f8;
41248	:douta	=	16'h	7434;
41249	:douta	=	16'h	29ca;
41250	:douta	=	16'h	10e5;
41251	:douta	=	16'h	1105;
41252	:douta	=	16'h	1927;
41253	:douta	=	16'h	1106;
41254	:douta	=	16'h	1926;
41255	:douta	=	16'h	1126;
41256	:douta	=	16'h	1105;
41257	:douta	=	16'h	10e5;
41258	:douta	=	16'h	1906;
41259	:douta	=	16'h	1126;
41260	:douta	=	16'h	1927;
41261	:douta	=	16'h	2147;
41262	:douta	=	16'h	1947;
41263	:douta	=	16'h	2188;
41264	:douta	=	16'h	21a8;
41265	:douta	=	16'h	10c4;
41266	:douta	=	16'h	10a4;
41267	:douta	=	16'h	2126;
41268	:douta	=	16'h	1926;
41269	:douta	=	16'h	3186;
41270	:douta	=	16'h	2126;
41271	:douta	=	16'h	10c5;
41272	:douta	=	16'h	2126;
41273	:douta	=	16'h	2126;
41274	:douta	=	16'h	2167;
41275	:douta	=	16'h	18a3;
41276	:douta	=	16'h	1081;
41277	:douta	=	16'h	1061;
41278	:douta	=	16'h	0841;
41279	:douta	=	16'h	18c4;
41280	:douta	=	16'h	2967;
41281	:douta	=	16'h	29a9;
41282	:douta	=	16'h	29a9;
41283	:douta	=	16'h	31ea;
41284	:douta	=	16'h	31e9;
41285	:douta	=	16'h	2968;
41286	:douta	=	16'h	2188;
41287	:douta	=	16'h	3a2a;
41288	:douta	=	16'h	29a8;
41289	:douta	=	16'h	3209;
41290	:douta	=	16'h	320a;
41291	:douta	=	16'h	424b;
41292	:douta	=	16'h	424b;
41293	:douta	=	16'h	422b;
41294	:douta	=	16'h	3a09;
41295	:douta	=	16'h	422a;
41296	:douta	=	16'h	422a;
41297	:douta	=	16'h	4acd;
41298	:douta	=	16'h	428c;
41299	:douta	=	16'h	4a8c;
41300	:douta	=	16'h	3a2a;
41301	:douta	=	16'h	52ab;
41302	:douta	=	16'h	62eb;
41303	:douta	=	16'h	6acb;
41304	:douta	=	16'h	72c9;
41305	:douta	=	16'h	7ac8;
41306	:douta	=	16'h	82c6;
41307	:douta	=	16'h	92c3;
41308	:douta	=	16'h	92c3;
41309	:douta	=	16'h	ab23;
41310	:douta	=	16'h	ab44;
41311	:douta	=	16'h	b384;
41312	:douta	=	16'h	b385;
41313	:douta	=	16'h	b385;
41314	:douta	=	16'h	b385;
41315	:douta	=	16'h	b3a5;
41316	:douta	=	16'h	b3a5;
41317	:douta	=	16'h	bba6;
41318	:douta	=	16'h	bba5;
41319	:douta	=	16'h	bbc4;
41320	:douta	=	16'h	bbc5;
41321	:douta	=	16'h	bbc5;
41322	:douta	=	16'h	c3e5;
41323	:douta	=	16'h	bbe5;
41324	:douta	=	16'h	c405;
41325	:douta	=	16'h	c405;
41326	:douta	=	16'h	c405;
41327	:douta	=	16'h	c404;
41328	:douta	=	16'h	c404;
41329	:douta	=	16'h	c404;
41330	:douta	=	16'h	cc05;
41331	:douta	=	16'h	cc46;
41332	:douta	=	16'h	cc25;
41333	:douta	=	16'h	cc25;
41334	:douta	=	16'h	cc25;
41335	:douta	=	16'h	cc45;
41336	:douta	=	16'h	cc45;
41337	:douta	=	16'h	cc25;
41338	:douta	=	16'h	cc45;
41339	:douta	=	16'h	cc45;
41340	:douta	=	16'h	cc45;
41341	:douta	=	16'h	cc45;
41342	:douta	=	16'h	cc46;
41343	:douta	=	16'h	cc45;
41344	:douta	=	16'h	cc45;
41345	:douta	=	16'h	cc46;
41346	:douta	=	16'h	cc66;
41347	:douta	=	16'h	d466;
41348	:douta	=	16'h	d445;
41349	:douta	=	16'h	cc46;
41350	:douta	=	16'h	cc66;
41351	:douta	=	16'h	d445;
41352	:douta	=	16'h	d444;
41353	:douta	=	16'h	d421;
41354	:douta	=	16'h	cc21;
41355	:douta	=	16'h	cc22;
41356	:douta	=	16'h	cc45;
41357	:douta	=	16'h	d4a9;
41358	:douta	=	16'h	d50b;
41359	:douta	=	16'h	ddaf;
41360	:douta	=	16'h	ddf1;
41361	:douta	=	16'h	eeb5;
41362	:douta	=	16'h	ef39;
41363	:douta	=	16'h	ff9a;
41364	:douta	=	16'h	e6f8;
41365	:douta	=	16'h	c5f5;
41366	:douta	=	16'h	8bcf;
41367	:douta	=	16'h	836e;
41368	:douta	=	16'h	834d;
41369	:douta	=	16'h	730c;
41370	:douta	=	16'h	7b6d;
41371	:douta	=	16'h	a490;
41372	:douta	=	16'h	d5b2;
41373	:douta	=	16'h	e656;
41374	:douta	=	16'h	e677;
41375	:douta	=	16'h	cdb3;
41376	:douta	=	16'h	f6f8;
41377	:douta	=	16'h	9cd6;
41378	:douta	=	16'h	bd97;
41379	:douta	=	16'h	cdd6;
41380	:douta	=	16'h	d616;
41381	:douta	=	16'h	b597;
41382	:douta	=	16'h	94b6;
41383	:douta	=	16'h	9cd6;
41384	:douta	=	16'h	a516;
41385	:douta	=	16'h	9cd5;
41386	:douta	=	16'h	9cb4;
41387	:douta	=	16'h	9cb4;
41388	:douta	=	16'h	8433;
41389	:douta	=	16'h	8c33;
41390	:douta	=	16'h	8412;
41391	:douta	=	16'h	7390;
41392	:douta	=	16'h	6b90;
41393	:douta	=	16'h	7390;
41394	:douta	=	16'h	8412;
41395	:douta	=	16'h	7bd0;
41396	:douta	=	16'h	6b6f;
41397	:douta	=	16'h	73b0;
41398	:douta	=	16'h	7390;
41399	:douta	=	16'h	5aac;
41400	:douta	=	16'h	4a08;
41401	:douta	=	16'h	49e7;
41402	:douta	=	16'h	5248;
41403	:douta	=	16'h	9c4f;
41404	:douta	=	16'h	bd0f;
41405	:douta	=	16'h	c550;
41406	:douta	=	16'h	d5f2;
41407	:douta	=	16'h	e635;
41408	:douta	=	16'h	e676;
41409	:douta	=	16'h	cdb2;
41410	:douta	=	16'h	c572;
41411	:douta	=	16'h	d5d4;
41412	:douta	=	16'h	de35;
41413	:douta	=	16'h	d5f4;
41414	:douta	=	16'h	ddd4;
41415	:douta	=	16'h	ddf5;
41416	:douta	=	16'h	d5d5;
41417	:douta	=	16'h	cdb5;
41418	:douta	=	16'h	c555;
41419	:douta	=	16'h	acd4;
41420	:douta	=	16'h	acd4;
41421	:douta	=	16'h	a4d5;
41422	:douta	=	16'h	a4d5;
41423	:douta	=	16'h	9cf5;
41424	:douta	=	16'h	9cf6;
41425	:douta	=	16'h	9cf5;
41426	:douta	=	16'h	94f6;
41427	:douta	=	16'h	94d5;
41428	:douta	=	16'h	8c75;
41429	:douta	=	16'h	7c34;
41430	:douta	=	16'h	7c54;
41431	:douta	=	16'h	7434;
41432	:douta	=	16'h	7434;
41433	:douta	=	16'h	6bf3;
41434	:douta	=	16'h	6392;
41435	:douta	=	16'h	5330;
41436	:douta	=	16'h	322c;
41437	:douta	=	16'h	3a2b;
41438	:douta	=	16'h	4acf;
41439	:douta	=	16'h	73f1;
41440	:douta	=	16'h	634f;
41441	:douta	=	16'h	2147;
41442	:douta	=	16'h	2126;
41443	:douta	=	16'h	2948;
41444	:douta	=	16'h	1906;
41445	:douta	=	16'h	6a46;
41446	:douta	=	16'h	6a25;
41447	:douta	=	16'h	6a25;
41448	:douta	=	16'h	6a05;
41449	:douta	=	16'h	6a25;
41450	:douta	=	16'h	6a05;
41451	:douta	=	16'h	61e5;
41452	:douta	=	16'h	61e5;
41453	:douta	=	16'h	61e5;
41454	:douta	=	16'h	59e5;
41455	:douta	=	16'h	59e5;
41456	:douta	=	16'h	59c5;
41457	:douta	=	16'h	59e6;
41458	:douta	=	16'h	51c5;
41459	:douta	=	16'h	51a5;
41460	:douta	=	16'h	51c5;
41461	:douta	=	16'h	51c6;
41462	:douta	=	16'h	51c6;
41463	:douta	=	16'h	49c6;
41464	:douta	=	16'h	49a6;
41465	:douta	=	16'h	49a6;
41466	:douta	=	16'h	49a6;
41467	:douta	=	16'h	4185;
41468	:douta	=	16'h	4186;
41469	:douta	=	16'h	4186;
41470	:douta	=	16'h	4186;
41471	:douta	=	16'h	4186;
41472	:douta	=	16'h	f6f8;
41473	:douta	=	16'h	f6f9;
41474	:douta	=	16'h	f6f8;
41475	:douta	=	16'h	f719;
41476	:douta	=	16'h	ff19;
41477	:douta	=	16'h	f719;
41478	:douta	=	16'h	ff19;
41479	:douta	=	16'h	ff19;
41480	:douta	=	16'h	ff7b;
41481	:douta	=	16'h	d5f5;
41482	:douta	=	16'h	d5d5;
41483	:douta	=	16'h	ad16;
41484	:douta	=	16'h	9cb4;
41485	:douta	=	16'h	a537;
41486	:douta	=	16'h	9cd5;
41487	:douta	=	16'h	a516;
41488	:douta	=	16'h	9cb4;
41489	:douta	=	16'h	a4b4;
41490	:douta	=	16'h	9cf5;
41491	:douta	=	16'h	a516;
41492	:douta	=	16'h	a516;
41493	:douta	=	16'h	6bf3;
41494	:douta	=	16'h	6bf3;
41495	:douta	=	16'h	7414;
41496	:douta	=	16'h	73f4;
41497	:douta	=	16'h	7435;
41498	:douta	=	16'h	7c76;
41499	:douta	=	16'h	8497;
41500	:douta	=	16'h	7c76;
41501	:douta	=	16'h	8497;
41502	:douta	=	16'h	8476;
41503	:douta	=	16'h	7c76;
41504	:douta	=	16'h	8497;
41505	:douta	=	16'h	8d39;
41506	:douta	=	16'h	0884;
41507	:douta	=	16'h	10c5;
41508	:douta	=	16'h	10c5;
41509	:douta	=	16'h	10e5;
41510	:douta	=	16'h	1105;
41511	:douta	=	16'h	1105;
41512	:douta	=	16'h	08c5;
41513	:douta	=	16'h	10e5;
41514	:douta	=	16'h	10e5;
41515	:douta	=	16'h	1906;
41516	:douta	=	16'h	1926;
41517	:douta	=	16'h	1105;
41518	:douta	=	16'h	1926;
41519	:douta	=	16'h	1927;
41520	:douta	=	16'h	2147;
41521	:douta	=	16'h	2126;
41522	:douta	=	16'h	18e5;
41523	:douta	=	16'h	10c4;
41524	:douta	=	16'h	18c4;
41525	:douta	=	16'h	10c3;
41526	:douta	=	16'h	2126;
41527	:douta	=	16'h	10c5;
41528	:douta	=	16'h	2126;
41529	:douta	=	16'h	1905;
41530	:douta	=	16'h	2146;
41531	:douta	=	16'h	2147;
41532	:douta	=	16'h	20e5;
41533	:douta	=	16'h	20e3;
41534	:douta	=	16'h	1083;
41535	:douta	=	16'h	2145;
41536	:douta	=	16'h	320b;
41537	:douta	=	16'h	322b;
41538	:douta	=	16'h	3a2c;
41539	:douta	=	16'h	3a2c;
41540	:douta	=	16'h	320a;
41541	:douta	=	16'h	424b;
41542	:douta	=	16'h	3a2b;
41543	:douta	=	16'h	4aad;
41544	:douta	=	16'h	4ace;
41545	:douta	=	16'h	42ae;
41546	:douta	=	16'h	4ace;
41547	:douta	=	16'h	426c;
41548	:douta	=	16'h	3a2a;
41549	:douta	=	16'h	320a;
41550	:douta	=	16'h	3a2b;
41551	:douta	=	16'h	4a8c;
41552	:douta	=	16'h	4aac;
41553	:douta	=	16'h	52ab;
41554	:douta	=	16'h	62cb;
41555	:douta	=	16'h	6aea;
41556	:douta	=	16'h	6267;
41557	:douta	=	16'h	7266;
41558	:douta	=	16'h	8263;
41559	:douta	=	16'h	8283;
41560	:douta	=	16'h	8aa2;
41561	:douta	=	16'h	92c2;
41562	:douta	=	16'h	9ac2;
41563	:douta	=	16'h	a325;
41564	:douta	=	16'h	a345;
41565	:douta	=	16'h	ab64;
41566	:douta	=	16'h	ab84;
41567	:douta	=	16'h	ab64;
41568	:douta	=	16'h	b365;
41569	:douta	=	16'h	b385;
41570	:douta	=	16'h	b3a5;
41571	:douta	=	16'h	b3a5;
41572	:douta	=	16'h	b3c5;
41573	:douta	=	16'h	bba5;
41574	:douta	=	16'h	b3c4;
41575	:douta	=	16'h	bbe5;
41576	:douta	=	16'h	bbc6;
41577	:douta	=	16'h	bbe5;
41578	:douta	=	16'h	bbe5;
41579	:douta	=	16'h	c3e5;
41580	:douta	=	16'h	c405;
41581	:douta	=	16'h	c405;
41582	:douta	=	16'h	c425;
41583	:douta	=	16'h	cc05;
41584	:douta	=	16'h	c406;
41585	:douta	=	16'h	cc25;
41586	:douta	=	16'h	cc25;
41587	:douta	=	16'h	cc46;
41588	:douta	=	16'h	cc47;
41589	:douta	=	16'h	cc26;
41590	:douta	=	16'h	cc46;
41591	:douta	=	16'h	cc66;
41592	:douta	=	16'h	cc25;
41593	:douta	=	16'h	cc45;
41594	:douta	=	16'h	cc25;
41595	:douta	=	16'h	cc46;
41596	:douta	=	16'h	cc45;
41597	:douta	=	16'h	cc45;
41598	:douta	=	16'h	cc45;
41599	:douta	=	16'h	cc46;
41600	:douta	=	16'h	cc44;
41601	:douta	=	16'h	cc65;
41602	:douta	=	16'h	cc45;
41603	:douta	=	16'h	cc24;
41604	:douta	=	16'h	cc02;
41605	:douta	=	16'h	cc20;
41606	:douta	=	16'h	cc00;
41607	:douta	=	16'h	cc44;
41608	:douta	=	16'h	cc87;
41609	:douta	=	16'h	d4ea;
41610	:douta	=	16'h	d56e;
41611	:douta	=	16'h	e5d0;
41612	:douta	=	16'h	e694;
41613	:douta	=	16'h	ef38;
41614	:douta	=	16'h	f77a;
41615	:douta	=	16'h	ffbc;
41616	:douta	=	16'h	f7dc;
41617	:douta	=	16'h	f779;
41618	:douta	=	16'h	f6f6;
41619	:douta	=	16'h	e693;
41620	:douta	=	16'h	f650;
41621	:douta	=	16'h	ee2f;
41622	:douta	=	16'h	bc29;
41623	:douta	=	16'h	a3ca;
41624	:douta	=	16'h	ac6f;
41625	:douta	=	16'h	940e;
41626	:douta	=	16'h	d5d4;
41627	:douta	=	16'h	de14;
41628	:douta	=	16'h	e656;
41629	:douta	=	16'h	e677;
41630	:douta	=	16'h	de36;
41631	:douta	=	16'h	d5f5;
41632	:douta	=	16'h	eeb7;
41633	:douta	=	16'h	94d6;
41634	:douta	=	16'h	bd76;
41635	:douta	=	16'h	c5d7;
41636	:douta	=	16'h	cdd7;
41637	:douta	=	16'h	a557;
41638	:douta	=	16'h	8c96;
41639	:douta	=	16'h	8454;
41640	:douta	=	16'h	94b5;
41641	:douta	=	16'h	8c74;
41642	:douta	=	16'h	8453;
41643	:douta	=	16'h	8c53;
41644	:douta	=	16'h	8412;
41645	:douta	=	16'h	7bf2;
41646	:douta	=	16'h	8412;
41647	:douta	=	16'h	6b6f;
41648	:douta	=	16'h	6b6f;
41649	:douta	=	16'h	6b4f;
41650	:douta	=	16'h	6b2f;
41651	:douta	=	16'h	73b0;
41652	:douta	=	16'h	6b70;
41653	:douta	=	16'h	7390;
41654	:douta	=	16'h	524a;
41655	:douta	=	16'h	41c6;
41656	:douta	=	16'h	5228;
41657	:douta	=	16'h	83cd;
41658	:douta	=	16'h	9c4e;
41659	:douta	=	16'h	c530;
41660	:douta	=	16'h	cd91;
41661	:douta	=	16'h	d5d3;
41662	:douta	=	16'h	d5f4;
41663	:douta	=	16'h	e655;
41664	:douta	=	16'h	c533;
41665	:douta	=	16'h	e676;
41666	:douta	=	16'h	cd93;
41667	:douta	=	16'h	d5b3;
41668	:douta	=	16'h	d5d4;
41669	:douta	=	16'h	d5b4;
41670	:douta	=	16'h	d5b3;
41671	:douta	=	16'h	d5b4;
41672	:douta	=	16'h	bd34;
41673	:douta	=	16'h	bd34;
41674	:douta	=	16'h	bd75;
41675	:douta	=	16'h	9cb3;
41676	:douta	=	16'h	9cb3;
41677	:douta	=	16'h	a4b5;
41678	:douta	=	16'h	9cd5;
41679	:douta	=	16'h	9cf5;
41680	:douta	=	16'h	9d16;
41681	:douta	=	16'h	94f6;
41682	:douta	=	16'h	8cb5;
41683	:douta	=	16'h	8cd5;
41684	:douta	=	16'h	8c95;
41685	:douta	=	16'h	7c34;
41686	:douta	=	16'h	7c54;
41687	:douta	=	16'h	7434;
41688	:douta	=	16'h	7434;
41689	:douta	=	16'h	7434;
41690	:douta	=	16'h	7c75;
41691	:douta	=	16'h	7414;
41692	:douta	=	16'h	63b2;
41693	:douta	=	16'h	5b72;
41694	:douta	=	16'h	52ef;
41695	:douta	=	16'h	31a7;
41696	:douta	=	16'h	7b90;
41697	:douta	=	16'h	1906;
41698	:douta	=	16'h	2127;
41699	:douta	=	16'h	1926;
41700	:douta	=	16'h	08c5;
41701	:douta	=	16'h	41a5;
41702	:douta	=	16'h	7245;
41703	:douta	=	16'h	6a25;
41704	:douta	=	16'h	6a25;
41705	:douta	=	16'h	6a05;
41706	:douta	=	16'h	61e5;
41707	:douta	=	16'h	59e5;
41708	:douta	=	16'h	61e5;
41709	:douta	=	16'h	6206;
41710	:douta	=	16'h	59e5;
41711	:douta	=	16'h	59e5;
41712	:douta	=	16'h	59c5;
41713	:douta	=	16'h	59e6;
41714	:douta	=	16'h	51c5;
41715	:douta	=	16'h	51c5;
41716	:douta	=	16'h	51c5;
41717	:douta	=	16'h	51c6;
41718	:douta	=	16'h	51c5;
41719	:douta	=	16'h	49a5;
41720	:douta	=	16'h	49a6;
41721	:douta	=	16'h	49a5;
41722	:douta	=	16'h	4986;
41723	:douta	=	16'h	49a6;
41724	:douta	=	16'h	4185;
41725	:douta	=	16'h	4166;
41726	:douta	=	16'h	4186;
41727	:douta	=	16'h	3966;
41728	:douta	=	16'h	ff19;
41729	:douta	=	16'h	f6d8;
41730	:douta	=	16'h	f6d8;
41731	:douta	=	16'h	ff19;
41732	:douta	=	16'h	ff19;
41733	:douta	=	16'h	f739;
41734	:douta	=	16'h	f719;
41735	:douta	=	16'h	ff19;
41736	:douta	=	16'h	ff9b;
41737	:douta	=	16'h	d593;
41738	:douta	=	16'h	cdb6;
41739	:douta	=	16'h	a4d5;
41740	:douta	=	16'h	9473;
41741	:douta	=	16'h	a536;
41742	:douta	=	16'h	a516;
41743	:douta	=	16'h	a4f5;
41744	:douta	=	16'h	a4d4;
41745	:douta	=	16'h	9cb4;
41746	:douta	=	16'h	9cf5;
41747	:douta	=	16'h	9cd5;
41748	:douta	=	16'h	8c95;
41749	:douta	=	16'h	7414;
41750	:douta	=	16'h	7414;
41751	:douta	=	16'h	7434;
41752	:douta	=	16'h	7c55;
41753	:douta	=	16'h	7435;
41754	:douta	=	16'h	7c35;
41755	:douta	=	16'h	7c76;
41756	:douta	=	16'h	84d7;
41757	:douta	=	16'h	8497;
41758	:douta	=	16'h	7c76;
41759	:douta	=	16'h	73f3;
41760	:douta	=	16'h	6bf4;
41761	:douta	=	16'h	6c35;
41762	:douta	=	16'h	0883;
41763	:douta	=	16'h	10c5;
41764	:douta	=	16'h	08a5;
41765	:douta	=	16'h	10e5;
41766	:douta	=	16'h	10e5;
41767	:douta	=	16'h	10e5;
41768	:douta	=	16'h	10c5;
41769	:douta	=	16'h	10e5;
41770	:douta	=	16'h	10e5;
41771	:douta	=	16'h	10e5;
41772	:douta	=	16'h	10c5;
41773	:douta	=	16'h	10c4;
41774	:douta	=	16'h	1105;
41775	:douta	=	16'h	1906;
41776	:douta	=	16'h	1905;
41777	:douta	=	16'h	10e5;
41778	:douta	=	16'h	18e5;
41779	:douta	=	16'h	18e5;
41780	:douta	=	16'h	2125;
41781	:douta	=	16'h	18e4;
41782	:douta	=	16'h	2106;
41783	:douta	=	16'h	10e4;
41784	:douta	=	16'h	18e5;
41785	:douta	=	16'h	1926;
41786	:douta	=	16'h	18e5;
41787	:douta	=	16'h	2125;
41788	:douta	=	16'h	2167;
41789	:douta	=	16'h	29a9;
41790	:douta	=	16'h	18e4;
41791	:douta	=	16'h	31ea;
41792	:douta	=	16'h	324c;
41793	:douta	=	16'h	322b;
41794	:douta	=	16'h	3a6c;
41795	:douta	=	16'h	3a2c;
41796	:douta	=	16'h	3a6c;
41797	:douta	=	16'h	322b;
41798	:douta	=	16'h	3a4c;
41799	:douta	=	16'h	42ce;
41800	:douta	=	16'h	42ad;
41801	:douta	=	16'h	4a4a;
41802	:douta	=	16'h	51a5;
41803	:douta	=	16'h	51a5;
41804	:douta	=	16'h	59e4;
41805	:douta	=	16'h	61e4;
41806	:douta	=	16'h	61a3;
41807	:douta	=	16'h	69e3;
41808	:douta	=	16'h	7203;
41809	:douta	=	16'h	7a24;
41810	:douta	=	16'h	7a44;
41811	:douta	=	16'h	8aa4;
41812	:douta	=	16'h	8ac4;
41813	:douta	=	16'h	92c4;
41814	:douta	=	16'h	92e4;
41815	:douta	=	16'h	92e4;
41816	:douta	=	16'h	9b04;
41817	:douta	=	16'h	9b05;
41818	:douta	=	16'h	9b04;
41819	:douta	=	16'h	a345;
41820	:douta	=	16'h	a344;
41821	:douta	=	16'h	ab65;
41822	:douta	=	16'h	ab64;
41823	:douta	=	16'h	ab85;
41824	:douta	=	16'h	b385;
41825	:douta	=	16'h	b385;
41826	:douta	=	16'h	ab84;
41827	:douta	=	16'h	b384;
41828	:douta	=	16'h	b3a5;
41829	:douta	=	16'h	bba5;
41830	:douta	=	16'h	bbc5;
41831	:douta	=	16'h	bbc5;
41832	:douta	=	16'h	bbc6;
41833	:douta	=	16'h	bbe5;
41834	:douta	=	16'h	c3e5;
41835	:douta	=	16'h	c3e5;
41836	:douta	=	16'h	c405;
41837	:douta	=	16'h	c425;
41838	:douta	=	16'h	c426;
41839	:douta	=	16'h	c426;
41840	:douta	=	16'h	cc46;
41841	:douta	=	16'h	d467;
41842	:douta	=	16'h	cc46;
41843	:douta	=	16'h	cc25;
41844	:douta	=	16'h	cc25;
41845	:douta	=	16'h	cc45;
41846	:douta	=	16'h	cc25;
41847	:douta	=	16'h	cc25;
41848	:douta	=	16'h	cc25;
41849	:douta	=	16'h	cc24;
41850	:douta	=	16'h	cc04;
41851	:douta	=	16'h	c3e2;
41852	:douta	=	16'h	c3e1;
41853	:douta	=	16'h	cc24;
41854	:douta	=	16'h	cc66;
41855	:douta	=	16'h	cca8;
41856	:douta	=	16'h	dd6e;
41857	:douta	=	16'h	ddae;
41858	:douta	=	16'h	e633;
41859	:douta	=	16'h	eed7;
41860	:douta	=	16'h	ef39;
41861	:douta	=	16'h	f7bc;
41862	:douta	=	16'h	ffdc;
41863	:douta	=	16'h	f7bb;
41864	:douta	=	16'h	f738;
41865	:douta	=	16'h	eed6;
41866	:douta	=	16'h	e611;
41867	:douta	=	16'h	ddaf;
41868	:douta	=	16'h	d50a;
41869	:douta	=	16'h	d487;
41870	:douta	=	16'h	cc65;
41871	:douta	=	16'h	cc22;
41872	:douta	=	16'h	cc02;
41873	:douta	=	16'h	d425;
41874	:douta	=	16'h	cc45;
41875	:douta	=	16'h	d466;
41876	:douta	=	16'h	d467;
41877	:douta	=	16'h	d466;
41878	:douta	=	16'h	d486;
41879	:douta	=	16'h	d466;
41880	:douta	=	16'h	d443;
41881	:douta	=	16'h	bd95;
41882	:douta	=	16'h	d5d6;
41883	:douta	=	16'h	d5d5;
41884	:douta	=	16'h	d5f5;
41885	:douta	=	16'h	cdb5;
41886	:douta	=	16'h	de56;
41887	:douta	=	16'h	de35;
41888	:douta	=	16'h	bd97;
41889	:douta	=	16'h	a537;
41890	:douta	=	16'h	ad77;
41891	:douta	=	16'h	bd98;
41892	:douta	=	16'h	b598;
41893	:douta	=	16'h	94b5;
41894	:douta	=	16'h	8453;
41895	:douta	=	16'h	7bf2;
41896	:douta	=	16'h	73b1;
41897	:douta	=	16'h	7bd1;
41898	:douta	=	16'h	73d0;
41899	:douta	=	16'h	7b90;
41900	:douta	=	16'h	6b6f;
41901	:douta	=	16'h	7b70;
41902	:douta	=	16'h	734e;
41903	:douta	=	16'h	630e;
41904	:douta	=	16'h	632e;
41905	:douta	=	16'h	6b6f;
41906	:douta	=	16'h	630e;
41907	:douta	=	16'h	4a49;
41908	:douta	=	16'h	49c6;
41909	:douta	=	16'h	49e7;
41910	:douta	=	16'h	7bad;
41911	:douta	=	16'h	c571;
41912	:douta	=	16'h	c571;
41913	:douta	=	16'h	d5d3;
41914	:douta	=	16'h	de14;
41915	:douta	=	16'h	de56;
41916	:douta	=	16'h	e656;
41917	:douta	=	16'h	de55;
41918	:douta	=	16'h	de36;
41919	:douta	=	16'h	de55;
41920	:douta	=	16'h	cdd4;
41921	:douta	=	16'h	a4b3;
41922	:douta	=	16'h	de36;
41923	:douta	=	16'h	de56;
41924	:douta	=	16'h	cdd4;
41925	:douta	=	16'h	bd34;
41926	:douta	=	16'h	b514;
41927	:douta	=	16'h	bd14;
41928	:douta	=	16'h	9493;
41929	:douta	=	16'h	9493;
41930	:douta	=	16'h	9c94;
41931	:douta	=	16'h	8c93;
41932	:douta	=	16'h	94b4;
41933	:douta	=	16'h	8c93;
41934	:douta	=	16'h	9493;
41935	:douta	=	16'h	7c32;
41936	:douta	=	16'h	7c33;
41937	:douta	=	16'h	7c13;
41938	:douta	=	16'h	7c33;
41939	:douta	=	16'h	7c33;
41940	:douta	=	16'h	8454;
41941	:douta	=	16'h	7c13;
41942	:douta	=	16'h	73f2;
41943	:douta	=	16'h	6bf2;
41944	:douta	=	16'h	6bf2;
41945	:douta	=	16'h	6b91;
41946	:douta	=	16'h	6bf2;
41947	:douta	=	16'h	6b91;
41948	:douta	=	16'h	3165;
41949	:douta	=	16'h	41a7;
41950	:douta	=	16'h	52cd;
41951	:douta	=	16'h	428d;
41952	:douta	=	16'h	29a9;
41953	:douta	=	16'h	5b0f;
41954	:douta	=	16'h	10c5;
41955	:douta	=	16'h	10e5;
41956	:douta	=	16'h	18e5;
41957	:douta	=	16'h	08a5;
41958	:douta	=	16'h	8a85;
41959	:douta	=	16'h	7245;
41960	:douta	=	16'h	6225;
41961	:douta	=	16'h	6205;
41962	:douta	=	16'h	6a05;
41963	:douta	=	16'h	6205;
41964	:douta	=	16'h	6205;
41965	:douta	=	16'h	59e5;
41966	:douta	=	16'h	59e5;
41967	:douta	=	16'h	5a05;
41968	:douta	=	16'h	59c5;
41969	:douta	=	16'h	51c5;
41970	:douta	=	16'h	51c5;
41971	:douta	=	16'h	51c6;
41972	:douta	=	16'h	51c6;
41973	:douta	=	16'h	49a5;
41974	:douta	=	16'h	49a6;
41975	:douta	=	16'h	49a6;
41976	:douta	=	16'h	49a6;
41977	:douta	=	16'h	49a5;
41978	:douta	=	16'h	49a6;
41979	:douta	=	16'h	4185;
41980	:douta	=	16'h	41a6;
41981	:douta	=	16'h	4186;
41982	:douta	=	16'h	4166;
41983	:douta	=	16'h	4166;
41984	:douta	=	16'h	f719;
41985	:douta	=	16'h	f6f8;
41986	:douta	=	16'h	f6d8;
41987	:douta	=	16'h	ff19;
41988	:douta	=	16'h	f6f8;
41989	:douta	=	16'h	f719;
41990	:douta	=	16'h	f73a;
41991	:douta	=	16'h	f719;
41992	:douta	=	16'h	ef18;
41993	:douta	=	16'h	d5d4;
41994	:douta	=	16'h	c575;
41995	:douta	=	16'h	9c94;
41996	:douta	=	16'h	9c93;
41997	:douta	=	16'h	a516;
41998	:douta	=	16'h	a4f5;
41999	:douta	=	16'h	a4d5;
42000	:douta	=	16'h	a4f5;
42001	:douta	=	16'h	a4b4;
42002	:douta	=	16'h	9cf5;
42003	:douta	=	16'h	9cd5;
42004	:douta	=	16'h	7c54;
42005	:douta	=	16'h	73f3;
42006	:douta	=	16'h	7c34;
42007	:douta	=	16'h	7414;
42008	:douta	=	16'h	7c35;
42009	:douta	=	16'h	7c55;
42010	:douta	=	16'h	8496;
42011	:douta	=	16'h	7c35;
42012	:douta	=	16'h	8cd7;
42013	:douta	=	16'h	7c76;
42014	:douta	=	16'h	7c75;
42015	:douta	=	16'h	7c55;
42016	:douta	=	16'h	8476;
42017	:douta	=	16'h	3a4c;
42018	:douta	=	16'h	10c4;
42019	:douta	=	16'h	10e5;
42020	:douta	=	16'h	10c4;
42021	:douta	=	16'h	10c5;
42022	:douta	=	16'h	10c5;
42023	:douta	=	16'h	1106;
42024	:douta	=	16'h	1106;
42025	:douta	=	16'h	10e5;
42026	:douta	=	16'h	1106;
42027	:douta	=	16'h	10e5;
42028	:douta	=	16'h	10c5;
42029	:douta	=	16'h	10e5;
42030	:douta	=	16'h	1906;
42031	:douta	=	16'h	10a4;
42032	:douta	=	16'h	10e4;
42033	:douta	=	16'h	10e5;
42034	:douta	=	16'h	1905;
42035	:douta	=	16'h	18c4;
42036	:douta	=	16'h	1905;
42037	:douta	=	16'h	2126;
42038	:douta	=	16'h	1906;
42039	:douta	=	16'h	18e5;
42040	:douta	=	16'h	1906;
42041	:douta	=	16'h	2126;
42042	:douta	=	16'h	2167;
42043	:douta	=	16'h	1926;
42044	:douta	=	16'h	2988;
42045	:douta	=	16'h	31ea;
42046	:douta	=	16'h	1905;
42047	:douta	=	16'h	322b;
42048	:douta	=	16'h	3a6c;
42049	:douta	=	16'h	3a6c;
42050	:douta	=	16'h	3a8e;
42051	:douta	=	16'h	430f;
42052	:douta	=	16'h	3a4c;
42053	:douta	=	16'h	426c;
42054	:douta	=	16'h	4a4b;
42055	:douta	=	16'h	4a07;
42056	:douta	=	16'h	51e6;
42057	:douta	=	16'h	59c4;
42058	:douta	=	16'h	61e3;
42059	:douta	=	16'h	61e3;
42060	:douta	=	16'h	59a2;
42061	:douta	=	16'h	61c3;
42062	:douta	=	16'h	69e3;
42063	:douta	=	16'h	7a44;
42064	:douta	=	16'h	7a64;
42065	:douta	=	16'h	8284;
42066	:douta	=	16'h	8284;
42067	:douta	=	16'h	8aa4;
42068	:douta	=	16'h	8aa3;
42069	:douta	=	16'h	8ac3;
42070	:douta	=	16'h	92e4;
42071	:douta	=	16'h	92e4;
42072	:douta	=	16'h	9b04;
42073	:douta	=	16'h	9b04;
42074	:douta	=	16'h	9b05;
42075	:douta	=	16'h	a345;
42076	:douta	=	16'h	a345;
42077	:douta	=	16'h	a344;
42078	:douta	=	16'h	ab64;
42079	:douta	=	16'h	ab64;
42080	:douta	=	16'h	b385;
42081	:douta	=	16'h	ab85;
42082	:douta	=	16'h	b3a4;
42083	:douta	=	16'h	b385;
42084	:douta	=	16'h	b3c5;
42085	:douta	=	16'h	b3a5;
42086	:douta	=	16'h	bbc5;
42087	:douta	=	16'h	bbc4;
42088	:douta	=	16'h	bbe5;
42089	:douta	=	16'h	bbc5;
42090	:douta	=	16'h	bbe5;
42091	:douta	=	16'h	c3e5;
42092	:douta	=	16'h	c3e6;
42093	:douta	=	16'h	c406;
42094	:douta	=	16'h	c405;
42095	:douta	=	16'h	c405;
42096	:douta	=	16'h	c405;
42097	:douta	=	16'h	c426;
42098	:douta	=	16'h	cc06;
42099	:douta	=	16'h	cc25;
42100	:douta	=	16'h	c404;
42101	:douta	=	16'h	c3e3;
42102	:douta	=	16'h	c3c2;
42103	:douta	=	16'h	c3c2;
42104	:douta	=	16'h	c3c2;
42105	:douta	=	16'h	cc25;
42106	:douta	=	16'h	cc67;
42107	:douta	=	16'h	d4eb;
42108	:douta	=	16'h	d52d;
42109	:douta	=	16'h	e5f1;
42110	:douta	=	16'h	e6b5;
42111	:douta	=	16'h	eef8;
42112	:douta	=	16'h	f79b;
42113	:douta	=	16'h	f7bc;
42114	:douta	=	16'h	ffbc;
42115	:douta	=	16'h	f759;
42116	:douta	=	16'h	f717;
42117	:douta	=	16'h	ee73;
42118	:douta	=	16'h	de11;
42119	:douta	=	16'h	dd6d;
42120	:douta	=	16'h	d4c9;
42121	:douta	=	16'h	d486;
42122	:douta	=	16'h	cc22;
42123	:douta	=	16'h	cc02;
42124	:douta	=	16'h	cc04;
42125	:douta	=	16'h	d445;
42126	:douta	=	16'h	d446;
42127	:douta	=	16'h	d467;
42128	:douta	=	16'h	d467;
42129	:douta	=	16'h	d486;
42130	:douta	=	16'h	d466;
42131	:douta	=	16'h	d467;
42132	:douta	=	16'h	d467;
42133	:douta	=	16'h	d466;
42134	:douta	=	16'h	cc86;
42135	:douta	=	16'h	d487;
42136	:douta	=	16'h	d466;
42137	:douta	=	16'h	ac6f;
42138	:douta	=	16'h	b514;
42139	:douta	=	16'h	c595;
42140	:douta	=	16'h	cdd7;
42141	:douta	=	16'h	c576;
42142	:douta	=	16'h	d5d7;
42143	:douta	=	16'h	cdd6;
42144	:douta	=	16'h	b577;
42145	:douta	=	16'h	ad57;
42146	:douta	=	16'h	ad77;
42147	:douta	=	16'h	bd97;
42148	:douta	=	16'h	94d6;
42149	:douta	=	16'h	8c73;
42150	:douta	=	16'h	8412;
42151	:douta	=	16'h	7bf2;
42152	:douta	=	16'h	6b70;
42153	:douta	=	16'h	73b0;
42154	:douta	=	16'h	7390;
42155	:douta	=	16'h	7390;
42156	:douta	=	16'h	6b4f;
42157	:douta	=	16'h	634e;
42158	:douta	=	16'h	6b4e;
42159	:douta	=	16'h	6b2f;
42160	:douta	=	16'h	6b2f;
42161	:douta	=	16'h	5a6b;
42162	:douta	=	16'h	41e7;
42163	:douta	=	16'h	5248;
42164	:douta	=	16'h	6b0c;
42165	:douta	=	16'h	736d;
42166	:douta	=	16'h	bd31;
42167	:douta	=	16'h	d5d3;
42168	:douta	=	16'h	cd72;
42169	:douta	=	16'h	de35;
42170	:douta	=	16'h	de56;
42171	:douta	=	16'h	de55;
42172	:douta	=	16'h	e656;
42173	:douta	=	16'h	de35;
42174	:douta	=	16'h	e635;
42175	:douta	=	16'h	de35;
42176	:douta	=	16'h	d5d4;
42177	:douta	=	16'h	9c93;
42178	:douta	=	16'h	a4d3;
42179	:douta	=	16'h	e616;
42180	:douta	=	16'h	c574;
42181	:douta	=	16'h	bd54;
42182	:douta	=	16'h	b514;
42183	:douta	=	16'h	acd4;
42184	:douta	=	16'h	9494;
42185	:douta	=	16'h	8432;
42186	:douta	=	16'h	8c73;
42187	:douta	=	16'h	8c52;
42188	:douta	=	16'h	8c73;
42189	:douta	=	16'h	8c53;
42190	:douta	=	16'h	8432;
42191	:douta	=	16'h	7bf2;
42192	:douta	=	16'h	73d1;
42193	:douta	=	16'h	73b0;
42194	:douta	=	16'h	73b1;
42195	:douta	=	16'h	73d2;
42196	:douta	=	16'h	73f2;
42197	:douta	=	16'h	6bb1;
42198	:douta	=	16'h	6bb1;
42199	:douta	=	16'h	6bb1;
42200	:douta	=	16'h	6bb2;
42201	:douta	=	16'h	5acd;
42202	:douta	=	16'h	39a6;
42203	:douta	=	16'h	49e8;
42204	:douta	=	16'h	5228;
42205	:douta	=	16'h	632d;
42206	:douta	=	16'h	52ce;
42207	:douta	=	16'h	4aad;
42208	:douta	=	16'h	320b;
42209	:douta	=	16'h	7c12;
42210	:douta	=	16'h	31c9;
42211	:douta	=	16'h	1906;
42212	:douta	=	16'h	18e5;
42213	:douta	=	16'h	1905;
42214	:douta	=	16'h	2925;
42215	:douta	=	16'h	59e4;
42216	:douta	=	16'h	6a25;
42217	:douta	=	16'h	6a05;
42218	:douta	=	16'h	6a26;
42219	:douta	=	16'h	6205;
42220	:douta	=	16'h	6205;
42221	:douta	=	16'h	59e5;
42222	:douta	=	16'h	59e6;
42223	:douta	=	16'h	5a06;
42224	:douta	=	16'h	51a5;
42225	:douta	=	16'h	51c5;
42226	:douta	=	16'h	51c5;
42227	:douta	=	16'h	51a5;
42228	:douta	=	16'h	51c6;
42229	:douta	=	16'h	51c5;
42230	:douta	=	16'h	51a6;
42231	:douta	=	16'h	49a5;
42232	:douta	=	16'h	49a6;
42233	:douta	=	16'h	49a5;
42234	:douta	=	16'h	49a6;
42235	:douta	=	16'h	4186;
42236	:douta	=	16'h	41a6;
42237	:douta	=	16'h	4186;
42238	:douta	=	16'h	4166;
42239	:douta	=	16'h	3966;
42240	:douta	=	16'h	f6f9;
42241	:douta	=	16'h	eeb7;
42242	:douta	=	16'h	f6d8;
42243	:douta	=	16'h	ff7b;
42244	:douta	=	16'h	f718;
42245	:douta	=	16'h	f6d8;
42246	:douta	=	16'h	fef9;
42247	:douta	=	16'h	ff7b;
42248	:douta	=	16'h	d5b4;
42249	:douta	=	16'h	cdb5;
42250	:douta	=	16'h	b515;
42251	:douta	=	16'h	9453;
42252	:douta	=	16'h	a515;
42253	:douta	=	16'h	ad56;
42254	:douta	=	16'h	a4f5;
42255	:douta	=	16'h	b515;
42256	:douta	=	16'h	b535;
42257	:douta	=	16'h	a4f5;
42258	:douta	=	16'h	9cd5;
42259	:douta	=	16'h	8c95;
42260	:douta	=	16'h	7413;
42261	:douta	=	16'h	7414;
42262	:douta	=	16'h	7414;
42263	:douta	=	16'h	8475;
42264	:douta	=	16'h	7c55;
42265	:douta	=	16'h	8476;
42266	:douta	=	16'h	8476;
42267	:douta	=	16'h	8496;
42268	:douta	=	16'h	7c55;
42269	:douta	=	16'h	7c54;
42270	:douta	=	16'h	7c34;
42271	:douta	=	16'h	8cb7;
42272	:douta	=	16'h	8d18;
42273	:douta	=	16'h	0042;
42274	:douta	=	16'h	10e5;
42275	:douta	=	16'h	10e5;
42276	:douta	=	16'h	10c5;
42277	:douta	=	16'h	10e5;
42278	:douta	=	16'h	10e5;
42279	:douta	=	16'h	10c4;
42280	:douta	=	16'h	10c4;
42281	:douta	=	16'h	1106;
42282	:douta	=	16'h	1105;
42283	:douta	=	16'h	10e5;
42284	:douta	=	16'h	1905;
42285	:douta	=	16'h	10e6;
42286	:douta	=	16'h	10e5;
42287	:douta	=	16'h	10c4;
42288	:douta	=	16'h	10e4;
42289	:douta	=	16'h	10e5;
42290	:douta	=	16'h	10c5;
42291	:douta	=	16'h	18e4;
42292	:douta	=	16'h	18e5;
42293	:douta	=	16'h	2947;
42294	:douta	=	16'h	18a4;
42295	:douta	=	16'h	18e5;
42296	:douta	=	16'h	29c9;
42297	:douta	=	16'h	29ca;
42298	:douta	=	16'h	2a2c;
42299	:douta	=	16'h	2168;
42300	:douta	=	16'h	2146;
42301	:douta	=	16'h	3209;
42302	:douta	=	16'h	31c8;
42303	:douta	=	16'h	39c8;
42304	:douta	=	16'h	5228;
42305	:douta	=	16'h	4963;
42306	:douta	=	16'h	4942;
42307	:douta	=	16'h	4901;
42308	:douta	=	16'h	5162;
42309	:douta	=	16'h	5183;
42310	:douta	=	16'h	5183;
42311	:douta	=	16'h	59c4;
42312	:douta	=	16'h	61c4;
42313	:douta	=	16'h	69e4;
42314	:douta	=	16'h	7224;
42315	:douta	=	16'h	7224;
42316	:douta	=	16'h	6a24;
42317	:douta	=	16'h	7224;
42318	:douta	=	16'h	7224;
42319	:douta	=	16'h	7a44;
42320	:douta	=	16'h	7a44;
42321	:douta	=	16'h	7a44;
42322	:douta	=	16'h	8284;
42323	:douta	=	16'h	8aa4;
42324	:douta	=	16'h	8ae4;
42325	:douta	=	16'h	8ac4;
42326	:douta	=	16'h	92e4;
42327	:douta	=	16'h	92e4;
42328	:douta	=	16'h	9b05;
42329	:douta	=	16'h	9b05;
42330	:douta	=	16'h	a325;
42331	:douta	=	16'h	a344;
42332	:douta	=	16'h	a345;
42333	:douta	=	16'h	ab86;
42334	:douta	=	16'h	ab64;
42335	:douta	=	16'h	b385;
42336	:douta	=	16'h	b365;
42337	:douta	=	16'h	b385;
42338	:douta	=	16'h	b3a5;
42339	:douta	=	16'h	b3c5;
42340	:douta	=	16'h	b3c4;
42341	:douta	=	16'h	bbc5;
42342	:douta	=	16'h	bbc6;
42343	:douta	=	16'h	bbc6;
42344	:douta	=	16'h	bbe6;
42345	:douta	=	16'h	bbe5;
42346	:douta	=	16'h	c3e4;
42347	:douta	=	16'h	bbc3;
42348	:douta	=	16'h	bba3;
42349	:douta	=	16'h	bb83;
42350	:douta	=	16'h	bbc2;
42351	:douta	=	16'h	c3e3;
42352	:douta	=	16'h	c426;
42353	:douta	=	16'h	ccaa;
42354	:douta	=	16'h	cd0c;
42355	:douta	=	16'h	d590;
42356	:douta	=	16'h	e674;
42357	:douta	=	16'h	e6d7;
42358	:douta	=	16'h	f77a;
42359	:douta	=	16'h	f79b;
42360	:douta	=	16'h	f7bb;
42361	:douta	=	16'h	ef58;
42362	:douta	=	16'h	ef17;
42363	:douta	=	16'h	e672;
42364	:douta	=	16'h	de30;
42365	:douta	=	16'h	dd6d;
42366	:douta	=	16'h	d4e8;
42367	:douta	=	16'h	d4a7;
42368	:douta	=	16'h	cc44;
42369	:douta	=	16'h	c420;
42370	:douta	=	16'h	c400;
42371	:douta	=	16'h	cc22;
42372	:douta	=	16'h	cc24;
42373	:douta	=	16'h	cc45;
42374	:douta	=	16'h	d446;
42375	:douta	=	16'h	d466;
42376	:douta	=	16'h	d467;
42377	:douta	=	16'h	d487;
42378	:douta	=	16'h	cc66;
42379	:douta	=	16'h	d486;
42380	:douta	=	16'h	d466;
42381	:douta	=	16'h	d466;
42382	:douta	=	16'h	d466;
42383	:douta	=	16'h	d466;
42384	:douta	=	16'h	d486;
42385	:douta	=	16'h	d466;
42386	:douta	=	16'h	d466;
42387	:douta	=	16'h	d466;
42388	:douta	=	16'h	d466;
42389	:douta	=	16'h	d466;
42390	:douta	=	16'h	d467;
42391	:douta	=	16'h	d486;
42392	:douta	=	16'h	d487;
42393	:douta	=	16'h	d465;
42394	:douta	=	16'h	b46d;
42395	:douta	=	16'h	a492;
42396	:douta	=	16'h	a516;
42397	:douta	=	16'h	ad56;
42398	:douta	=	16'h	a516;
42399	:douta	=	16'h	a537;
42400	:douta	=	16'h	ad37;
42401	:douta	=	16'h	9cd6;
42402	:douta	=	16'h	a537;
42403	:douta	=	16'h	b577;
42404	:douta	=	16'h	8c74;
42405	:douta	=	16'h	73b1;
42406	:douta	=	16'h	8c33;
42407	:douta	=	16'h	7bb1;
42408	:douta	=	16'h	73b1;
42409	:douta	=	16'h	6b70;
42410	:douta	=	16'h	632e;
42411	:douta	=	16'h	7370;
42412	:douta	=	16'h	632e;
42413	:douta	=	16'h	5aac;
42414	:douta	=	16'h	526a;
42415	:douta	=	16'h	39a7;
42416	:douta	=	16'h	41c7;
42417	:douta	=	16'h	7bae;
42418	:douta	=	16'h	a4b0;
42419	:douta	=	16'h	9c4f;
42420	:douta	=	16'h	c572;
42421	:douta	=	16'h	d614;
42422	:douta	=	16'h	de15;
42423	:douta	=	16'h	de35;
42424	:douta	=	16'h	cd72;
42425	:douta	=	16'h	ee97;
42426	:douta	=	16'h	e656;
42427	:douta	=	16'h	de15;
42428	:douta	=	16'h	d5f5;
42429	:douta	=	16'h	d5f5;
42430	:douta	=	16'h	d5f5;
42431	:douta	=	16'h	cd94;
42432	:douta	=	16'h	bd34;
42433	:douta	=	16'h	9cd4;
42434	:douta	=	16'h	9cb4;
42435	:douta	=	16'h	8432;
42436	:douta	=	16'h	9cd4;
42437	:douta	=	16'h	a4d5;
42438	:douta	=	16'h	9c93;
42439	:douta	=	16'h	8c52;
42440	:douta	=	16'h	8433;
42441	:douta	=	16'h	8c53;
42442	:douta	=	16'h	7bd1;
42443	:douta	=	16'h	7bd1;
42444	:douta	=	16'h	7bd1;
42445	:douta	=	16'h	73b0;
42446	:douta	=	16'h	73b0;
42447	:douta	=	16'h	632e;
42448	:douta	=	16'h	632e;
42449	:douta	=	16'h	632e;
42450	:douta	=	16'h	632f;
42451	:douta	=	16'h	630e;
42452	:douta	=	16'h	6b4f;
42453	:douta	=	16'h	632e;
42454	:douta	=	16'h	5acb;
42455	:douta	=	16'h	28e4;
42456	:douta	=	16'h	20a2;
42457	:douta	=	16'h	62ca;
42458	:douta	=	16'h	734d;
42459	:douta	=	16'h	83ee;
42460	:douta	=	16'h	736e;
42461	:douta	=	16'h	630e;
42462	:douta	=	16'h	428d;
42463	:douta	=	16'h	52cf;
42464	:douta	=	16'h	5b30;
42465	:douta	=	16'h	3a4a;
42466	:douta	=	16'h	634f;
42467	:douta	=	16'h	29a9;
42468	:douta	=	16'h	29aa;
42469	:douta	=	16'h	29a9;
42470	:douta	=	16'h	1105;
42471	:douta	=	16'h	10e5;
42472	:douta	=	16'h	7245;
42473	:douta	=	16'h	6226;
42474	:douta	=	16'h	6205;
42475	:douta	=	16'h	6226;
42476	:douta	=	16'h	6206;
42477	:douta	=	16'h	59e5;
42478	:douta	=	16'h	59e5;
42479	:douta	=	16'h	59e6;
42480	:douta	=	16'h	59e6;
42481	:douta	=	16'h	51c6;
42482	:douta	=	16'h	51c5;
42483	:douta	=	16'h	51a5;
42484	:douta	=	16'h	49a5;
42485	:douta	=	16'h	51a6;
42486	:douta	=	16'h	49a6;
42487	:douta	=	16'h	49a6;
42488	:douta	=	16'h	49a6;
42489	:douta	=	16'h	49a6;
42490	:douta	=	16'h	4185;
42491	:douta	=	16'h	41a6;
42492	:douta	=	16'h	4186;
42493	:douta	=	16'h	4186;
42494	:douta	=	16'h	4166;
42495	:douta	=	16'h	3965;
42496	:douta	=	16'h	f6f8;
42497	:douta	=	16'h	eeb7;
42498	:douta	=	16'h	f6f9;
42499	:douta	=	16'h	ff5b;
42500	:douta	=	16'h	ff3a;
42501	:douta	=	16'h	f6f8;
42502	:douta	=	16'h	f6f8;
42503	:douta	=	16'h	ff5a;
42504	:douta	=	16'h	cd73;
42505	:douta	=	16'h	c5b6;
42506	:douta	=	16'h	acf5;
42507	:douta	=	16'h	9473;
42508	:douta	=	16'h	ad36;
42509	:douta	=	16'h	b556;
42510	:douta	=	16'h	a4f5;
42511	:douta	=	16'h	b556;
42512	:douta	=	16'h	b535;
42513	:douta	=	16'h	ad15;
42514	:douta	=	16'h	9cd6;
42515	:douta	=	16'h	8474;
42516	:douta	=	16'h	7413;
42517	:douta	=	16'h	7414;
42518	:douta	=	16'h	7c55;
42519	:douta	=	16'h	7c35;
42520	:douta	=	16'h	7c55;
42521	:douta	=	16'h	7c55;
42522	:douta	=	16'h	8496;
42523	:douta	=	16'h	8496;
42524	:douta	=	16'h	7c54;
42525	:douta	=	16'h	7c14;
42526	:douta	=	16'h	7c34;
42527	:douta	=	16'h	9518;
42528	:douta	=	16'h	4b0f;
42529	:douta	=	16'h	10a4;
42530	:douta	=	16'h	10e5;
42531	:douta	=	16'h	1906;
42532	:douta	=	16'h	10a5;
42533	:douta	=	16'h	08a5;
42534	:douta	=	16'h	08e5;
42535	:douta	=	16'h	10e6;
42536	:douta	=	16'h	10e6;
42537	:douta	=	16'h	10e5;
42538	:douta	=	16'h	10e5;
42539	:douta	=	16'h	08a4;
42540	:douta	=	16'h	10e5;
42541	:douta	=	16'h	10e5;
42542	:douta	=	16'h	10e5;
42543	:douta	=	16'h	10c4;
42544	:douta	=	16'h	10c4;
42545	:douta	=	16'h	18e5;
42546	:douta	=	16'h	2127;
42547	:douta	=	16'h	1906;
42548	:douta	=	16'h	2126;
42549	:douta	=	16'h	2987;
42550	:douta	=	16'h	10a3;
42551	:douta	=	16'h	29ca;
42552	:douta	=	16'h	320a;
42553	:douta	=	16'h	3a4c;
42554	:douta	=	16'h	3166;
42555	:douta	=	16'h	30e3;
42556	:douta	=	16'h	3103;
42557	:douta	=	16'h	4123;
42558	:douta	=	16'h	4143;
42559	:douta	=	16'h	28c2;
42560	:douta	=	16'h	4100;
42561	:douta	=	16'h	4942;
42562	:douta	=	16'h	4964;
42563	:douta	=	16'h	4984;
42564	:douta	=	16'h	51a4;
42565	:douta	=	16'h	59c4;
42566	:douta	=	16'h	61e4;
42567	:douta	=	16'h	6a04;
42568	:douta	=	16'h	6a24;
42569	:douta	=	16'h	6a24;
42570	:douta	=	16'h	6a24;
42571	:douta	=	16'h	6a04;
42572	:douta	=	16'h	7204;
42573	:douta	=	16'h	7224;
42574	:douta	=	16'h	7244;
42575	:douta	=	16'h	7a44;
42576	:douta	=	16'h	7a44;
42577	:douta	=	16'h	8264;
42578	:douta	=	16'h	82a4;
42579	:douta	=	16'h	8aa4;
42580	:douta	=	16'h	8ac5;
42581	:douta	=	16'h	8ac4;
42582	:douta	=	16'h	92e4;
42583	:douta	=	16'h	9305;
42584	:douta	=	16'h	9b05;
42585	:douta	=	16'h	9b25;
42586	:douta	=	16'h	9b25;
42587	:douta	=	16'h	a344;
42588	:douta	=	16'h	a345;
42589	:douta	=	16'h	ab65;
42590	:douta	=	16'h	ab65;
42591	:douta	=	16'h	b385;
42592	:douta	=	16'h	b385;
42593	:douta	=	16'h	b3a5;
42594	:douta	=	16'h	b3c4;
42595	:douta	=	16'h	bbc4;
42596	:douta	=	16'h	b3c4;
42597	:douta	=	16'h	b3a4;
42598	:douta	=	16'h	b3a4;
42599	:douta	=	16'h	bb83;
42600	:douta	=	16'h	b363;
42601	:douta	=	16'h	b363;
42602	:douta	=	16'h	bbe4;
42603	:douta	=	16'h	c405;
42604	:douta	=	16'h	c489;
42605	:douta	=	16'h	ccca;
42606	:douta	=	16'h	d590;
42607	:douta	=	16'h	e654;
42608	:douta	=	16'h	eeb6;
42609	:douta	=	16'h	f759;
42610	:douta	=	16'h	f79b;
42611	:douta	=	16'h	f79a;
42612	:douta	=	16'h	ef59;
42613	:douta	=	16'h	ef17;
42614	:douta	=	16'h	e673;
42615	:douta	=	16'h	de31;
42616	:douta	=	16'h	dd8d;
42617	:douta	=	16'h	ccc9;
42618	:douta	=	16'h	d487;
42619	:douta	=	16'h	cc24;
42620	:douta	=	16'h	cbe3;
42621	:douta	=	16'h	cbe3;
42622	:douta	=	16'h	cc04;
42623	:douta	=	16'h	cc25;
42624	:douta	=	16'h	cc25;
42625	:douta	=	16'h	d446;
42626	:douta	=	16'h	cc46;
42627	:douta	=	16'h	d446;
42628	:douta	=	16'h	d466;
42629	:douta	=	16'h	cc66;
42630	:douta	=	16'h	d467;
42631	:douta	=	16'h	cc66;
42632	:douta	=	16'h	d467;
42633	:douta	=	16'h	d467;
42634	:douta	=	16'h	d467;
42635	:douta	=	16'h	d466;
42636	:douta	=	16'h	cc66;
42637	:douta	=	16'h	d487;
42638	:douta	=	16'h	cc66;
42639	:douta	=	16'h	d466;
42640	:douta	=	16'h	d466;
42641	:douta	=	16'h	d466;
42642	:douta	=	16'h	d467;
42643	:douta	=	16'h	d466;
42644	:douta	=	16'h	d466;
42645	:douta	=	16'h	d486;
42646	:douta	=	16'h	d467;
42647	:douta	=	16'h	cc66;
42648	:douta	=	16'h	d467;
42649	:douta	=	16'h	d485;
42650	:douta	=	16'h	cc66;
42651	:douta	=	16'h	9c52;
42652	:douta	=	16'h	a4f5;
42653	:douta	=	16'h	a536;
42654	:douta	=	16'h	9cd5;
42655	:douta	=	16'h	9cd5;
42656	:douta	=	16'h	9cb5;
42657	:douta	=	16'h	9494;
42658	:douta	=	16'h	9cd5;
42659	:douta	=	16'h	9cd4;
42660	:douta	=	16'h	8432;
42661	:douta	=	16'h	736f;
42662	:douta	=	16'h	9494;
42663	:douta	=	16'h	8432;
42664	:douta	=	16'h	7390;
42665	:douta	=	16'h	7390;
42666	:douta	=	16'h	6b2f;
42667	:douta	=	16'h	6b2f;
42668	:douta	=	16'h	630e;
42669	:douta	=	16'h	5a6a;
42670	:douta	=	16'h	49e7;
42671	:douta	=	16'h	6b0c;
42672	:douta	=	16'h	7b8d;
42673	:douta	=	16'h	c593;
42674	:douta	=	16'h	b511;
42675	:douta	=	16'h	acd1;
42676	:douta	=	16'h	de15;
42677	:douta	=	16'h	de56;
42678	:douta	=	16'h	de55;
42679	:douta	=	16'h	de35;
42680	:douta	=	16'h	cd92;
42681	:douta	=	16'h	e697;
42682	:douta	=	16'h	de56;
42683	:douta	=	16'h	d5d5;
42684	:douta	=	16'h	d5f5;
42685	:douta	=	16'h	cdb5;
42686	:douta	=	16'h	bd55;
42687	:douta	=	16'h	ad14;
42688	:douta	=	16'h	acf5;
42689	:douta	=	16'h	9cf5;
42690	:douta	=	16'h	8c73;
42691	:douta	=	16'h	8412;
42692	:douta	=	16'h	8433;
42693	:douta	=	16'h	94b5;
42694	:douta	=	16'h	8c73;
42695	:douta	=	16'h	8412;
42696	:douta	=	16'h	7bd1;
42697	:douta	=	16'h	7bd1;
42698	:douta	=	16'h	6b90;
42699	:douta	=	16'h	7bf1;
42700	:douta	=	16'h	73b0;
42701	:douta	=	16'h	6b4f;
42702	:douta	=	16'h	632e;
42703	:douta	=	16'h	632e;
42704	:douta	=	16'h	632f;
42705	:douta	=	16'h	632e;
42706	:douta	=	16'h	62cd;
42707	:douta	=	16'h	5acd;
42708	:douta	=	16'h	49e8;
42709	:douta	=	16'h	49c5;
42710	:douta	=	16'h	62a8;
42711	:douta	=	16'h	6b0b;
42712	:douta	=	16'h	732b;
42713	:douta	=	16'h	8bed;
42714	:douta	=	16'h	acb0;
42715	:douta	=	16'h	b4f0;
42716	:douta	=	16'h	62ed;
42717	:douta	=	16'h	4a6c;
42718	:douta	=	16'h	3a2b;
42719	:douta	=	16'h	422a;
42720	:douta	=	16'h	422b;
42721	:douta	=	16'h	2147;
42722	:douta	=	16'h	52ae;
42723	:douta	=	16'h	29ca;
42724	:douta	=	16'h	29c9;
42725	:douta	=	16'h	29ca;
42726	:douta	=	16'h	2147;
42727	:douta	=	16'h	08a4;
42728	:douta	=	16'h	7245;
42729	:douta	=	16'h	6a46;
42730	:douta	=	16'h	6a26;
42731	:douta	=	16'h	6226;
42732	:douta	=	16'h	6206;
42733	:douta	=	16'h	59e5;
42734	:douta	=	16'h	59c5;
42735	:douta	=	16'h	59e6;
42736	:douta	=	16'h	59c6;
42737	:douta	=	16'h	51c6;
42738	:douta	=	16'h	51c5;
42739	:douta	=	16'h	49a5;
42740	:douta	=	16'h	51c5;
42741	:douta	=	16'h	49a6;
42742	:douta	=	16'h	51a6;
42743	:douta	=	16'h	4986;
42744	:douta	=	16'h	49a6;
42745	:douta	=	16'h	49a5;
42746	:douta	=	16'h	4185;
42747	:douta	=	16'h	41a6;
42748	:douta	=	16'h	4186;
42749	:douta	=	16'h	4166;
42750	:douta	=	16'h	4186;
42751	:douta	=	16'h	3966;
42752	:douta	=	16'h	f6f9;
42753	:douta	=	16'h	ff19;
42754	:douta	=	16'h	ff5b;
42755	:douta	=	16'h	ff7b;
42756	:douta	=	16'h	ff7b;
42757	:douta	=	16'h	ff5a;
42758	:douta	=	16'h	ff5a;
42759	:douta	=	16'h	eeb9;
42760	:douta	=	16'h	ddf5;
42761	:douta	=	16'h	acf5;
42762	:douta	=	16'h	acf5;
42763	:douta	=	16'h	a4d5;
42764	:douta	=	16'h	b577;
42765	:douta	=	16'h	ad36;
42766	:douta	=	16'h	b555;
42767	:douta	=	16'h	b514;
42768	:douta	=	16'h	b535;
42769	:douta	=	16'h	ad16;
42770	:douta	=	16'h	9cd6;
42771	:douta	=	16'h	73f3;
42772	:douta	=	16'h	7413;
42773	:douta	=	16'h	7c34;
42774	:douta	=	16'h	7c55;
42775	:douta	=	16'h	7c55;
42776	:douta	=	16'h	7c55;
42777	:douta	=	16'h	8476;
42778	:douta	=	16'h	8cb6;
42779	:douta	=	16'h	8476;
42780	:douta	=	16'h	7413;
42781	:douta	=	16'h	7c54;
42782	:douta	=	16'h	8496;
42783	:douta	=	16'h	322a;
42784	:douta	=	16'h	0001;
42785	:douta	=	16'h	10c4;
42786	:douta	=	16'h	0863;
42787	:douta	=	16'h	0883;
42788	:douta	=	16'h	08a4;
42789	:douta	=	16'h	08a4;
42790	:douta	=	16'h	10a4;
42791	:douta	=	16'h	10a5;
42792	:douta	=	16'h	10e5;
42793	:douta	=	16'h	1967;
42794	:douta	=	16'h	2168;
42795	:douta	=	16'h	2188;
42796	:douta	=	16'h	2168;
42797	:douta	=	16'h	29ca;
42798	:douta	=	16'h	29ca;
42799	:douta	=	16'h	29ca;
42800	:douta	=	16'h	29cb;
42801	:douta	=	16'h	29c9;
42802	:douta	=	16'h	2105;
42803	:douta	=	16'h	20e4;
42804	:douta	=	16'h	2126;
42805	:douta	=	16'h	2967;
42806	:douta	=	16'h	18c4;
42807	:douta	=	16'h	28a1;
42808	:douta	=	16'h	30e2;
42809	:douta	=	16'h	30c2;
42810	:douta	=	16'h	3902;
42811	:douta	=	16'h	4143;
42812	:douta	=	16'h	4143;
42813	:douta	=	16'h	4963;
42814	:douta	=	16'h	5184;
42815	:douta	=	16'h	3102;
42816	:douta	=	16'h	59c4;
42817	:douta	=	16'h	59c4;
42818	:douta	=	16'h	61c4;
42819	:douta	=	16'h	59c4;
42820	:douta	=	16'h	59e3;
42821	:douta	=	16'h	6203;
42822	:douta	=	16'h	6204;
42823	:douta	=	16'h	61e4;
42824	:douta	=	16'h	6a04;
42825	:douta	=	16'h	7224;
42826	:douta	=	16'h	6a24;
42827	:douta	=	16'h	7224;
42828	:douta	=	16'h	7224;
42829	:douta	=	16'h	7224;
42830	:douta	=	16'h	7a44;
42831	:douta	=	16'h	7a64;
42832	:douta	=	16'h	7a64;
42833	:douta	=	16'h	8284;
42834	:douta	=	16'h	8284;
42835	:douta	=	16'h	8aa4;
42836	:douta	=	16'h	8ac4;
42837	:douta	=	16'h	8ae4;
42838	:douta	=	16'h	9304;
42839	:douta	=	16'h	9b05;
42840	:douta	=	16'h	9b05;
42841	:douta	=	16'h	9b25;
42842	:douta	=	16'h	9b25;
42843	:douta	=	16'h	a345;
42844	:douta	=	16'h	a324;
42845	:douta	=	16'h	a303;
42846	:douta	=	16'h	a323;
42847	:douta	=	16'h	ab22;
42848	:douta	=	16'h	ab43;
42849	:douta	=	16'h	ab65;
42850	:douta	=	16'h	bc07;
42851	:douta	=	16'h	bc48;
42852	:douta	=	16'h	cd2e;
42853	:douta	=	16'h	de13;
42854	:douta	=	16'h	e675;
42855	:douta	=	16'h	ef18;
42856	:douta	=	16'h	ef59;
42857	:douta	=	16'h	f79a;
42858	:douta	=	16'h	ef58;
42859	:douta	=	16'h	ef17;
42860	:douta	=	16'h	e672;
42861	:douta	=	16'h	de31;
42862	:douta	=	16'h	d56d;
42863	:douta	=	16'h	cce9;
42864	:douta	=	16'h	cc87;
42865	:douta	=	16'h	c403;
42866	:douta	=	16'h	c3e2;
42867	:douta	=	16'h	c3e2;
42868	:douta	=	16'h	c3e2;
42869	:douta	=	16'h	c404;
42870	:douta	=	16'h	cc05;
42871	:douta	=	16'h	cc25;
42872	:douta	=	16'h	cc45;
42873	:douta	=	16'h	cc46;
42874	:douta	=	16'h	cc47;
42875	:douta	=	16'h	cc66;
42876	:douta	=	16'h	cc45;
42877	:douta	=	16'h	cc46;
42878	:douta	=	16'h	cc46;
42879	:douta	=	16'h	cc45;
42880	:douta	=	16'h	cc46;
42881	:douta	=	16'h	cc65;
42882	:douta	=	16'h	cc66;
42883	:douta	=	16'h	cc66;
42884	:douta	=	16'h	cc66;
42885	:douta	=	16'h	d466;
42886	:douta	=	16'h	cc46;
42887	:douta	=	16'h	d466;
42888	:douta	=	16'h	d466;
42889	:douta	=	16'h	d466;
42890	:douta	=	16'h	d467;
42891	:douta	=	16'h	d466;
42892	:douta	=	16'h	d466;
42893	:douta	=	16'h	d466;
42894	:douta	=	16'h	d487;
42895	:douta	=	16'h	d466;
42896	:douta	=	16'h	d466;
42897	:douta	=	16'h	d466;
42898	:douta	=	16'h	d467;
42899	:douta	=	16'h	d467;
42900	:douta	=	16'h	d466;
42901	:douta	=	16'h	d466;
42902	:douta	=	16'h	d467;
42903	:douta	=	16'h	d467;
42904	:douta	=	16'h	cc86;
42905	:douta	=	16'h	d466;
42906	:douta	=	16'h	d486;
42907	:douta	=	16'h	d465;
42908	:douta	=	16'h	8c10;
42909	:douta	=	16'h	9451;
42910	:douta	=	16'h	9cd4;
42911	:douta	=	16'h	9453;
42912	:douta	=	16'h	8c11;
42913	:douta	=	16'h	9473;
42914	:douta	=	16'h	9453;
42915	:douta	=	16'h	83f1;
42916	:douta	=	16'h	8412;
42917	:douta	=	16'h	7bd1;
42918	:douta	=	16'h	7bd1;
42919	:douta	=	16'h	7391;
42920	:douta	=	16'h	7390;
42921	:douta	=	16'h	630e;
42922	:douta	=	16'h	41c8;
42923	:douta	=	16'h	49e7;
42924	:douta	=	16'h	acd0;
42925	:douta	=	16'h	7b4b;
42926	:douta	=	16'h	a46e;
42927	:douta	=	16'h	c592;
42928	:douta	=	16'h	d5f4;
42929	:douta	=	16'h	de55;
42930	:douta	=	16'h	b532;
42931	:douta	=	16'h	e6b7;
42932	:douta	=	16'h	e656;
42933	:douta	=	16'h	e696;
42934	:douta	=	16'h	de55;
42935	:douta	=	16'h	e656;
42936	:douta	=	16'h	cdb4;
42937	:douta	=	16'h	d616;
42938	:douta	=	16'h	d5f6;
42939	:douta	=	16'h	cd95;
42940	:douta	=	16'h	bd75;
42941	:douta	=	16'h	b555;
42942	:douta	=	16'h	a4f6;
42943	:douta	=	16'h	9cd5;
42944	:douta	=	16'h	8c74;
42945	:douta	=	16'h	9474;
42946	:douta	=	16'h	94b4;
42947	:douta	=	16'h	8c53;
42948	:douta	=	16'h	8c74;
42949	:douta	=	16'h	8433;
42950	:douta	=	16'h	8452;
42951	:douta	=	16'h	7bf1;
42952	:douta	=	16'h	73d1;
42953	:douta	=	16'h	6b4f;
42954	:douta	=	16'h	6b4f;
42955	:douta	=	16'h	8411;
42956	:douta	=	16'h	6b6f;
42957	:douta	=	16'h	6b2e;
42958	:douta	=	16'h	630d;
42959	:douta	=	16'h	630c;
42960	:douta	=	16'h	5229;
42961	:douta	=	16'h	5a48;
42962	:douta	=	16'h	93ed;
42963	:douta	=	16'h	940d;
42964	:douta	=	16'h	940e;
42965	:douta	=	16'h	8bcd;
42966	:douta	=	16'h	8bcd;
42967	:douta	=	16'h	a46e;
42968	:douta	=	16'h	a48f;
42969	:douta	=	16'h	acb0;
42970	:douta	=	16'h	b4f1;
42971	:douta	=	16'h	b4d1;
42972	:douta	=	16'h	5acd;
42973	:douta	=	16'h	3a2a;
42974	:douta	=	16'h	4209;
42975	:douta	=	16'h	31a8;
42976	:douta	=	16'h	3188;
42977	:douta	=	16'h	2948;
42978	:douta	=	16'h	31ea;
42979	:douta	=	16'h	10e6;
42980	:douta	=	16'h	10e4;
42981	:douta	=	16'h	10c5;
42982	:douta	=	16'h	18e5;
42983	:douta	=	16'h	18e5;
42984	:douta	=	16'h	3966;
42985	:douta	=	16'h	6206;
42986	:douta	=	16'h	6206;
42987	:douta	=	16'h	6205;
42988	:douta	=	16'h	59e5;
42989	:douta	=	16'h	59e5;
42990	:douta	=	16'h	59e6;
42991	:douta	=	16'h	59e6;
42992	:douta	=	16'h	51c5;
42993	:douta	=	16'h	51c5;
42994	:douta	=	16'h	51a5;
42995	:douta	=	16'h	49a5;
42996	:douta	=	16'h	49a5;
42997	:douta	=	16'h	49a6;
42998	:douta	=	16'h	49a6;
42999	:douta	=	16'h	49a6;
43000	:douta	=	16'h	4165;
43001	:douta	=	16'h	4185;
43002	:douta	=	16'h	41a6;
43003	:douta	=	16'h	4185;
43004	:douta	=	16'h	4186;
43005	:douta	=	16'h	4186;
43006	:douta	=	16'h	4166;
43007	:douta	=	16'h	4166;
43008	:douta	=	16'h	f6d8;
43009	:douta	=	16'h	f73a;
43010	:douta	=	16'h	ff7b;
43011	:douta	=	16'h	ff9c;
43012	:douta	=	16'h	ffbd;
43013	:douta	=	16'h	ffbd;
43014	:douta	=	16'h	ff3a;
43015	:douta	=	16'h	de57;
43016	:douta	=	16'h	de16;
43017	:douta	=	16'h	a4f5;
43018	:douta	=	16'h	9c94;
43019	:douta	=	16'h	b536;
43020	:douta	=	16'h	b577;
43021	:douta	=	16'h	ad15;
43022	:douta	=	16'h	bd75;
43023	:douta	=	16'h	b535;
43024	:douta	=	16'h	ad15;
43025	:douta	=	16'h	acf5;
43026	:douta	=	16'h	9cb5;
43027	:douta	=	16'h	73f3;
43028	:douta	=	16'h	7c34;
43029	:douta	=	16'h	7c35;
43030	:douta	=	16'h	7c54;
43031	:douta	=	16'h	8475;
43032	:douta	=	16'h	8496;
43033	:douta	=	16'h	8cb7;
43034	:douta	=	16'h	8496;
43035	:douta	=	16'h	7c75;
43036	:douta	=	16'h	7c33;
43037	:douta	=	16'h	7c74;
43038	:douta	=	16'h	94f7;
43039	:douta	=	16'h	0084;
43040	:douta	=	16'h	1063;
43041	:douta	=	16'h	10e5;
43042	:douta	=	16'h	1967;
43043	:douta	=	16'h	10e5;
43044	:douta	=	16'h	10e5;
43045	:douta	=	16'h	10e5;
43046	:douta	=	16'h	10e6;
43047	:douta	=	16'h	1928;
43048	:douta	=	16'h	29ca;
43049	:douta	=	16'h	2a0c;
43050	:douta	=	16'h	220c;
43051	:douta	=	16'h	21aa;
43052	:douta	=	16'h	21ca;
43053	:douta	=	16'h	29eb;
43054	:douta	=	16'h	2167;
43055	:douta	=	16'h	2105;
43056	:douta	=	16'h	20e4;
43057	:douta	=	16'h	20a2;
43058	:douta	=	16'h	2081;
43059	:douta	=	16'h	2081;
43060	:douta	=	16'h	20e3;
43061	:douta	=	16'h	2947;
43062	:douta	=	16'h	20c3;
43063	:douta	=	16'h	3103;
43064	:douta	=	16'h	3923;
43065	:douta	=	16'h	3923;
43066	:douta	=	16'h	4144;
43067	:douta	=	16'h	4163;
43068	:douta	=	16'h	4964;
43069	:douta	=	16'h	4964;
43070	:douta	=	16'h	4984;
43071	:douta	=	16'h	3923;
43072	:douta	=	16'h	61c4;
43073	:douta	=	16'h	59c4;
43074	:douta	=	16'h	59c4;
43075	:douta	=	16'h	61c4;
43076	:douta	=	16'h	59e4;
43077	:douta	=	16'h	61e4;
43078	:douta	=	16'h	61e4;
43079	:douta	=	16'h	61e4;
43080	:douta	=	16'h	6a04;
43081	:douta	=	16'h	7224;
43082	:douta	=	16'h	7204;
43083	:douta	=	16'h	7224;
43084	:douta	=	16'h	7224;
43085	:douta	=	16'h	7224;
43086	:douta	=	16'h	7a44;
43087	:douta	=	16'h	7a64;
43088	:douta	=	16'h	7a64;
43089	:douta	=	16'h	8264;
43090	:douta	=	16'h	82a4;
43091	:douta	=	16'h	8aa4;
43092	:douta	=	16'h	8ac4;
43093	:douta	=	16'h	92c4;
43094	:douta	=	16'h	92c4;
43095	:douta	=	16'h	92c4;
43096	:douta	=	16'h	92c4;
43097	:douta	=	16'h	92c3;
43098	:douta	=	16'h	92a2;
43099	:douta	=	16'h	9ae3;
43100	:douta	=	16'h	a324;
43101	:douta	=	16'h	abc7;
43102	:douta	=	16'h	b408;
43103	:douta	=	16'h	bcac;
43104	:douta	=	16'h	d5d1;
43105	:douta	=	16'h	de33;
43106	:douta	=	16'h	e6d6;
43107	:douta	=	16'h	ef18;
43108	:douta	=	16'h	f77a;
43109	:douta	=	16'h	ef58;
43110	:douta	=	16'h	ef16;
43111	:douta	=	16'h	e652;
43112	:douta	=	16'h	de11;
43113	:douta	=	16'h	d56e;
43114	:douta	=	16'h	cce9;
43115	:douta	=	16'h	c486;
43116	:douta	=	16'h	c423;
43117	:douta	=	16'h	c3e3;
43118	:douta	=	16'h	c3a3;
43119	:douta	=	16'h	c3c3;
43120	:douta	=	16'h	c3c3;
43121	:douta	=	16'h	c405;
43122	:douta	=	16'h	c405;
43123	:douta	=	16'h	cc26;
43124	:douta	=	16'h	cc25;
43125	:douta	=	16'h	cc46;
43126	:douta	=	16'h	c445;
43127	:douta	=	16'h	cc45;
43128	:douta	=	16'h	cc45;
43129	:douta	=	16'h	cc45;
43130	:douta	=	16'h	cc45;
43131	:douta	=	16'h	cc45;
43132	:douta	=	16'h	d466;
43133	:douta	=	16'h	cc46;
43134	:douta	=	16'h	cc46;
43135	:douta	=	16'h	cc46;
43136	:douta	=	16'h	d446;
43137	:douta	=	16'h	cc46;
43138	:douta	=	16'h	cc46;
43139	:douta	=	16'h	d466;
43140	:douta	=	16'h	cc66;
43141	:douta	=	16'h	d466;
43142	:douta	=	16'h	cc66;
43143	:douta	=	16'h	d466;
43144	:douta	=	16'h	d467;
43145	:douta	=	16'h	d467;
43146	:douta	=	16'h	d466;
43147	:douta	=	16'h	cc66;
43148	:douta	=	16'h	d466;
43149	:douta	=	16'h	d466;
43150	:douta	=	16'h	cc66;
43151	:douta	=	16'h	d466;
43152	:douta	=	16'h	d466;
43153	:douta	=	16'h	d466;
43154	:douta	=	16'h	d467;
43155	:douta	=	16'h	d466;
43156	:douta	=	16'h	d466;
43157	:douta	=	16'h	d467;
43158	:douta	=	16'h	d487;
43159	:douta	=	16'h	d467;
43160	:douta	=	16'h	d485;
43161	:douta	=	16'h	d466;
43162	:douta	=	16'h	d466;
43163	:douta	=	16'h	dc65;
43164	:douta	=	16'h	b44c;
43165	:douta	=	16'h	8c31;
43166	:douta	=	16'h	9473;
43167	:douta	=	16'h	9c93;
43168	:douta	=	16'h	8bf2;
43169	:douta	=	16'h	83d0;
43170	:douta	=	16'h	83d1;
43171	:douta	=	16'h	7bb0;
43172	:douta	=	16'h	83d1;
43173	:douta	=	16'h	7bf2;
43174	:douta	=	16'h	73b1;
43175	:douta	=	16'h	6b6f;
43176	:douta	=	16'h	5269;
43177	:douta	=	16'h	5248;
43178	:douta	=	16'h	5a49;
43179	:douta	=	16'h	acf1;
43180	:douta	=	16'h	836c;
43181	:douta	=	16'h	bd52;
43182	:douta	=	16'h	c5b2;
43183	:douta	=	16'h	d614;
43184	:douta	=	16'h	de35;
43185	:douta	=	16'h	cdd5;
43186	:douta	=	16'h	b512;
43187	:douta	=	16'h	e696;
43188	:douta	=	16'h	e656;
43189	:douta	=	16'h	e676;
43190	:douta	=	16'h	de35;
43191	:douta	=	16'h	e675;
43192	:douta	=	16'h	d5f4;
43193	:douta	=	16'h	c595;
43194	:douta	=	16'h	c595;
43195	:douta	=	16'h	bd54;
43196	:douta	=	16'h	b515;
43197	:douta	=	16'h	acf5;
43198	:douta	=	16'h	9cb5;
43199	:douta	=	16'h	9cd5;
43200	:douta	=	16'h	8c74;
43201	:douta	=	16'h	8412;
43202	:douta	=	16'h	8412;
43203	:douta	=	16'h	8453;
43204	:douta	=	16'h	8c73;
43205	:douta	=	16'h	8c53;
43206	:douta	=	16'h	8432;
43207	:douta	=	16'h	73d1;
43208	:douta	=	16'h	7390;
43209	:douta	=	16'h	6b4f;
43210	:douta	=	16'h	632f;
43211	:douta	=	16'h	8c32;
43212	:douta	=	16'h	8c12;
43213	:douta	=	16'h	524a;
43214	:douta	=	16'h	4a28;
43215	:douta	=	16'h	3103;
43216	:douta	=	16'h	41a5;
43217	:douta	=	16'h	41c5;
43218	:douta	=	16'h	93ec;
43219	:douta	=	16'h	b4ef;
43220	:douta	=	16'h	c572;
43221	:douta	=	16'h	b531;
43222	:douta	=	16'h	a4b0;
43223	:douta	=	16'h	a46f;
43224	:douta	=	16'h	a48f;
43225	:douta	=	16'h	acd0;
43226	:douta	=	16'h	b4d1;
43227	:douta	=	16'h	acd1;
43228	:douta	=	16'h	630d;
43229	:douta	=	16'h	422b;
43230	:douta	=	16'h	3a09;
43231	:douta	=	16'h	39e8;
43232	:douta	=	16'h	31a9;
43233	:douta	=	16'h	2147;
43234	:douta	=	16'h	1906;
43235	:douta	=	16'h	18e4;
43236	:douta	=	16'h	18e5;
43237	:douta	=	16'h	10e4;
43238	:douta	=	16'h	1926;
43239	:douta	=	16'h	1926;
43240	:douta	=	16'h	18e5;
43241	:douta	=	16'h	7246;
43242	:douta	=	16'h	6226;
43243	:douta	=	16'h	59e5;
43244	:douta	=	16'h	6206;
43245	:douta	=	16'h	6206;
43246	:douta	=	16'h	59c5;
43247	:douta	=	16'h	59e6;
43248	:douta	=	16'h	51c6;
43249	:douta	=	16'h	51c5;
43250	:douta	=	16'h	51a5;
43251	:douta	=	16'h	49a5;
43252	:douta	=	16'h	49a5;
43253	:douta	=	16'h	49a6;
43254	:douta	=	16'h	49a6;
43255	:douta	=	16'h	4986;
43256	:douta	=	16'h	4186;
43257	:douta	=	16'h	4185;
43258	:douta	=	16'h	41a6;
43259	:douta	=	16'h	41a6;
43260	:douta	=	16'h	4186;
43261	:douta	=	16'h	3965;
43262	:douta	=	16'h	4186;
43263	:douta	=	16'h	4166;
43264	:douta	=	16'h	f719;
43265	:douta	=	16'h	ff7b;
43266	:douta	=	16'h	ffbc;
43267	:douta	=	16'h	ffbd;
43268	:douta	=	16'h	ffbc;
43269	:douta	=	16'h	ffdd;
43270	:douta	=	16'h	de56;
43271	:douta	=	16'h	e657;
43272	:douta	=	16'h	d5f6;
43273	:douta	=	16'h	a4b4;
43274	:douta	=	16'h	9473;
43275	:douta	=	16'h	b556;
43276	:douta	=	16'h	b576;
43277	:douta	=	16'h	b535;
43278	:douta	=	16'h	bd75;
43279	:douta	=	16'h	bd76;
43280	:douta	=	16'h	ad36;
43281	:douta	=	16'h	a4f5;
43282	:douta	=	16'h	8c75;
43283	:douta	=	16'h	7413;
43284	:douta	=	16'h	7c54;
43285	:douta	=	16'h	8455;
43286	:douta	=	16'h	8475;
43287	:douta	=	16'h	8475;
43288	:douta	=	16'h	8476;
43289	:douta	=	16'h	8475;
43290	:douta	=	16'h	7c75;
43291	:douta	=	16'h	7c34;
43292	:douta	=	16'h	7c34;
43293	:douta	=	16'h	8c96;
43294	:douta	=	16'h	4aae;
43295	:douta	=	16'h	326e;
43296	:douta	=	16'h	2a4e;
43297	:douta	=	16'h	21cb;
43298	:douta	=	16'h	220d;
43299	:douta	=	16'h	2a2d;
43300	:douta	=	16'h	21ec;
43301	:douta	=	16'h	21cb;
43302	:douta	=	16'h	21a9;
43303	:douta	=	16'h	18a3;
43304	:douta	=	16'h	18a3;
43305	:douta	=	16'h	1881;
43306	:douta	=	16'h	1061;
43307	:douta	=	16'h	1861;
43308	:douta	=	16'h	1881;
43309	:douta	=	16'h	1881;
43310	:douta	=	16'h	20a2;
43311	:douta	=	16'h	20a2;
43312	:douta	=	16'h	20c2;
43313	:douta	=	16'h	28c2;
43314	:douta	=	16'h	28e3;
43315	:douta	=	16'h	2903;
43316	:douta	=	16'h	2925;
43317	:douta	=	16'h	2126;
43318	:douta	=	16'h	2904;
43319	:douta	=	16'h	4123;
43320	:douta	=	16'h	3923;
43321	:douta	=	16'h	3923;
43322	:douta	=	16'h	4143;
43323	:douta	=	16'h	4144;
43324	:douta	=	16'h	4984;
43325	:douta	=	16'h	4964;
43326	:douta	=	16'h	5184;
43327	:douta	=	16'h	51a4;
43328	:douta	=	16'h	4143;
43329	:douta	=	16'h	61c4;
43330	:douta	=	16'h	59c4;
43331	:douta	=	16'h	59c4;
43332	:douta	=	16'h	61e4;
43333	:douta	=	16'h	61e4;
43334	:douta	=	16'h	61e4;
43335	:douta	=	16'h	6a04;
43336	:douta	=	16'h	6a04;
43337	:douta	=	16'h	7224;
43338	:douta	=	16'h	7204;
43339	:douta	=	16'h	7204;
43340	:douta	=	16'h	7224;
43341	:douta	=	16'h	7224;
43342	:douta	=	16'h	7224;
43343	:douta	=	16'h	7203;
43344	:douta	=	16'h	7203;
43345	:douta	=	16'h	7223;
43346	:douta	=	16'h	8244;
43347	:douta	=	16'h	8ac6;
43348	:douta	=	16'h	9b89;
43349	:douta	=	16'h	a40a;
43350	:douta	=	16'h	bd2f;
43351	:douta	=	16'h	c591;
43352	:douta	=	16'h	d654;
43353	:douta	=	16'h	de95;
43354	:douta	=	16'h	e716;
43355	:douta	=	16'h	e6f6;
43356	:douta	=	16'h	e6b5;
43357	:douta	=	16'h	de32;
43358	:douta	=	16'h	d5f0;
43359	:douta	=	16'h	cd4e;
43360	:douta	=	16'h	bc89;
43361	:douta	=	16'h	bc27;
43362	:douta	=	16'h	bbe5;
43363	:douta	=	16'h	b3a2;
43364	:douta	=	16'h	b363;
43365	:douta	=	16'h	bb83;
43366	:douta	=	16'h	bbc3;
43367	:douta	=	16'h	bbc4;
43368	:douta	=	16'h	bbc5;
43369	:douta	=	16'h	c3e5;
43370	:douta	=	16'h	c406;
43371	:douta	=	16'h	c405;
43372	:douta	=	16'h	c405;
43373	:douta	=	16'h	c405;
43374	:douta	=	16'h	c405;
43375	:douta	=	16'h	c425;
43376	:douta	=	16'h	c405;
43377	:douta	=	16'h	cc25;
43378	:douta	=	16'h	cc25;
43379	:douta	=	16'h	cc26;
43380	:douta	=	16'h	cc26;
43381	:douta	=	16'h	cc26;
43382	:douta	=	16'h	cc46;
43383	:douta	=	16'h	cc46;
43384	:douta	=	16'h	cc46;
43385	:douta	=	16'h	cc45;
43386	:douta	=	16'h	cc45;
43387	:douta	=	16'h	cc45;
43388	:douta	=	16'h	cc45;
43389	:douta	=	16'h	cc45;
43390	:douta	=	16'h	cc47;
43391	:douta	=	16'h	d467;
43392	:douta	=	16'h	cc66;
43393	:douta	=	16'h	d466;
43394	:douta	=	16'h	cc66;
43395	:douta	=	16'h	cc46;
43396	:douta	=	16'h	cc66;
43397	:douta	=	16'h	cc66;
43398	:douta	=	16'h	cc66;
43399	:douta	=	16'h	d466;
43400	:douta	=	16'h	d466;
43401	:douta	=	16'h	cc66;
43402	:douta	=	16'h	d467;
43403	:douta	=	16'h	d466;
43404	:douta	=	16'h	d466;
43405	:douta	=	16'h	d466;
43406	:douta	=	16'h	d466;
43407	:douta	=	16'h	d466;
43408	:douta	=	16'h	d466;
43409	:douta	=	16'h	d466;
43410	:douta	=	16'h	d466;
43411	:douta	=	16'h	d466;
43412	:douta	=	16'h	d466;
43413	:douta	=	16'h	d466;
43414	:douta	=	16'h	d467;
43415	:douta	=	16'h	d466;
43416	:douta	=	16'h	d467;
43417	:douta	=	16'h	d467;
43418	:douta	=	16'h	d466;
43419	:douta	=	16'h	d488;
43420	:douta	=	16'h	cc86;
43421	:douta	=	16'h	dc84;
43422	:douta	=	16'h	bc8c;
43423	:douta	=	16'h	8c52;
43424	:douta	=	16'h	9452;
43425	:douta	=	16'h	8411;
43426	:douta	=	16'h	7bb1;
43427	:douta	=	16'h	7b90;
43428	:douta	=	16'h	736f;
43429	:douta	=	16'h	5a69;
43430	:douta	=	16'h	5a89;
43431	:douta	=	16'h	734b;
43432	:douta	=	16'h	944e;
43433	:douta	=	16'h	940d;
43434	:douta	=	16'h	f6f7;
43435	:douta	=	16'h	c552;
43436	:douta	=	16'h	d615;
43437	:douta	=	16'h	de35;
43438	:douta	=	16'h	de36;
43439	:douta	=	16'h	d635;
43440	:douta	=	16'h	de56;
43441	:douta	=	16'h	bd33;
43442	:douta	=	16'h	b513;
43443	:douta	=	16'h	cdd5;
43444	:douta	=	16'h	c595;
43445	:douta	=	16'h	c595;
43446	:douta	=	16'h	bd36;
43447	:douta	=	16'h	acf5;
43448	:douta	=	16'h	a4d4;
43449	:douta	=	16'h	a4f4;
43450	:douta	=	16'h	9cd4;
43451	:douta	=	16'h	94b4;
43452	:douta	=	16'h	8c53;
43453	:douta	=	16'h	7c12;
43454	:douta	=	16'h	8453;
43455	:douta	=	16'h	8c94;
43456	:douta	=	16'h	7c12;
43457	:douta	=	16'h	8c33;
43458	:douta	=	16'h	83f2;
43459	:douta	=	16'h	632f;
43460	:douta	=	16'h	73d1;
43461	:douta	=	16'h	8c32;
43462	:douta	=	16'h	8433;
43463	:douta	=	16'h	73f1;
43464	:douta	=	16'h	8412;
43465	:douta	=	16'h	6b4e;
43466	:douta	=	16'h	4a28;
43467	:douta	=	16'h	1060;
43468	:douta	=	16'h	18c1;
43469	:douta	=	16'h	7b2b;
43470	:douta	=	16'h	ac8f;
43471	:douta	=	16'h	bd53;
43472	:douta	=	16'h	9c50;
43473	:douta	=	16'h	8c0d;
43474	:douta	=	16'h	732a;
43475	:douta	=	16'h	5248;
43476	:douta	=	16'h	5269;
43477	:douta	=	16'h	ac8f;
43478	:douta	=	16'h	c552;
43479	:douta	=	16'h	d5d4;
43480	:douta	=	16'h	d5d4;
43481	:douta	=	16'h	c553;
43482	:douta	=	16'h	acf1;
43483	:douta	=	16'h	a470;
43484	:douta	=	16'h	734e;
43485	:douta	=	16'h	62ed;
43486	:douta	=	16'h	6b0c;
43487	:douta	=	16'h	31e9;
43488	:douta	=	16'h	2147;
43489	:douta	=	16'h	18e5;
43490	:douta	=	16'h	1905;
43491	:douta	=	16'h	420a;
43492	:douta	=	16'h	1926;
43493	:douta	=	16'h	29a9;
43494	:douta	=	16'h	29c9;
43495	:douta	=	16'h	29a8;
43496	:douta	=	16'h	1906;
43497	:douta	=	16'h	6a46;
43498	:douta	=	16'h	6226;
43499	:douta	=	16'h	59e5;
43500	:douta	=	16'h	59e5;
43501	:douta	=	16'h	59e5;
43502	:douta	=	16'h	59e6;
43503	:douta	=	16'h	59e6;
43504	:douta	=	16'h	51c6;
43505	:douta	=	16'h	51c6;
43506	:douta	=	16'h	51a5;
43507	:douta	=	16'h	49a5;
43508	:douta	=	16'h	49a5;
43509	:douta	=	16'h	49a6;
43510	:douta	=	16'h	49a6;
43511	:douta	=	16'h	49a6;
43512	:douta	=	16'h	49a6;
43513	:douta	=	16'h	4186;
43514	:douta	=	16'h	41a6;
43515	:douta	=	16'h	4186;
43516	:douta	=	16'h	4186;
43517	:douta	=	16'h	3965;
43518	:douta	=	16'h	3966;
43519	:douta	=	16'h	3986;
43520	:douta	=	16'h	ff3a;
43521	:douta	=	16'h	ff9c;
43522	:douta	=	16'h	ff9d;
43523	:douta	=	16'h	ffbc;
43524	:douta	=	16'h	ff9c;
43525	:douta	=	16'h	ffbd;
43526	:douta	=	16'h	de35;
43527	:douta	=	16'h	d5f5;
43528	:douta	=	16'h	d617;
43529	:douta	=	16'h	9c93;
43530	:douta	=	16'h	9c93;
43531	:douta	=	16'h	b556;
43532	:douta	=	16'h	b576;
43533	:douta	=	16'h	b535;
43534	:douta	=	16'h	b534;
43535	:douta	=	16'h	bd75;
43536	:douta	=	16'h	ad15;
43537	:douta	=	16'h	9cd5;
43538	:douta	=	16'h	8c75;
43539	:douta	=	16'h	7c34;
43540	:douta	=	16'h	8455;
43541	:douta	=	16'h	8475;
43542	:douta	=	16'h	8475;
43543	:douta	=	16'h	8455;
43544	:douta	=	16'h	8476;
43545	:douta	=	16'h	8475;
43546	:douta	=	16'h	8455;
43547	:douta	=	16'h	8475;
43548	:douta	=	16'h	7c13;
43549	:douta	=	16'h	7413;
43550	:douta	=	16'h	1082;
43551	:douta	=	16'h	2126;
43552	:douta	=	16'h	21c9;
43553	:douta	=	16'h	220c;
43554	:douta	=	16'h	2189;
43555	:douta	=	16'h	2168;
43556	:douta	=	16'h	18e5;
43557	:douta	=	16'h	18c3;
43558	:douta	=	16'h	1882;
43559	:douta	=	16'h	1861;
43560	:douta	=	16'h	1882;
43561	:douta	=	16'h	1882;
43562	:douta	=	16'h	1882;
43563	:douta	=	16'h	2082;
43564	:douta	=	16'h	20a2;
43565	:douta	=	16'h	20a2;
43566	:douta	=	16'h	20a2;
43567	:douta	=	16'h	20a2;
43568	:douta	=	16'h	20c2;
43569	:douta	=	16'h	28e2;
43570	:douta	=	16'h	28e2;
43571	:douta	=	16'h	2903;
43572	:douta	=	16'h	2946;
43573	:douta	=	16'h	1906;
43574	:douta	=	16'h	3103;
43575	:douta	=	16'h	4143;
43576	:douta	=	16'h	4144;
43577	:douta	=	16'h	4123;
43578	:douta	=	16'h	4143;
43579	:douta	=	16'h	4964;
43580	:douta	=	16'h	4963;
43581	:douta	=	16'h	4984;
43582	:douta	=	16'h	4984;
43583	:douta	=	16'h	59c4;
43584	:douta	=	16'h	3923;
43585	:douta	=	16'h	61c5;
43586	:douta	=	16'h	59c4;
43587	:douta	=	16'h	59c4;
43588	:douta	=	16'h	61e4;
43589	:douta	=	16'h	61e4;
43590	:douta	=	16'h	61e4;
43591	:douta	=	16'h	6a04;
43592	:douta	=	16'h	6a24;
43593	:douta	=	16'h	69e3;
43594	:douta	=	16'h	69e3;
43595	:douta	=	16'h	61a3;
43596	:douta	=	16'h	61a3;
43597	:douta	=	16'h	61a3;
43598	:douta	=	16'h	7244;
43599	:douta	=	16'h	8307;
43600	:douta	=	16'h	9369;
43601	:douta	=	16'h	a44c;
43602	:douta	=	16'h	b4ae;
43603	:douta	=	16'h	c5b1;
43604	:douta	=	16'h	de74;
43605	:douta	=	16'h	e6b5;
43606	:douta	=	16'h	e6b5;
43607	:douta	=	16'h	de94;
43608	:douta	=	16'h	d612;
43609	:douta	=	16'h	cdb0;
43610	:douta	=	16'h	c4ec;
43611	:douta	=	16'h	b429;
43612	:douta	=	16'h	b3e8;
43613	:douta	=	16'h	ab84;
43614	:douta	=	16'h	ab64;
43615	:douta	=	16'h	ab43;
43616	:douta	=	16'h	b343;
43617	:douta	=	16'h	b384;
43618	:douta	=	16'h	b364;
43619	:douta	=	16'h	bbc4;
43620	:douta	=	16'h	bbe5;
43621	:douta	=	16'h	c405;
43622	:douta	=	16'h	c405;
43623	:douta	=	16'h	c405;
43624	:douta	=	16'h	c406;
43625	:douta	=	16'h	c405;
43626	:douta	=	16'h	c426;
43627	:douta	=	16'h	c426;
43628	:douta	=	16'h	c425;
43629	:douta	=	16'h	c425;
43630	:douta	=	16'h	c425;
43631	:douta	=	16'h	c425;
43632	:douta	=	16'h	cc25;
43633	:douta	=	16'h	c405;
43634	:douta	=	16'h	c425;
43635	:douta	=	16'h	cc25;
43636	:douta	=	16'h	cc26;
43637	:douta	=	16'h	cc26;
43638	:douta	=	16'h	cc46;
43639	:douta	=	16'h	cc46;
43640	:douta	=	16'h	cc46;
43641	:douta	=	16'h	cc45;
43642	:douta	=	16'h	cc45;
43643	:douta	=	16'h	cc46;
43644	:douta	=	16'h	cc66;
43645	:douta	=	16'h	cc45;
43646	:douta	=	16'h	cc66;
43647	:douta	=	16'h	cc47;
43648	:douta	=	16'h	cc66;
43649	:douta	=	16'h	cc66;
43650	:douta	=	16'h	cc66;
43651	:douta	=	16'h	cc66;
43652	:douta	=	16'h	d466;
43653	:douta	=	16'h	cc66;
43654	:douta	=	16'h	cc66;
43655	:douta	=	16'h	d466;
43656	:douta	=	16'h	d466;
43657	:douta	=	16'h	cc66;
43658	:douta	=	16'h	d466;
43659	:douta	=	16'h	d466;
43660	:douta	=	16'h	d466;
43661	:douta	=	16'h	d466;
43662	:douta	=	16'h	d466;
43663	:douta	=	16'h	cc66;
43664	:douta	=	16'h	d466;
43665	:douta	=	16'h	d466;
43666	:douta	=	16'h	d467;
43667	:douta	=	16'h	d466;
43668	:douta	=	16'h	d467;
43669	:douta	=	16'h	d487;
43670	:douta	=	16'h	d467;
43671	:douta	=	16'h	d466;
43672	:douta	=	16'h	d466;
43673	:douta	=	16'h	d466;
43674	:douta	=	16'h	d466;
43675	:douta	=	16'h	d468;
43676	:douta	=	16'h	d466;
43677	:douta	=	16'h	cc68;
43678	:douta	=	16'h	dc84;
43679	:douta	=	16'h	cc69;
43680	:douta	=	16'h	7c12;
43681	:douta	=	16'h	7bd0;
43682	:douta	=	16'h	83b0;
43683	:douta	=	16'h	62ab;
43684	:douta	=	16'h	5249;
43685	:douta	=	16'h	6acb;
43686	:douta	=	16'h	acd0;
43687	:douta	=	16'h	a4b0;
43688	:douta	=	16'h	9c4e;
43689	:douta	=	16'h	c592;
43690	:douta	=	16'h	de35;
43691	:douta	=	16'h	83ac;
43692	:douta	=	16'h	f6f8;
43693	:douta	=	16'h	de16;
43694	:douta	=	16'h	de36;
43695	:douta	=	16'h	d615;
43696	:douta	=	16'h	de35;
43697	:douta	=	16'h	bd54;
43698	:douta	=	16'h	acd3;
43699	:douta	=	16'h	c575;
43700	:douta	=	16'h	b575;
43701	:douta	=	16'h	b536;
43702	:douta	=	16'h	acf5;
43703	:douta	=	16'h	9495;
43704	:douta	=	16'h	8c94;
43705	:douta	=	16'h	94b4;
43706	:douta	=	16'h	94b4;
43707	:douta	=	16'h	8c74;
43708	:douta	=	16'h	8453;
43709	:douta	=	16'h	7bf2;
43710	:douta	=	16'h	7bd1;
43711	:douta	=	16'h	7bf1;
43712	:douta	=	16'h	73d0;
43713	:douta	=	16'h	8412;
43714	:douta	=	16'h	7c12;
43715	:douta	=	16'h	5b2f;
43716	:douta	=	16'h	52cd;
43717	:douta	=	16'h	8412;
43718	:douta	=	16'h	7bf1;
43719	:douta	=	16'h	6b2c;
43720	:douta	=	16'h	3965;
43721	:douta	=	16'h	49e5;
43722	:douta	=	16'h	6ac9;
43723	:douta	=	16'h	62c9;
43724	:douta	=	16'h	5269;
43725	:douta	=	16'h	2903;
43726	:douta	=	16'h	49c6;
43727	:douta	=	16'h	acb0;
43728	:douta	=	16'h	cd93;
43729	:douta	=	16'h	c572;
43730	:douta	=	16'h	acaf;
43731	:douta	=	16'h	a46e;
43732	:douta	=	16'h	5aa9;
43733	:douta	=	16'h	6aaa;
43734	:douta	=	16'h	838c;
43735	:douta	=	16'h	bd31;
43736	:douta	=	16'h	cdd3;
43737	:douta	=	16'h	d614;
43738	:douta	=	16'h	b511;
43739	:douta	=	16'h	ac91;
43740	:douta	=	16'h	83cf;
43741	:douta	=	16'h	7b6f;
43742	:douta	=	16'h	6b4e;
43743	:douta	=	16'h	31c8;
43744	:douta	=	16'h	2126;
43745	:douta	=	16'h	2147;
43746	:douta	=	16'h	2126;
43747	:douta	=	16'h	2126;
43748	:douta	=	16'h	10e5;
43749	:douta	=	16'h	18e5;
43750	:douta	=	16'h	29a8;
43751	:douta	=	16'h	29a9;
43752	:douta	=	16'h	1926;
43753	:douta	=	16'h	6a46;
43754	:douta	=	16'h	6226;
43755	:douta	=	16'h	6206;
43756	:douta	=	16'h	59e5;
43757	:douta	=	16'h	59e5;
43758	:douta	=	16'h	59e6;
43759	:douta	=	16'h	59e6;
43760	:douta	=	16'h	51c5;
43761	:douta	=	16'h	51c5;
43762	:douta	=	16'h	51a5;
43763	:douta	=	16'h	4985;
43764	:douta	=	16'h	4985;
43765	:douta	=	16'h	4985;
43766	:douta	=	16'h	49a6;
43767	:douta	=	16'h	4986;
43768	:douta	=	16'h	49a6;
43769	:douta	=	16'h	4186;
43770	:douta	=	16'h	49a6;
43771	:douta	=	16'h	4186;
43772	:douta	=	16'h	4166;
43773	:douta	=	16'h	3966;
43774	:douta	=	16'h	3966;
43775	:douta	=	16'h	4166;
43776	:douta	=	16'h	f73a;
43777	:douta	=	16'h	ff9c;
43778	:douta	=	16'h	ff9c;
43779	:douta	=	16'h	ffbc;
43780	:douta	=	16'h	ffbd;
43781	:douta	=	16'h	ffdd;
43782	:douta	=	16'h	d593;
43783	:douta	=	16'h	d5b3;
43784	:douta	=	16'h	b555;
43785	:douta	=	16'h	9c73;
43786	:douta	=	16'h	b556;
43787	:douta	=	16'h	b556;
43788	:douta	=	16'h	b556;
43789	:douta	=	16'h	bd95;
43790	:douta	=	16'h	bd75;
43791	:douta	=	16'h	b555;
43792	:douta	=	16'h	a516;
43793	:douta	=	16'h	8c74;
43794	:douta	=	16'h	8c95;
43795	:douta	=	16'h	8454;
43796	:douta	=	16'h	8455;
43797	:douta	=	16'h	8475;
43798	:douta	=	16'h	8c96;
43799	:douta	=	16'h	7c34;
43800	:douta	=	16'h	8496;
43801	:douta	=	16'h	7c55;
43802	:douta	=	16'h	7c34;
43803	:douta	=	16'h	8454;
43804	:douta	=	16'h	94d6;
43805	:douta	=	16'h	1020;
43806	:douta	=	16'h	1882;
43807	:douta	=	16'h	18c3;
43808	:douta	=	16'h	20a3;
43809	:douta	=	16'h	1041;
43810	:douta	=	16'h	1061;
43811	:douta	=	16'h	1861;
43812	:douta	=	16'h	1882;
43813	:douta	=	16'h	1882;
43814	:douta	=	16'h	1862;
43815	:douta	=	16'h	1883;
43816	:douta	=	16'h	18a2;
43817	:douta	=	16'h	1882;
43818	:douta	=	16'h	18a2;
43819	:douta	=	16'h	20a2;
43820	:douta	=	16'h	20a2;
43821	:douta	=	16'h	20a2;
43822	:douta	=	16'h	20a2;
43823	:douta	=	16'h	28c3;
43824	:douta	=	16'h	20c2;
43825	:douta	=	16'h	28e2;
43826	:douta	=	16'h	28e3;
43827	:douta	=	16'h	2904;
43828	:douta	=	16'h	2947;
43829	:douta	=	16'h	18e5;
43830	:douta	=	16'h	3903;
43831	:douta	=	16'h	3903;
43832	:douta	=	16'h	4124;
43833	:douta	=	16'h	4143;
43834	:douta	=	16'h	4163;
43835	:douta	=	16'h	4964;
43836	:douta	=	16'h	4984;
43837	:douta	=	16'h	4984;
43838	:douta	=	16'h	49a4;
43839	:douta	=	16'h	5984;
43840	:douta	=	16'h	30e2;
43841	:douta	=	16'h	5163;
43842	:douta	=	16'h	5162;
43843	:douta	=	16'h	5983;
43844	:douta	=	16'h	59c3;
43845	:douta	=	16'h	6a46;
43846	:douta	=	16'h	72a7;
43847	:douta	=	16'h	8329;
43848	:douta	=	16'h	8b8a;
43849	:douta	=	16'h	acae;
43850	:douta	=	16'h	bd50;
43851	:douta	=	16'h	bd91;
43852	:douta	=	16'h	c5d2;
43853	:douta	=	16'h	c5d1;
43854	:douta	=	16'h	c591;
43855	:douta	=	16'h	b4ee;
43856	:douta	=	16'h	ac6c;
43857	:douta	=	16'h	a40a;
43858	:douta	=	16'h	9bc9;
43859	:douta	=	16'h	9306;
43860	:douta	=	16'h	8ac3;
43861	:douta	=	16'h	8aa2;
43862	:douta	=	16'h	92a2;
43863	:douta	=	16'h	9282;
43864	:douta	=	16'h	9b04;
43865	:douta	=	16'h	9b04;
43866	:douta	=	16'h	a345;
43867	:douta	=	16'h	ab85;
43868	:douta	=	16'h	a364;
43869	:douta	=	16'h	ab85;
43870	:douta	=	16'h	ab65;
43871	:douta	=	16'h	b3a5;
43872	:douta	=	16'h	b3a5;
43873	:douta	=	16'h	b3a4;
43874	:douta	=	16'h	bbc4;
43875	:douta	=	16'h	c405;
43876	:douta	=	16'h	bbe5;
43877	:douta	=	16'h	c405;
43878	:douta	=	16'h	c405;
43879	:douta	=	16'h	c405;
43880	:douta	=	16'h	c406;
43881	:douta	=	16'h	c425;
43882	:douta	=	16'h	c425;
43883	:douta	=	16'h	c425;
43884	:douta	=	16'h	c425;
43885	:douta	=	16'h	c445;
43886	:douta	=	16'h	c425;
43887	:douta	=	16'h	c425;
43888	:douta	=	16'h	c425;
43889	:douta	=	16'h	c425;
43890	:douta	=	16'h	c425;
43891	:douta	=	16'h	cc25;
43892	:douta	=	16'h	cc25;
43893	:douta	=	16'h	cc26;
43894	:douta	=	16'h	cc46;
43895	:douta	=	16'h	cc26;
43896	:douta	=	16'h	cc45;
43897	:douta	=	16'h	cc45;
43898	:douta	=	16'h	cc45;
43899	:douta	=	16'h	cc46;
43900	:douta	=	16'h	cc45;
43901	:douta	=	16'h	cc46;
43902	:douta	=	16'h	cc66;
43903	:douta	=	16'h	cc46;
43904	:douta	=	16'h	cc47;
43905	:douta	=	16'h	cc47;
43906	:douta	=	16'h	cc66;
43907	:douta	=	16'h	cc66;
43908	:douta	=	16'h	cc66;
43909	:douta	=	16'h	cc66;
43910	:douta	=	16'h	cc66;
43911	:douta	=	16'h	cc66;
43912	:douta	=	16'h	d467;
43913	:douta	=	16'h	d467;
43914	:douta	=	16'h	d466;
43915	:douta	=	16'h	cc66;
43916	:douta	=	16'h	d466;
43917	:douta	=	16'h	d467;
43918	:douta	=	16'h	d467;
43919	:douta	=	16'h	d467;
43920	:douta	=	16'h	d466;
43921	:douta	=	16'h	cc66;
43922	:douta	=	16'h	d466;
43923	:douta	=	16'h	d466;
43924	:douta	=	16'h	d466;
43925	:douta	=	16'h	d466;
43926	:douta	=	16'h	d466;
43927	:douta	=	16'h	d467;
43928	:douta	=	16'h	d466;
43929	:douta	=	16'h	d466;
43930	:douta	=	16'h	d466;
43931	:douta	=	16'h	d467;
43932	:douta	=	16'h	d467;
43933	:douta	=	16'h	cc66;
43934	:douta	=	16'h	cc86;
43935	:douta	=	16'h	d487;
43936	:douta	=	16'h	cc89;
43937	:douta	=	16'h	9c4f;
43938	:douta	=	16'h	940d;
43939	:douta	=	16'h	9c4e;
43940	:douta	=	16'h	acb0;
43941	:douta	=	16'h	bd31;
43942	:douta	=	16'h	bd51;
43943	:douta	=	16'h	c573;
43944	:douta	=	16'h	e676;
43945	:douta	=	16'h	eeb7;
43946	:douta	=	16'h	9c0f;
43947	:douta	=	16'h	de16;
43948	:douta	=	16'h	d5f5;
43949	:douta	=	16'h	d615;
43950	:douta	=	16'h	d615;
43951	:douta	=	16'h	cdd5;
43952	:douta	=	16'h	cdd6;
43953	:douta	=	16'h	cdb5;
43954	:douta	=	16'h	a4b3;
43955	:douta	=	16'h	a4d3;
43956	:douta	=	16'h	a4f5;
43957	:douta	=	16'h	9cd5;
43958	:douta	=	16'h	8c94;
43959	:douta	=	16'h	9494;
43960	:douta	=	16'h	8433;
43961	:douta	=	16'h	7bd1;
43962	:douta	=	16'h	8c74;
43963	:douta	=	16'h	7bf2;
43964	:douta	=	16'h	7bd1;
43965	:douta	=	16'h	7bd1;
43966	:douta	=	16'h	73b1;
43967	:douta	=	16'h	73d1;
43968	:douta	=	16'h	634e;
43969	:douta	=	16'h	73d1;
43970	:douta	=	16'h	6b6f;
43971	:douta	=	16'h	4a28;
43972	:douta	=	16'h	41a8;
43973	:douta	=	16'h	3964;
43974	:douta	=	16'h	5247;
43975	:douta	=	16'h	83cd;
43976	:douta	=	16'h	942e;
43977	:douta	=	16'h	7bac;
43978	:douta	=	16'h	7b8b;
43979	:douta	=	16'h	b4f1;
43980	:douta	=	16'h	c551;
43981	:douta	=	16'h	b531;
43982	:douta	=	16'h	acd0;
43983	:douta	=	16'h	83ac;
43984	:douta	=	16'h	730b;
43985	:douta	=	16'h	83ad;
43986	:douta	=	16'h	cd93;
43987	:douta	=	16'h	d5d4;
43988	:douta	=	16'h	de36;
43989	:douta	=	16'h	cdb2;
43990	:douta	=	16'h	bd31;
43991	:douta	=	16'h	9c6f;
43992	:douta	=	16'h	ac6f;
43993	:douta	=	16'h	b512;
43994	:douta	=	16'h	c532;
43995	:douta	=	16'h	acd2;
43996	:douta	=	16'h	8431;
43997	:douta	=	16'h	7bd1;
43998	:douta	=	16'h	6b4f;
43999	:douta	=	16'h	4ace;
44000	:douta	=	16'h	4a8d;
44001	:douta	=	16'h	3a0a;
44002	:douta	=	16'h	3a0a;
44003	:douta	=	16'h	18e5;
44004	:douta	=	16'h	52ee;
44005	:douta	=	16'h	2968;
44006	:douta	=	16'h	1906;
44007	:douta	=	16'h	1926;
44008	:douta	=	16'h	1927;
44009	:douta	=	16'h	6a26;
44010	:douta	=	16'h	6226;
44011	:douta	=	16'h	59e6;
44012	:douta	=	16'h	6206;
44013	:douta	=	16'h	59e6;
44014	:douta	=	16'h	59e6;
44015	:douta	=	16'h	51c5;
44016	:douta	=	16'h	51c6;
44017	:douta	=	16'h	51c5;
44018	:douta	=	16'h	51a5;
44019	:douta	=	16'h	49a5;
44020	:douta	=	16'h	49a5;
44021	:douta	=	16'h	49a5;
44022	:douta	=	16'h	49a5;
44023	:douta	=	16'h	4986;
44024	:douta	=	16'h	4185;
44025	:douta	=	16'h	4186;
44026	:douta	=	16'h	4185;
44027	:douta	=	16'h	4186;
44028	:douta	=	16'h	4186;
44029	:douta	=	16'h	4186;
44030	:douta	=	16'h	4166;
44031	:douta	=	16'h	3986;
44032	:douta	=	16'h	ff5a;
44033	:douta	=	16'h	ff7c;
44034	:douta	=	16'h	ff9c;
44035	:douta	=	16'h	ff9c;
44036	:douta	=	16'h	ff7b;
44037	:douta	=	16'h	ffdc;
44038	:douta	=	16'h	cd94;
44039	:douta	=	16'h	ee78;
44040	:douta	=	16'h	ad35;
44041	:douta	=	16'h	9c93;
44042	:douta	=	16'h	b576;
44043	:douta	=	16'h	bd97;
44044	:douta	=	16'h	bd77;
44045	:douta	=	16'h	bd95;
44046	:douta	=	16'h	bd95;
44047	:douta	=	16'h	b555;
44048	:douta	=	16'h	9cf6;
44049	:douta	=	16'h	8454;
44050	:douta	=	16'h	8c74;
44051	:douta	=	16'h	8475;
44052	:douta	=	16'h	8454;
44053	:douta	=	16'h	8475;
44054	:douta	=	16'h	8496;
44055	:douta	=	16'h	7c54;
44056	:douta	=	16'h	8475;
44057	:douta	=	16'h	7c55;
44058	:douta	=	16'h	8454;
44059	:douta	=	16'h	8433;
44060	:douta	=	16'h	8454;
44061	:douta	=	16'h	1040;
44062	:douta	=	16'h	20c3;
44063	:douta	=	16'h	18a2;
44064	:douta	=	16'h	18a3;
44065	:douta	=	16'h	1861;
44066	:douta	=	16'h	1882;
44067	:douta	=	16'h	1082;
44068	:douta	=	16'h	1882;
44069	:douta	=	16'h	1861;
44070	:douta	=	16'h	18a2;
44071	:douta	=	16'h	1882;
44072	:douta	=	16'h	1882;
44073	:douta	=	16'h	1882;
44074	:douta	=	16'h	2082;
44075	:douta	=	16'h	20a2;
44076	:douta	=	16'h	20a2;
44077	:douta	=	16'h	20a2;
44078	:douta	=	16'h	20c2;
44079	:douta	=	16'h	20c2;
44080	:douta	=	16'h	28e2;
44081	:douta	=	16'h	28e2;
44082	:douta	=	16'h	30e2;
44083	:douta	=	16'h	2924;
44084	:douta	=	16'h	2967;
44085	:douta	=	16'h	18e5;
44086	:douta	=	16'h	3923;
44087	:douta	=	16'h	3923;
44088	:douta	=	16'h	4143;
44089	:douta	=	16'h	4123;
44090	:douta	=	16'h	4123;
44091	:douta	=	16'h	4122;
44092	:douta	=	16'h	4122;
44093	:douta	=	16'h	4922;
44094	:douta	=	16'h	4922;
44095	:douta	=	16'h	5184;
44096	:douta	=	16'h	3924;
44097	:douta	=	16'h	59e5;
44098	:douta	=	16'h	8329;
44099	:douta	=	16'h	8bab;
44100	:douta	=	16'h	944d;
44101	:douta	=	16'h	acf0;
44102	:douta	=	16'h	b531;
44103	:douta	=	16'h	bd72;
44104	:douta	=	16'h	bd71;
44105	:douta	=	16'h	bd30;
44106	:douta	=	16'h	ac8e;
44107	:douta	=	16'h	9c2c;
44108	:douta	=	16'h	8b69;
44109	:douta	=	16'h	8b27;
44110	:douta	=	16'h	82c6;
44111	:douta	=	16'h	7a63;
44112	:douta	=	16'h	7a43;
44113	:douta	=	16'h	7a43;
44114	:douta	=	16'h	8244;
44115	:douta	=	16'h	8284;
44116	:douta	=	16'h	8ac5;
44117	:douta	=	16'h	92c4;
44118	:douta	=	16'h	9b05;
44119	:douta	=	16'h	9b05;
44120	:douta	=	16'h	a325;
44121	:douta	=	16'h	9b25;
44122	:douta	=	16'h	a345;
44123	:douta	=	16'h	ab65;
44124	:douta	=	16'h	ab65;
44125	:douta	=	16'h	ab85;
44126	:douta	=	16'h	ab85;
44127	:douta	=	16'h	b3a5;
44128	:douta	=	16'h	b3a5;
44129	:douta	=	16'h	b3a5;
44130	:douta	=	16'h	bc05;
44131	:douta	=	16'h	c406;
44132	:douta	=	16'h	c406;
44133	:douta	=	16'h	bc06;
44134	:douta	=	16'h	c406;
44135	:douta	=	16'h	c405;
44136	:douta	=	16'h	c405;
44137	:douta	=	16'h	cc46;
44138	:douta	=	16'h	cc66;
44139	:douta	=	16'h	c446;
44140	:douta	=	16'h	cc46;
44141	:douta	=	16'h	cc46;
44142	:douta	=	16'h	c405;
44143	:douta	=	16'h	c405;
44144	:douta	=	16'h	c405;
44145	:douta	=	16'h	c405;
44146	:douta	=	16'h	cc25;
44147	:douta	=	16'h	cc46;
44148	:douta	=	16'h	cc25;
44149	:douta	=	16'h	cc46;
44150	:douta	=	16'h	cc25;
44151	:douta	=	16'h	cc26;
44152	:douta	=	16'h	cc45;
44153	:douta	=	16'h	cc45;
44154	:douta	=	16'h	cc45;
44155	:douta	=	16'h	cc46;
44156	:douta	=	16'h	cc45;
44157	:douta	=	16'h	cc46;
44158	:douta	=	16'h	cc46;
44159	:douta	=	16'h	cc66;
44160	:douta	=	16'h	d467;
44161	:douta	=	16'h	cc47;
44162	:douta	=	16'h	cc47;
44163	:douta	=	16'h	cc47;
44164	:douta	=	16'h	d466;
44165	:douta	=	16'h	cc66;
44166	:douta	=	16'h	cc66;
44167	:douta	=	16'h	cc66;
44168	:douta	=	16'h	d467;
44169	:douta	=	16'h	d467;
44170	:douta	=	16'h	cc66;
44171	:douta	=	16'h	cc66;
44172	:douta	=	16'h	d466;
44173	:douta	=	16'h	d466;
44174	:douta	=	16'h	d467;
44175	:douta	=	16'h	d467;
44176	:douta	=	16'h	d467;
44177	:douta	=	16'h	d466;
44178	:douta	=	16'h	d467;
44179	:douta	=	16'h	d466;
44180	:douta	=	16'h	d487;
44181	:douta	=	16'h	d467;
44182	:douta	=	16'h	d467;
44183	:douta	=	16'h	d467;
44184	:douta	=	16'h	d467;
44185	:douta	=	16'h	d467;
44186	:douta	=	16'h	d467;
44187	:douta	=	16'h	d467;
44188	:douta	=	16'h	d487;
44189	:douta	=	16'h	d486;
44190	:douta	=	16'h	d468;
44191	:douta	=	16'h	d467;
44192	:douta	=	16'h	d466;
44193	:douta	=	16'h	b4d0;
44194	:douta	=	16'h	ac8f;
44195	:douta	=	16'h	bd11;
44196	:douta	=	16'h	bd11;
44197	:douta	=	16'h	d5f4;
44198	:douta	=	16'h	c592;
44199	:douta	=	16'h	d5f4;
44200	:douta	=	16'h	e697;
44201	:douta	=	16'h	d635;
44202	:douta	=	16'h	bd31;
44203	:douta	=	16'h	eeb7;
44204	:douta	=	16'h	d5f6;
44205	:douta	=	16'h	d5b6;
44206	:douta	=	16'h	d5d5;
44207	:douta	=	16'h	cdb5;
44208	:douta	=	16'h	c596;
44209	:douta	=	16'h	c576;
44210	:douta	=	16'h	9c93;
44211	:douta	=	16'h	9c73;
44212	:douta	=	16'h	9494;
44213	:douta	=	16'h	8c94;
44214	:douta	=	16'h	8c53;
44215	:douta	=	16'h	8433;
44216	:douta	=	16'h	8412;
44217	:douta	=	16'h	7bb1;
44218	:douta	=	16'h	7bf2;
44219	:douta	=	16'h	8433;
44220	:douta	=	16'h	7390;
44221	:douta	=	16'h	7bd1;
44222	:douta	=	16'h	6b90;
44223	:douta	=	16'h	73b1;
44224	:douta	=	16'h	6b90;
44225	:douta	=	16'h	5acb;
44226	:douta	=	16'h	5228;
44227	:douta	=	16'h	3143;
44228	:douta	=	16'h	49c5;
44229	:douta	=	16'h	6aeb;
44230	:douta	=	16'h	732c;
44231	:douta	=	16'h	7b6c;
44232	:douta	=	16'h	b510;
44233	:douta	=	16'h	a48f;
44234	:douta	=	16'h	9c2e;
44235	:douta	=	16'h	9c4f;
44236	:douta	=	16'h	b4d0;
44237	:douta	=	16'h	cdd3;
44238	:douta	=	16'h	cdd3;
44239	:douta	=	16'h	cdb3;
44240	:douta	=	16'h	a46f;
44241	:douta	=	16'h	8bee;
44242	:douta	=	16'h	a46e;
44243	:douta	=	16'h	c551;
44244	:douta	=	16'h	d5f4;
44245	:douta	=	16'h	e636;
44246	:douta	=	16'h	e615;
44247	:douta	=	16'h	d5d4;
44248	:douta	=	16'h	cd73;
44249	:douta	=	16'h	b512;
44250	:douta	=	16'h	acd2;
44251	:douta	=	16'h	acb1;
44252	:douta	=	16'h	8c73;
44253	:douta	=	16'h	7bf1;
44254	:douta	=	16'h	6b6f;
44255	:douta	=	16'h	52ce;
44256	:douta	=	16'h	4a8d;
44257	:douta	=	16'h	39ea;
44258	:douta	=	16'h	3a2b;
44259	:douta	=	16'h	2167;
44260	:douta	=	16'h	3a0a;
44261	:douta	=	16'h	31ea;
44262	:douta	=	16'h	1926;
44263	:douta	=	16'h	2126;
44264	:douta	=	16'h	2188;
44265	:douta	=	16'h	5a27;
44266	:douta	=	16'h	6a46;
44267	:douta	=	16'h	6206;
44268	:douta	=	16'h	5a06;
44269	:douta	=	16'h	59e6;
44270	:douta	=	16'h	59c6;
44271	:douta	=	16'h	51e5;
44272	:douta	=	16'h	51c6;
44273	:douta	=	16'h	51c5;
44274	:douta	=	16'h	49a5;
44275	:douta	=	16'h	4985;
44276	:douta	=	16'h	49a5;
44277	:douta	=	16'h	49a5;
44278	:douta	=	16'h	49a5;
44279	:douta	=	16'h	49a6;
44280	:douta	=	16'h	4185;
44281	:douta	=	16'h	4186;
44282	:douta	=	16'h	41a6;
44283	:douta	=	16'h	4186;
44284	:douta	=	16'h	4186;
44285	:douta	=	16'h	3965;
44286	:douta	=	16'h	3986;
44287	:douta	=	16'h	3986;
44288	:douta	=	16'h	ff7b;
44289	:douta	=	16'h	ff9c;
44290	:douta	=	16'h	ffbc;
44291	:douta	=	16'h	ff9c;
44292	:douta	=	16'h	fffe;
44293	:douta	=	16'h	e6b8;
44294	:douta	=	16'h	ee98;
44295	:douta	=	16'h	e657;
44296	:douta	=	16'h	9c93;
44297	:douta	=	16'h	ad36;
44298	:douta	=	16'h	bd97;
44299	:douta	=	16'h	b556;
44300	:douta	=	16'h	bd56;
44301	:douta	=	16'h	c596;
44302	:douta	=	16'h	bd95;
44303	:douta	=	16'h	ad55;
44304	:douta	=	16'h	8c75;
44305	:douta	=	16'h	8cb6;
44306	:douta	=	16'h	8454;
44307	:douta	=	16'h	8475;
44308	:douta	=	16'h	8c75;
44309	:douta	=	16'h	8454;
44310	:douta	=	16'h	8475;
44311	:douta	=	16'h	8495;
44312	:douta	=	16'h	7c54;
44313	:douta	=	16'h	8433;
44314	:douta	=	16'h	7c13;
44315	:douta	=	16'h	94f7;
44316	:douta	=	16'h	0841;
44317	:douta	=	16'h	18a3;
44318	:douta	=	16'h	20e3;
44319	:douta	=	16'h	18a3;
44320	:douta	=	16'h	20c3;
44321	:douta	=	16'h	1061;
44322	:douta	=	16'h	1082;
44323	:douta	=	16'h	18a2;
44324	:douta	=	16'h	1082;
44325	:douta	=	16'h	1882;
44326	:douta	=	16'h	1862;
44327	:douta	=	16'h	1882;
44328	:douta	=	16'h	1882;
44329	:douta	=	16'h	20a2;
44330	:douta	=	16'h	1882;
44331	:douta	=	16'h	20a2;
44332	:douta	=	16'h	20a2;
44333	:douta	=	16'h	2082;
44334	:douta	=	16'h	20c2;
44335	:douta	=	16'h	28c2;
44336	:douta	=	16'h	20c2;
44337	:douta	=	16'h	28c2;
44338	:douta	=	16'h	28a1;
44339	:douta	=	16'h	2925;
44340	:douta	=	16'h	2987;
44341	:douta	=	16'h	18c4;
44342	:douta	=	16'h	4184;
44343	:douta	=	16'h	49a5;
44344	:douta	=	16'h	62a8;
44345	:douta	=	16'h	62ca;
44346	:douta	=	16'h	7b8d;
44347	:douta	=	16'h	8c2f;
44348	:douta	=	16'h	9490;
44349	:douta	=	16'h	9490;
44350	:douta	=	16'h	9c8f;
44351	:douta	=	16'h	8c2e;
44352	:douta	=	16'h	8c2e;
44353	:douta	=	16'h	6a87;
44354	:douta	=	16'h	7ae8;
44355	:douta	=	16'h	72a7;
44356	:douta	=	16'h	6a24;
44357	:douta	=	16'h	61e4;
44358	:douta	=	16'h	6a04;
44359	:douta	=	16'h	61a3;
44360	:douta	=	16'h	69c3;
44361	:douta	=	16'h	6a04;
44362	:douta	=	16'h	6a03;
44363	:douta	=	16'h	7203;
44364	:douta	=	16'h	7224;
44365	:douta	=	16'h	7244;
44366	:douta	=	16'h	7a64;
44367	:douta	=	16'h	7a63;
44368	:douta	=	16'h	8284;
44369	:douta	=	16'h	82a4;
44370	:douta	=	16'h	8aa4;
44371	:douta	=	16'h	8ac4;
44372	:douta	=	16'h	92e4;
44373	:douta	=	16'h	92e5;
44374	:douta	=	16'h	9b05;
44375	:douta	=	16'h	9b25;
44376	:douta	=	16'h	9b24;
44377	:douta	=	16'h	a325;
44378	:douta	=	16'h	a345;
44379	:douta	=	16'h	ab64;
44380	:douta	=	16'h	ab64;
44381	:douta	=	16'h	ab65;
44382	:douta	=	16'h	ab65;
44383	:douta	=	16'h	ab84;
44384	:douta	=	16'h	b3a5;
44385	:douta	=	16'h	bbc6;
44386	:douta	=	16'h	bbe5;
44387	:douta	=	16'h	c406;
44388	:douta	=	16'h	c426;
44389	:douta	=	16'h	c405;
44390	:douta	=	16'h	bbe5;
44391	:douta	=	16'h	c426;
44392	:douta	=	16'h	c426;
44393	:douta	=	16'h	c425;
44394	:douta	=	16'h	c425;
44395	:douta	=	16'h	c425;
44396	:douta	=	16'h	cc46;
44397	:douta	=	16'h	c405;
44398	:douta	=	16'h	c405;
44399	:douta	=	16'h	c425;
44400	:douta	=	16'h	c425;
44401	:douta	=	16'h	cc26;
44402	:douta	=	16'h	c425;
44403	:douta	=	16'h	cc26;
44404	:douta	=	16'h	cc26;
44405	:douta	=	16'h	cc25;
44406	:douta	=	16'h	cc46;
44407	:douta	=	16'h	cc46;
44408	:douta	=	16'h	cc46;
44409	:douta	=	16'h	cc46;
44410	:douta	=	16'h	cc46;
44411	:douta	=	16'h	cc46;
44412	:douta	=	16'h	cc46;
44413	:douta	=	16'h	cc46;
44414	:douta	=	16'h	cc66;
44415	:douta	=	16'h	cc46;
44416	:douta	=	16'h	cc66;
44417	:douta	=	16'h	cc46;
44418	:douta	=	16'h	d467;
44419	:douta	=	16'h	d467;
44420	:douta	=	16'h	cc66;
44421	:douta	=	16'h	cc66;
44422	:douta	=	16'h	d467;
44423	:douta	=	16'h	d467;
44424	:douta	=	16'h	d467;
44425	:douta	=	16'h	d467;
44426	:douta	=	16'h	d467;
44427	:douta	=	16'h	cc66;
44428	:douta	=	16'h	d466;
44429	:douta	=	16'h	d466;
44430	:douta	=	16'h	d466;
44431	:douta	=	16'h	d467;
44432	:douta	=	16'h	d467;
44433	:douta	=	16'h	d467;
44434	:douta	=	16'h	cc66;
44435	:douta	=	16'h	d467;
44436	:douta	=	16'h	d467;
44437	:douta	=	16'h	d467;
44438	:douta	=	16'h	d467;
44439	:douta	=	16'h	d467;
44440	:douta	=	16'h	d467;
44441	:douta	=	16'h	d467;
44442	:douta	=	16'h	d467;
44443	:douta	=	16'h	d467;
44444	:douta	=	16'h	d467;
44445	:douta	=	16'h	d467;
44446	:douta	=	16'h	d487;
44447	:douta	=	16'h	d467;
44448	:douta	=	16'h	d467;
44449	:douta	=	16'h	c448;
44450	:douta	=	16'h	9c2e;
44451	:douta	=	16'h	acb1;
44452	:douta	=	16'h	b4d2;
44453	:douta	=	16'h	d5d4;
44454	:douta	=	16'h	c573;
44455	:douta	=	16'h	cdb4;
44456	:douta	=	16'h	d636;
44457	:douta	=	16'h	c574;
44458	:douta	=	16'h	d5f5;
44459	:douta	=	16'h	c555;
44460	:douta	=	16'h	bd76;
44461	:douta	=	16'h	c576;
44462	:douta	=	16'h	b556;
44463	:douta	=	16'h	b536;
44464	:douta	=	16'h	a516;
44465	:douta	=	16'h	9cf6;
44466	:douta	=	16'h	73d1;
44467	:douta	=	16'h	7c12;
44468	:douta	=	16'h	7bf1;
44469	:douta	=	16'h	8432;
44470	:douta	=	16'h	8452;
44471	:douta	=	16'h	73b0;
44472	:douta	=	16'h	8432;
44473	:douta	=	16'h	7bd1;
44474	:douta	=	16'h	7bd1;
44475	:douta	=	16'h	6b90;
44476	:douta	=	16'h	73b1;
44477	:douta	=	16'h	630e;
44478	:douta	=	16'h	41a6;
44479	:douta	=	16'h	41c6;
44480	:douta	=	16'h	49c6;
44481	:douta	=	16'h	732c;
44482	:douta	=	16'h	7b4c;
44483	:douta	=	16'h	8bed;
44484	:douta	=	16'h	8bcd;
44485	:douta	=	16'h	b530;
44486	:douta	=	16'h	bd51;
44487	:douta	=	16'h	9c4f;
44488	:douta	=	16'h	8bed;
44489	:douta	=	16'h	c531;
44490	:douta	=	16'h	c572;
44491	:douta	=	16'h	bd51;
44492	:douta	=	16'h	bd31;
44493	:douta	=	16'h	b4f0;
44494	:douta	=	16'h	c572;
44495	:douta	=	16'h	d635;
44496	:douta	=	16'h	de35;
44497	:douta	=	16'h	de56;
44498	:douta	=	16'h	e656;
44499	:douta	=	16'h	d5f4;
44500	:douta	=	16'h	d5b4;
44501	:douta	=	16'h	d5b3;
44502	:douta	=	16'h	cd93;
44503	:douta	=	16'h	c553;
44504	:douta	=	16'h	c553;
44505	:douta	=	16'h	acf3;
44506	:douta	=	16'h	9493;
44507	:douta	=	16'h	9493;
44508	:douta	=	16'h	8432;
44509	:douta	=	16'h	8412;
44510	:douta	=	16'h	73b1;
44511	:douta	=	16'h	5b4f;
44512	:douta	=	16'h	5b2f;
44513	:douta	=	16'h	52ce;
44514	:douta	=	16'h	4a8c;
44515	:douta	=	16'h	424c;
44516	:douta	=	16'h	18e5;
44517	:douta	=	16'h	5aac;
44518	:douta	=	16'h	08a3;
44519	:douta	=	16'h	18e5;
44520	:douta	=	16'h	2125;
44521	:douta	=	16'h	2127;
44522	:douta	=	16'h	59e6;
44523	:douta	=	16'h	6205;
44524	:douta	=	16'h	59e6;
44525	:douta	=	16'h	59e6;
44526	:douta	=	16'h	51c6;
44527	:douta	=	16'h	51e5;
44528	:douta	=	16'h	51c5;
44529	:douta	=	16'h	51a5;
44530	:douta	=	16'h	49a5;
44531	:douta	=	16'h	49a5;
44532	:douta	=	16'h	49a6;
44533	:douta	=	16'h	49a6;
44534	:douta	=	16'h	49a5;
44535	:douta	=	16'h	49a6;
44536	:douta	=	16'h	4186;
44537	:douta	=	16'h	49a6;
44538	:douta	=	16'h	4185;
44539	:douta	=	16'h	4186;
44540	:douta	=	16'h	4165;
44541	:douta	=	16'h	4186;
44542	:douta	=	16'h	3966;
44543	:douta	=	16'h	3966;
44544	:douta	=	16'h	ff7b;
44545	:douta	=	16'h	ffbd;
44546	:douta	=	16'h	ffbd;
44547	:douta	=	16'h	ffbc;
44548	:douta	=	16'h	ff7c;
44549	:douta	=	16'h	de15;
44550	:douta	=	16'h	ee98;
44551	:douta	=	16'h	d616;
44552	:douta	=	16'h	9c93;
44553	:douta	=	16'h	bd97;
44554	:douta	=	16'h	b596;
44555	:douta	=	16'h	b576;
44556	:douta	=	16'h	b555;
44557	:douta	=	16'h	c596;
44558	:douta	=	16'h	bd75;
44559	:douta	=	16'h	ad36;
44560	:douta	=	16'h	8474;
44561	:douta	=	16'h	8cb5;
44562	:douta	=	16'h	8454;
44563	:douta	=	16'h	8455;
44564	:douta	=	16'h	8475;
44565	:douta	=	16'h	8475;
44566	:douta	=	16'h	8475;
44567	:douta	=	16'h	8496;
44568	:douta	=	16'h	7c54;
44569	:douta	=	16'h	8433;
44570	:douta	=	16'h	8c96;
44571	:douta	=	16'h	8c96;
44572	:douta	=	16'h	1020;
44573	:douta	=	16'h	20c3;
44574	:douta	=	16'h	20c3;
44575	:douta	=	16'h	18a2;
44576	:douta	=	16'h	18c3;
44577	:douta	=	16'h	1062;
44578	:douta	=	16'h	1882;
44579	:douta	=	16'h	1882;
44580	:douta	=	16'h	1882;
44581	:douta	=	16'h	1882;
44582	:douta	=	16'h	1882;
44583	:douta	=	16'h	1882;
44584	:douta	=	16'h	1882;
44585	:douta	=	16'h	2082;
44586	:douta	=	16'h	2082;
44587	:douta	=	16'h	20a2;
44588	:douta	=	16'h	2082;
44589	:douta	=	16'h	2081;
44590	:douta	=	16'h	2081;
44591	:douta	=	16'h	2081;
44592	:douta	=	16'h	28c2;
44593	:douta	=	16'h	3103;
44594	:douta	=	16'h	3124;
44595	:douta	=	16'h	2967;
44596	:douta	=	16'h	2967;
44597	:douta	=	16'h	18c3;
44598	:douta	=	16'h	7bae;
44599	:douta	=	16'h	7bae;
44600	:douta	=	16'h	840f;
44601	:douta	=	16'h	8c2f;
44602	:douta	=	16'h	83cd;
44603	:douta	=	16'h	734a;
44604	:douta	=	16'h	6ae9;
44605	:douta	=	16'h	6286;
44606	:douta	=	16'h	6245;
44607	:douta	=	16'h	6aa8;
44608	:douta	=	16'h	83cc;
44609	:douta	=	16'h	3102;
44610	:douta	=	16'h	5983;
44611	:douta	=	16'h	5983;
44612	:douta	=	16'h	61a3;
44613	:douta	=	16'h	61e3;
44614	:douta	=	16'h	61e4;
44615	:douta	=	16'h	6a04;
44616	:douta	=	16'h	6a24;
44617	:douta	=	16'h	7244;
44618	:douta	=	16'h	7223;
44619	:douta	=	16'h	7223;
44620	:douta	=	16'h	7244;
44621	:douta	=	16'h	7244;
44622	:douta	=	16'h	7a64;
44623	:douta	=	16'h	7a63;
44624	:douta	=	16'h	8284;
44625	:douta	=	16'h	82a4;
44626	:douta	=	16'h	8aa4;
44627	:douta	=	16'h	8ac4;
44628	:douta	=	16'h	92e5;
44629	:douta	=	16'h	9305;
44630	:douta	=	16'h	9b05;
44631	:douta	=	16'h	9b26;
44632	:douta	=	16'h	9b25;
44633	:douta	=	16'h	a325;
44634	:douta	=	16'h	a345;
44635	:douta	=	16'h	ab64;
44636	:douta	=	16'h	ab65;
44637	:douta	=	16'h	ab65;
44638	:douta	=	16'h	b385;
44639	:douta	=	16'h	b385;
44640	:douta	=	16'h	bbc6;
44641	:douta	=	16'h	bbc5;
44642	:douta	=	16'h	bc05;
44643	:douta	=	16'h	bbe5;
44644	:douta	=	16'h	bbe5;
44645	:douta	=	16'h	bc06;
44646	:douta	=	16'h	c406;
44647	:douta	=	16'h	c406;
44648	:douta	=	16'h	c406;
44649	:douta	=	16'h	c425;
44650	:douta	=	16'h	c425;
44651	:douta	=	16'h	c445;
44652	:douta	=	16'h	c425;
44653	:douta	=	16'h	c425;
44654	:douta	=	16'h	c405;
44655	:douta	=	16'h	c425;
44656	:douta	=	16'h	cc25;
44657	:douta	=	16'h	c425;
44658	:douta	=	16'h	c425;
44659	:douta	=	16'h	c425;
44660	:douta	=	16'h	cc26;
44661	:douta	=	16'h	cc25;
44662	:douta	=	16'h	cc25;
44663	:douta	=	16'h	cc26;
44664	:douta	=	16'h	cc46;
44665	:douta	=	16'h	cc46;
44666	:douta	=	16'h	cc46;
44667	:douta	=	16'h	cc47;
44668	:douta	=	16'h	cc46;
44669	:douta	=	16'h	cc46;
44670	:douta	=	16'h	cc46;
44671	:douta	=	16'h	cc47;
44672	:douta	=	16'h	cc66;
44673	:douta	=	16'h	cc46;
44674	:douta	=	16'h	cc46;
44675	:douta	=	16'h	cc47;
44676	:douta	=	16'h	d467;
44677	:douta	=	16'h	cc66;
44678	:douta	=	16'h	cc66;
44679	:douta	=	16'h	cc47;
44680	:douta	=	16'h	d467;
44681	:douta	=	16'h	d467;
44682	:douta	=	16'h	d467;
44683	:douta	=	16'h	d467;
44684	:douta	=	16'h	d466;
44685	:douta	=	16'h	d467;
44686	:douta	=	16'h	d466;
44687	:douta	=	16'h	d467;
44688	:douta	=	16'h	d467;
44689	:douta	=	16'h	d467;
44690	:douta	=	16'h	d467;
44691	:douta	=	16'h	d467;
44692	:douta	=	16'h	d467;
44693	:douta	=	16'h	d467;
44694	:douta	=	16'h	d467;
44695	:douta	=	16'h	d467;
44696	:douta	=	16'h	d467;
44697	:douta	=	16'h	d467;
44698	:douta	=	16'h	d466;
44699	:douta	=	16'h	d467;
44700	:douta	=	16'h	d467;
44701	:douta	=	16'h	d467;
44702	:douta	=	16'h	d467;
44703	:douta	=	16'h	d467;
44704	:douta	=	16'h	d487;
44705	:douta	=	16'h	d486;
44706	:douta	=	16'h	ac4d;
44707	:douta	=	16'h	ac91;
44708	:douta	=	16'h	a491;
44709	:douta	=	16'h	c553;
44710	:douta	=	16'h	c573;
44711	:douta	=	16'h	c594;
44712	:douta	=	16'h	d616;
44713	:douta	=	16'h	bd74;
44714	:douta	=	16'h	c5b6;
44715	:douta	=	16'h	ad16;
44716	:douta	=	16'h	ad36;
44717	:douta	=	16'h	ad36;
44718	:douta	=	16'h	a516;
44719	:douta	=	16'h	9cd6;
44720	:douta	=	16'h	9495;
44721	:douta	=	16'h	8c94;
44722	:douta	=	16'h	73f2;
44723	:douta	=	16'h	6b91;
44724	:douta	=	16'h	8c52;
44725	:douta	=	16'h	73b1;
44726	:douta	=	16'h	7c11;
44727	:douta	=	16'h	73b1;
44728	:douta	=	16'h	73b0;
44729	:douta	=	16'h	7390;
44730	:douta	=	16'h	6b70;
44731	:douta	=	16'h	630d;
44732	:douta	=	16'h	41e7;
44733	:douta	=	16'h	39a5;
44734	:douta	=	16'h	5aa9;
44735	:douta	=	16'h	62ca;
44736	:douta	=	16'h	8bcd;
44737	:douta	=	16'h	83ac;
44738	:douta	=	16'h	8c0e;
44739	:douta	=	16'h	9c6f;
44740	:douta	=	16'h	942e;
44741	:douta	=	16'h	b4f0;
44742	:douta	=	16'h	c572;
44743	:douta	=	16'h	bd31;
44744	:douta	=	16'h	836c;
44745	:douta	=	16'h	9c2e;
44746	:douta	=	16'h	cdd4;
44747	:douta	=	16'h	cdd3;
44748	:douta	=	16'h	cdd4;
44749	:douta	=	16'h	cd92;
44750	:douta	=	16'h	c572;
44751	:douta	=	16'h	cdb4;
44752	:douta	=	16'h	d615;
44753	:douta	=	16'h	de36;
44754	:douta	=	16'h	de35;
44755	:douta	=	16'h	e656;
44756	:douta	=	16'h	d614;
44757	:douta	=	16'h	cd93;
44758	:douta	=	16'h	cd93;
44759	:douta	=	16'h	c533;
44760	:douta	=	16'h	bcf3;
44761	:douta	=	16'h	a4d3;
44762	:douta	=	16'h	8c93;
44763	:douta	=	16'h	8c74;
44764	:douta	=	16'h	9494;
44765	:douta	=	16'h	8433;
44766	:douta	=	16'h	73b1;
44767	:douta	=	16'h	6350;
44768	:douta	=	16'h	634f;
44769	:douta	=	16'h	5b0f;
44770	:douta	=	16'h	5b0f;
44771	:douta	=	16'h	4aae;
44772	:douta	=	16'h	21a8;
44773	:douta	=	16'h	62ed;
44774	:douta	=	16'h	08a5;
44775	:douta	=	16'h	10e4;
44776	:douta	=	16'h	10e4;
44777	:douta	=	16'h	1107;
44778	:douta	=	16'h	3965;
44779	:douta	=	16'h	59e5;
44780	:douta	=	16'h	5a26;
44781	:douta	=	16'h	59e6;
44782	:douta	=	16'h	51c6;
44783	:douta	=	16'h	59c6;
44784	:douta	=	16'h	51c5;
44785	:douta	=	16'h	49a5;
44786	:douta	=	16'h	49a5;
44787	:douta	=	16'h	49a6;
44788	:douta	=	16'h	49a6;
44789	:douta	=	16'h	49a5;
44790	:douta	=	16'h	49a6;
44791	:douta	=	16'h	49a6;
44792	:douta	=	16'h	4185;
44793	:douta	=	16'h	4185;
44794	:douta	=	16'h	4186;
44795	:douta	=	16'h	4166;
44796	:douta	=	16'h	4186;
44797	:douta	=	16'h	4186;
44798	:douta	=	16'h	3966;
44799	:douta	=	16'h	3986;
44800	:douta	=	16'h	ff7c;
44801	:douta	=	16'h	ffdd;
44802	:douta	=	16'h	ffdd;
44803	:douta	=	16'h	fffe;
44804	:douta	=	16'h	de15;
44805	:douta	=	16'h	e677;
44806	:douta	=	16'h	e657;
44807	:douta	=	16'h	b555;
44808	:douta	=	16'h	9453;
44809	:douta	=	16'h	bdb7;
44810	:douta	=	16'h	b576;
44811	:douta	=	16'h	bd75;
44812	:douta	=	16'h	c596;
44813	:douta	=	16'h	c595;
44814	:douta	=	16'h	bd76;
44815	:douta	=	16'h	a516;
44816	:douta	=	16'h	9495;
44817	:douta	=	16'h	8c95;
44818	:douta	=	16'h	8475;
44819	:douta	=	16'h	8c75;
44820	:douta	=	16'h	8474;
44821	:douta	=	16'h	8454;
44822	:douta	=	16'h	8455;
44823	:douta	=	16'h	8475;
44824	:douta	=	16'h	7c33;
44825	:douta	=	16'h	7c33;
44826	:douta	=	16'h	8495;
44827	:douta	=	16'h	324b;
44828	:douta	=	16'h	29c8;
44829	:douta	=	16'h	1881;
44830	:douta	=	16'h	1861;
44831	:douta	=	16'h	18a2;
44832	:douta	=	16'h	1882;
44833	:douta	=	16'h	1062;
44834	:douta	=	16'h	1061;
44835	:douta	=	16'h	1040;
44836	:douta	=	16'h	1061;
44837	:douta	=	16'h	1061;
44838	:douta	=	16'h	1861;
44839	:douta	=	16'h	20c3;
44840	:douta	=	16'h	20c3;
44841	:douta	=	16'h	2924;
44842	:douta	=	16'h	3145;
44843	:douta	=	16'h	39a6;
44844	:douta	=	16'h	39c7;
44845	:douta	=	16'h	4a28;
44846	:douta	=	16'h	5269;
44847	:douta	=	16'h	5269;
44848	:douta	=	16'h	5248;
44849	:douta	=	16'h	4a27;
44850	:douta	=	16'h	4a27;
44851	:douta	=	16'h	2967;
44852	:douta	=	16'h	2967;
44853	:douta	=	16'h	20e3;
44854	:douta	=	16'h	4123;
44855	:douta	=	16'h	3902;
44856	:douta	=	16'h	3902;
44857	:douta	=	16'h	4122;
44858	:douta	=	16'h	4142;
44859	:douta	=	16'h	4963;
44860	:douta	=	16'h	4964;
44861	:douta	=	16'h	51a4;
44862	:douta	=	16'h	51a4;
44863	:douta	=	16'h	6aea;
44864	:douta	=	16'h	834a;
44865	:douta	=	16'h	3102;
44866	:douta	=	16'h	6a04;
44867	:douta	=	16'h	61e4;
44868	:douta	=	16'h	61e4;
44869	:douta	=	16'h	6a04;
44870	:douta	=	16'h	6a24;
44871	:douta	=	16'h	7224;
44872	:douta	=	16'h	6a24;
44873	:douta	=	16'h	7244;
44874	:douta	=	16'h	7224;
44875	:douta	=	16'h	7244;
44876	:douta	=	16'h	7224;
44877	:douta	=	16'h	7a44;
44878	:douta	=	16'h	8284;
44879	:douta	=	16'h	7a63;
44880	:douta	=	16'h	8284;
44881	:douta	=	16'h	8aa4;
44882	:douta	=	16'h	8aa4;
44883	:douta	=	16'h	8ac5;
44884	:douta	=	16'h	92e5;
44885	:douta	=	16'h	9305;
44886	:douta	=	16'h	9b05;
44887	:douta	=	16'h	9b05;
44888	:douta	=	16'h	a325;
44889	:douta	=	16'h	9b25;
44890	:douta	=	16'h	ab65;
44891	:douta	=	16'h	ab65;
44892	:douta	=	16'h	ab65;
44893	:douta	=	16'h	ab65;
44894	:douta	=	16'h	b385;
44895	:douta	=	16'h	b3a5;
44896	:douta	=	16'h	b3a5;
44897	:douta	=	16'h	b3c5;
44898	:douta	=	16'h	bbc4;
44899	:douta	=	16'h	bbc5;
44900	:douta	=	16'h	bbc6;
44901	:douta	=	16'h	bbe5;
44902	:douta	=	16'h	bbc5;
44903	:douta	=	16'h	c405;
44904	:douta	=	16'h	c405;
44905	:douta	=	16'h	bbe5;
44906	:douta	=	16'h	c405;
44907	:douta	=	16'h	c405;
44908	:douta	=	16'h	c426;
44909	:douta	=	16'h	c426;
44910	:douta	=	16'h	c405;
44911	:douta	=	16'h	c405;
44912	:douta	=	16'h	c405;
44913	:douta	=	16'h	c425;
44914	:douta	=	16'h	cc26;
44915	:douta	=	16'h	c425;
44916	:douta	=	16'h	cc25;
44917	:douta	=	16'h	cc26;
44918	:douta	=	16'h	cc26;
44919	:douta	=	16'h	cc26;
44920	:douta	=	16'h	cc46;
44921	:douta	=	16'h	cc46;
44922	:douta	=	16'h	cc46;
44923	:douta	=	16'h	cc46;
44924	:douta	=	16'h	cc46;
44925	:douta	=	16'h	cc46;
44926	:douta	=	16'h	cc66;
44927	:douta	=	16'h	cc46;
44928	:douta	=	16'h	cc66;
44929	:douta	=	16'h	cc66;
44930	:douta	=	16'h	cc47;
44931	:douta	=	16'h	d467;
44932	:douta	=	16'h	d467;
44933	:douta	=	16'h	d467;
44934	:douta	=	16'h	d467;
44935	:douta	=	16'h	d466;
44936	:douta	=	16'h	cc47;
44937	:douta	=	16'h	d467;
44938	:douta	=	16'h	d466;
44939	:douta	=	16'h	d466;
44940	:douta	=	16'h	d466;
44941	:douta	=	16'h	d466;
44942	:douta	=	16'h	cc66;
44943	:douta	=	16'h	d466;
44944	:douta	=	16'h	cc66;
44945	:douta	=	16'h	d467;
44946	:douta	=	16'h	d467;
44947	:douta	=	16'h	d467;
44948	:douta	=	16'h	d467;
44949	:douta	=	16'h	d467;
44950	:douta	=	16'h	d467;
44951	:douta	=	16'h	d467;
44952	:douta	=	16'h	d467;
44953	:douta	=	16'h	d467;
44954	:douta	=	16'h	d467;
44955	:douta	=	16'h	d467;
44956	:douta	=	16'h	d467;
44957	:douta	=	16'h	d467;
44958	:douta	=	16'h	d487;
44959	:douta	=	16'h	d487;
44960	:douta	=	16'h	d467;
44961	:douta	=	16'h	d466;
44962	:douta	=	16'h	d486;
44963	:douta	=	16'h	942f;
44964	:douta	=	16'h	a4b1;
44965	:douta	=	16'h	a492;
44966	:douta	=	16'h	a493;
44967	:douta	=	16'h	a4d3;
44968	:douta	=	16'h	c596;
44969	:douta	=	16'h	c575;
44970	:douta	=	16'h	ad16;
44971	:douta	=	16'h	94b5;
44972	:douta	=	16'h	9cd5;
44973	:douta	=	16'h	8c74;
44974	:douta	=	16'h	83f2;
44975	:douta	=	16'h	7bf2;
44976	:douta	=	16'h	7bf1;
44977	:douta	=	16'h	7bd1;
44978	:douta	=	16'h	73d1;
44979	:douta	=	16'h	6bb1;
44980	:douta	=	16'h	6b70;
44981	:douta	=	16'h	8432;
44982	:douta	=	16'h	6b70;
44983	:douta	=	16'h	5acb;
44984	:douta	=	16'h	526a;
44985	:douta	=	16'h	39a6;
44986	:douta	=	16'h	41e7;
44987	:douta	=	16'h	5a8a;
44988	:douta	=	16'h	940e;
44989	:douta	=	16'h	942e;
44990	:douta	=	16'h	9c2e;
44991	:douta	=	16'h	b4d0;
44992	:douta	=	16'h	9c4e;
44993	:douta	=	16'h	bd10;
44994	:douta	=	16'h	c550;
44995	:douta	=	16'h	bd10;
44996	:douta	=	16'h	c551;
44997	:douta	=	16'h	bd31;
44998	:douta	=	16'h	c552;
44999	:douta	=	16'h	bd52;
45000	:douta	=	16'h	d5f4;
45001	:douta	=	16'h	cdd4;
45002	:douta	=	16'h	bd30;
45003	:douta	=	16'h	d635;
45004	:douta	=	16'h	de35;
45005	:douta	=	16'h	de15;
45006	:douta	=	16'h	de35;
45007	:douta	=	16'h	de35;
45008	:douta	=	16'h	d615;
45009	:douta	=	16'h	cdb4;
45010	:douta	=	16'h	cd94;
45011	:douta	=	16'h	c573;
45012	:douta	=	16'h	bd53;
45013	:douta	=	16'h	b514;
45014	:douta	=	16'h	b4f4;
45015	:douta	=	16'h	9cb4;
45016	:douta	=	16'h	9cb4;
45017	:douta	=	16'h	9cb4;
45018	:douta	=	16'h	8c73;
45019	:douta	=	16'h	8c93;
45020	:douta	=	16'h	8c74;
45021	:douta	=	16'h	8c74;
45022	:douta	=	16'h	7bf3;
45023	:douta	=	16'h	6b6f;
45024	:douta	=	16'h	5b2e;
45025	:douta	=	16'h	4acd;
45026	:douta	=	16'h	4aad;
45027	:douta	=	16'h	424b;
45028	:douta	=	16'h	39ea;
45029	:douta	=	16'h	2167;
45030	:douta	=	16'h	83f1;
45031	:douta	=	16'h	3189;
45032	:douta	=	16'h	1905;
45033	:douta	=	16'h	1905;
45034	:douta	=	16'h	1905;
45035	:douta	=	16'h	1905;
45036	:douta	=	16'h	51c5;
45037	:douta	=	16'h	59e6;
45038	:douta	=	16'h	51c6;
45039	:douta	=	16'h	51c5;
45040	:douta	=	16'h	51c6;
45041	:douta	=	16'h	51c5;
45042	:douta	=	16'h	51e6;
45043	:douta	=	16'h	49a6;
45044	:douta	=	16'h	49a6;
45045	:douta	=	16'h	49a6;
45046	:douta	=	16'h	49a6;
45047	:douta	=	16'h	49a6;
45048	:douta	=	16'h	4165;
45049	:douta	=	16'h	41a6;
45050	:douta	=	16'h	4186;
45051	:douta	=	16'h	4166;
45052	:douta	=	16'h	4166;
45053	:douta	=	16'h	3966;
45054	:douta	=	16'h	4166;
45055	:douta	=	16'h	3986;
45056	:douta	=	16'h	ff7c;
45057	:douta	=	16'h	ffdd;
45058	:douta	=	16'h	ffbd;
45059	:douta	=	16'h	ffff;
45060	:douta	=	16'h	d5d5;
45061	:douta	=	16'h	eeb8;
45062	:douta	=	16'h	d617;
45063	:douta	=	16'h	ad15;
45064	:douta	=	16'h	9c73;
45065	:douta	=	16'h	bdb7;
45066	:douta	=	16'h	bd96;
45067	:douta	=	16'h	bd75;
45068	:douta	=	16'h	c5b6;
45069	:douta	=	16'h	c595;
45070	:douta	=	16'h	b556;
45071	:douta	=	16'h	9cb5;
45072	:douta	=	16'h	94b5;
45073	:douta	=	16'h	8c74;
45074	:douta	=	16'h	8c75;
45075	:douta	=	16'h	8475;
45076	:douta	=	16'h	8454;
45077	:douta	=	16'h	8454;
45078	:douta	=	16'h	8475;
45079	:douta	=	16'h	7c54;
45080	:douta	=	16'h	7c33;
45081	:douta	=	16'h	8454;
45082	:douta	=	16'h	4a8b;
45083	:douta	=	16'h	1062;
45084	:douta	=	16'h	3a6a;
45085	:douta	=	16'h	31c9;
45086	:douta	=	16'h	2126;
45087	:douta	=	16'h	1882;
45088	:douta	=	16'h	1841;
45089	:douta	=	16'h	1882;
45090	:douta	=	16'h	18a3;
45091	:douta	=	16'h	18c3;
45092	:douta	=	16'h	2124;
45093	:douta	=	16'h	2124;
45094	:douta	=	16'h	2965;
45095	:douta	=	16'h	29a6;
45096	:douta	=	16'h	31a7;
45097	:douta	=	16'h	39e7;
45098	:douta	=	16'h	39e8;
45099	:douta	=	16'h	39c7;
45100	:douta	=	16'h	39a6;
45101	:douta	=	16'h	3966;
45102	:douta	=	16'h	3965;
45103	:douta	=	16'h	3144;
45104	:douta	=	16'h	3103;
45105	:douta	=	16'h	28e2;
45106	:douta	=	16'h	30e2;
45107	:douta	=	16'h	31a7;
45108	:douta	=	16'h	2967;
45109	:douta	=	16'h	28e3;
45110	:douta	=	16'h	3903;
45111	:douta	=	16'h	4123;
45112	:douta	=	16'h	4143;
45113	:douta	=	16'h	4123;
45114	:douta	=	16'h	4963;
45115	:douta	=	16'h	5184;
45116	:douta	=	16'h	49a4;
45117	:douta	=	16'h	51a4;
45118	:douta	=	16'h	51a3;
45119	:douta	=	16'h	734c;
45120	:douta	=	16'h	7b08;
45121	:douta	=	16'h	4122;
45122	:douta	=	16'h	6a03;
45123	:douta	=	16'h	61e4;
45124	:douta	=	16'h	69e4;
45125	:douta	=	16'h	6a24;
45126	:douta	=	16'h	6a04;
45127	:douta	=	16'h	7224;
45128	:douta	=	16'h	7224;
45129	:douta	=	16'h	7244;
45130	:douta	=	16'h	7224;
45131	:douta	=	16'h	7224;
45132	:douta	=	16'h	7244;
45133	:douta	=	16'h	7a44;
45134	:douta	=	16'h	7a64;
45135	:douta	=	16'h	82a4;
45136	:douta	=	16'h	8284;
45137	:douta	=	16'h	8aa4;
45138	:douta	=	16'h	8aa4;
45139	:douta	=	16'h	8ac4;
45140	:douta	=	16'h	92e4;
45141	:douta	=	16'h	92e4;
45142	:douta	=	16'h	9b26;
45143	:douta	=	16'h	9b25;
45144	:douta	=	16'h	9b25;
45145	:douta	=	16'h	9b25;
45146	:douta	=	16'h	a365;
45147	:douta	=	16'h	ab65;
45148	:douta	=	16'h	ab65;
45149	:douta	=	16'h	ab85;
45150	:douta	=	16'h	b385;
45151	:douta	=	16'h	b385;
45152	:douta	=	16'h	b3c5;
45153	:douta	=	16'h	b3a5;
45154	:douta	=	16'h	bbc5;
45155	:douta	=	16'h	b3c5;
45156	:douta	=	16'h	bbc6;
45157	:douta	=	16'h	bbe6;
45158	:douta	=	16'h	bbe5;
45159	:douta	=	16'h	bbe5;
45160	:douta	=	16'h	bbe5;
45161	:douta	=	16'h	c405;
45162	:douta	=	16'h	c405;
45163	:douta	=	16'h	c405;
45164	:douta	=	16'h	c426;
45165	:douta	=	16'h	c406;
45166	:douta	=	16'h	c425;
45167	:douta	=	16'h	c425;
45168	:douta	=	16'h	c425;
45169	:douta	=	16'h	c425;
45170	:douta	=	16'h	c425;
45171	:douta	=	16'h	c425;
45172	:douta	=	16'h	cc25;
45173	:douta	=	16'h	cc25;
45174	:douta	=	16'h	cc46;
45175	:douta	=	16'h	cc46;
45176	:douta	=	16'h	cc46;
45177	:douta	=	16'h	cc46;
45178	:douta	=	16'h	cc46;
45179	:douta	=	16'h	cc46;
45180	:douta	=	16'h	cc47;
45181	:douta	=	16'h	cc45;
45182	:douta	=	16'h	cc66;
45183	:douta	=	16'h	cc46;
45184	:douta	=	16'h	cc66;
45185	:douta	=	16'h	cc66;
45186	:douta	=	16'h	cc47;
45187	:douta	=	16'h	cc46;
45188	:douta	=	16'h	cc47;
45189	:douta	=	16'h	d467;
45190	:douta	=	16'h	d467;
45191	:douta	=	16'h	cc66;
45192	:douta	=	16'h	d467;
45193	:douta	=	16'h	d467;
45194	:douta	=	16'h	cc66;
45195	:douta	=	16'h	d466;
45196	:douta	=	16'h	d467;
45197	:douta	=	16'h	d466;
45198	:douta	=	16'h	d466;
45199	:douta	=	16'h	d466;
45200	:douta	=	16'h	cc66;
45201	:douta	=	16'h	d467;
45202	:douta	=	16'h	d467;
45203	:douta	=	16'h	d487;
45204	:douta	=	16'h	d467;
45205	:douta	=	16'h	d467;
45206	:douta	=	16'h	d467;
45207	:douta	=	16'h	d467;
45208	:douta	=	16'h	d467;
45209	:douta	=	16'h	d467;
45210	:douta	=	16'h	d467;
45211	:douta	=	16'h	d467;
45212	:douta	=	16'h	d467;
45213	:douta	=	16'h	d487;
45214	:douta	=	16'h	d487;
45215	:douta	=	16'h	d466;
45216	:douta	=	16'h	d487;
45217	:douta	=	16'h	d466;
45218	:douta	=	16'h	d487;
45219	:douta	=	16'h	9c0d;
45220	:douta	=	16'h	9430;
45221	:douta	=	16'h	a4d2;
45222	:douta	=	16'h	9c72;
45223	:douta	=	16'h	9c72;
45224	:douta	=	16'h	b536;
45225	:douta	=	16'h	b515;
45226	:douta	=	16'h	a4d5;
45227	:douta	=	16'h	9495;
45228	:douta	=	16'h	8c74;
45229	:douta	=	16'h	7bf2;
45230	:douta	=	16'h	7390;
45231	:douta	=	16'h	73d1;
45232	:douta	=	16'h	73d0;
45233	:douta	=	16'h	73b1;
45234	:douta	=	16'h	73b0;
45235	:douta	=	16'h	6b90;
45236	:douta	=	16'h	6b90;
45237	:douta	=	16'h	7390;
45238	:douta	=	16'h	634e;
45239	:douta	=	16'h	1881;
45240	:douta	=	16'h	3124;
45241	:douta	=	16'h	6aeb;
45242	:douta	=	16'h	7b6e;
45243	:douta	=	16'h	942f;
45244	:douta	=	16'h	a46e;
45245	:douta	=	16'h	9c2e;
45246	:douta	=	16'h	b531;
45247	:douta	=	16'h	c571;
45248	:douta	=	16'h	b4ef;
45249	:douta	=	16'h	c551;
45250	:douta	=	16'h	cd92;
45251	:douta	=	16'h	c531;
45252	:douta	=	16'h	d5b3;
45253	:douta	=	16'h	c593;
45254	:douta	=	16'h	c573;
45255	:douta	=	16'h	c573;
45256	:douta	=	16'h	de36;
45257	:douta	=	16'h	de36;
45258	:douta	=	16'h	cdd4;
45259	:douta	=	16'h	d616;
45260	:douta	=	16'h	cdb4;
45261	:douta	=	16'h	de15;
45262	:douta	=	16'h	de15;
45263	:douta	=	16'h	cdd4;
45264	:douta	=	16'h	de35;
45265	:douta	=	16'h	d615;
45266	:douta	=	16'h	d5b4;
45267	:douta	=	16'h	c554;
45268	:douta	=	16'h	b514;
45269	:douta	=	16'h	a4d4;
45270	:douta	=	16'h	a4d5;
45271	:douta	=	16'h	9494;
45272	:douta	=	16'h	9c94;
45273	:douta	=	16'h	9cb4;
45274	:douta	=	16'h	9494;
45275	:douta	=	16'h	8c93;
45276	:douta	=	16'h	8c74;
45277	:douta	=	16'h	8c53;
45278	:douta	=	16'h	7bf3;
45279	:douta	=	16'h	6b91;
45280	:douta	=	16'h	634f;
45281	:douta	=	16'h	52ce;
45282	:douta	=	16'h	424c;
45283	:douta	=	16'h	31a8;
45284	:douta	=	16'h	39ea;
45285	:douta	=	16'h	29a9;
45286	:douta	=	16'h	9c92;
45287	:douta	=	16'h	424b;
45288	:douta	=	16'h	2189;
45289	:douta	=	16'h	18e5;
45290	:douta	=	16'h	1905;
45291	:douta	=	16'h	1926;
45292	:douta	=	16'h	41a6;
45293	:douta	=	16'h	51c5;
45294	:douta	=	16'h	51c6;
45295	:douta	=	16'h	51c6;
45296	:douta	=	16'h	51c6;
45297	:douta	=	16'h	51c6;
45298	:douta	=	16'h	51c5;
45299	:douta	=	16'h	49a6;
45300	:douta	=	16'h	49a6;
45301	:douta	=	16'h	49a6;
45302	:douta	=	16'h	49a6;
45303	:douta	=	16'h	4185;
45304	:douta	=	16'h	4185;
45305	:douta	=	16'h	4185;
45306	:douta	=	16'h	4166;
45307	:douta	=	16'h	4186;
45308	:douta	=	16'h	3945;
45309	:douta	=	16'h	4166;
45310	:douta	=	16'h	4166;
45311	:douta	=	16'h	4186;
45312	:douta	=	16'h	ff9c;
45313	:douta	=	16'h	ff9d;
45314	:douta	=	16'h	ff9d;
45315	:douta	=	16'h	ffbd;
45316	:douta	=	16'h	de37;
45317	:douta	=	16'h	eeb8;
45318	:douta	=	16'h	bd96;
45319	:douta	=	16'h	a4f4;
45320	:douta	=	16'h	9c93;
45321	:douta	=	16'h	bd96;
45322	:douta	=	16'h	b535;
45323	:douta	=	16'h	c5b5;
45324	:douta	=	16'h	bd95;
45325	:douta	=	16'h	bd55;
45326	:douta	=	16'h	a516;
45327	:douta	=	16'h	8c53;
45328	:douta	=	16'h	8cb5;
45329	:douta	=	16'h	8454;
45330	:douta	=	16'h	8c95;
45331	:douta	=	16'h	8c75;
45332	:douta	=	16'h	8c75;
45333	:douta	=	16'h	8474;
45334	:douta	=	16'h	8474;
45335	:douta	=	16'h	7bf3;
45336	:douta	=	16'h	8c74;
45337	:douta	=	16'h	94f7;
45338	:douta	=	16'h	0820;
45339	:douta	=	16'h	18a3;
45340	:douta	=	16'h	18a2;
45341	:douta	=	16'h	18e3;
45342	:douta	=	16'h	2966;
45343	:douta	=	16'h	29a8;
45344	:douta	=	16'h	2147;
45345	:douta	=	16'h	2946;
45346	:douta	=	16'h	2124;
45347	:douta	=	16'h	1904;
45348	:douta	=	16'h	18e3;
45349	:douta	=	16'h	20e3;
45350	:douta	=	16'h	2082;
45351	:douta	=	16'h	2082;
45352	:douta	=	16'h	2082;
45353	:douta	=	16'h	1881;
45354	:douta	=	16'h	1881;
45355	:douta	=	16'h	2082;
45356	:douta	=	16'h	20a1;
45357	:douta	=	16'h	20c2;
45358	:douta	=	16'h	28c2;
45359	:douta	=	16'h	28e2;
45360	:douta	=	16'h	30e3;
45361	:douta	=	16'h	30e3;
45362	:douta	=	16'h	3103;
45363	:douta	=	16'h	29a8;
45364	:douta	=	16'h	2126;
45365	:douta	=	16'h	30e3;
45366	:douta	=	16'h	4143;
45367	:douta	=	16'h	4143;
45368	:douta	=	16'h	4963;
45369	:douta	=	16'h	4963;
45370	:douta	=	16'h	4984;
45371	:douta	=	16'h	4964;
45372	:douta	=	16'h	51a4;
45373	:douta	=	16'h	51a4;
45374	:douta	=	16'h	5183;
45375	:douta	=	16'h	83ef;
45376	:douta	=	16'h	6a44;
45377	:douta	=	16'h	59a3;
45378	:douta	=	16'h	61e4;
45379	:douta	=	16'h	69e4;
45380	:douta	=	16'h	6a04;
45381	:douta	=	16'h	7224;
45382	:douta	=	16'h	7224;
45383	:douta	=	16'h	7224;
45384	:douta	=	16'h	7244;
45385	:douta	=	16'h	7244;
45386	:douta	=	16'h	7224;
45387	:douta	=	16'h	7244;
45388	:douta	=	16'h	7224;
45389	:douta	=	16'h	7224;
45390	:douta	=	16'h	8284;
45391	:douta	=	16'h	8285;
45392	:douta	=	16'h	8284;
45393	:douta	=	16'h	8aa4;
45394	:douta	=	16'h	8aa4;
45395	:douta	=	16'h	92e5;
45396	:douta	=	16'h	9305;
45397	:douta	=	16'h	9305;
45398	:douta	=	16'h	9b05;
45399	:douta	=	16'h	9b05;
45400	:douta	=	16'h	9b25;
45401	:douta	=	16'h	a345;
45402	:douta	=	16'h	a365;
45403	:douta	=	16'h	ab64;
45404	:douta	=	16'h	ab65;
45405	:douta	=	16'h	b385;
45406	:douta	=	16'h	ab85;
45407	:douta	=	16'h	b3a5;
45408	:douta	=	16'h	b3a5;
45409	:douta	=	16'h	b3c5;
45410	:douta	=	16'h	bbc5;
45411	:douta	=	16'h	bbe6;
45412	:douta	=	16'h	bbc6;
45413	:douta	=	16'h	bbc6;
45414	:douta	=	16'h	bbe5;
45415	:douta	=	16'h	bbe5;
45416	:douta	=	16'h	c406;
45417	:douta	=	16'h	c405;
45418	:douta	=	16'h	c405;
45419	:douta	=	16'h	c406;
45420	:douta	=	16'h	c426;
45421	:douta	=	16'h	c406;
45422	:douta	=	16'h	c405;
45423	:douta	=	16'h	c425;
45424	:douta	=	16'h	c425;
45425	:douta	=	16'h	c425;
45426	:douta	=	16'h	cc26;
45427	:douta	=	16'h	c425;
45428	:douta	=	16'h	cc26;
45429	:douta	=	16'h	cc26;
45430	:douta	=	16'h	cc46;
45431	:douta	=	16'h	cc46;
45432	:douta	=	16'h	cc46;
45433	:douta	=	16'h	cc46;
45434	:douta	=	16'h	cc46;
45435	:douta	=	16'h	cc46;
45436	:douta	=	16'h	cc46;
45437	:douta	=	16'h	d467;
45438	:douta	=	16'h	cc47;
45439	:douta	=	16'h	d467;
45440	:douta	=	16'h	d467;
45441	:douta	=	16'h	cc46;
45442	:douta	=	16'h	d467;
45443	:douta	=	16'h	d467;
45444	:douta	=	16'h	d467;
45445	:douta	=	16'h	cc46;
45446	:douta	=	16'h	d466;
45447	:douta	=	16'h	d467;
45448	:douta	=	16'h	d467;
45449	:douta	=	16'h	d467;
45450	:douta	=	16'h	d467;
45451	:douta	=	16'h	d467;
45452	:douta	=	16'h	d466;
45453	:douta	=	16'h	d466;
45454	:douta	=	16'h	d467;
45455	:douta	=	16'h	d467;
45456	:douta	=	16'h	d467;
45457	:douta	=	16'h	d467;
45458	:douta	=	16'h	d467;
45459	:douta	=	16'h	d467;
45460	:douta	=	16'h	d467;
45461	:douta	=	16'h	d467;
45462	:douta	=	16'h	d467;
45463	:douta	=	16'h	d467;
45464	:douta	=	16'h	d487;
45465	:douta	=	16'h	d467;
45466	:douta	=	16'h	d467;
45467	:douta	=	16'h	d467;
45468	:douta	=	16'h	d467;
45469	:douta	=	16'h	d487;
45470	:douta	=	16'h	d467;
45471	:douta	=	16'h	d487;
45472	:douta	=	16'h	cc67;
45473	:douta	=	16'h	cc87;
45474	:douta	=	16'h	d467;
45475	:douta	=	16'h	cd6f;
45476	:douta	=	16'h	9c90;
45477	:douta	=	16'h	acd3;
45478	:douta	=	16'h	8c10;
45479	:douta	=	16'h	9452;
45480	:douta	=	16'h	9c73;
45481	:douta	=	16'h	9473;
45482	:douta	=	16'h	7bf1;
45483	:douta	=	16'h	83f1;
45484	:douta	=	16'h	8432;
45485	:douta	=	16'h	7bd0;
45486	:douta	=	16'h	736f;
45487	:douta	=	16'h	6b4f;
45488	:douta	=	16'h	632f;
45489	:douta	=	16'h	6b4f;
45490	:douta	=	16'h	6b4f;
45491	:douta	=	16'h	5acd;
45492	:douta	=	16'h	39a5;
45493	:douta	=	16'h	5a68;
45494	:douta	=	16'h	732b;
45495	:douta	=	16'h	8bcd;
45496	:douta	=	16'h	942e;
45497	:douta	=	16'h	a4b0;
45498	:douta	=	16'h	acf1;
45499	:douta	=	16'h	c573;
45500	:douta	=	16'h	b511;
45501	:douta	=	16'h	c572;
45502	:douta	=	16'h	cdb3;
45503	:douta	=	16'h	c573;
45504	:douta	=	16'h	cd93;
45505	:douta	=	16'h	ddf4;
45506	:douta	=	16'h	d5f4;
45507	:douta	=	16'h	d5d3;
45508	:douta	=	16'h	de15;
45509	:douta	=	16'h	de35;
45510	:douta	=	16'h	c574;
45511	:douta	=	16'h	c5b4;
45512	:douta	=	16'h	e676;
45513	:douta	=	16'h	c594;
45514	:douta	=	16'h	cdb4;
45515	:douta	=	16'h	cdf4;
45516	:douta	=	16'h	cdf4;
45517	:douta	=	16'h	c5b4;
45518	:douta	=	16'h	c594;
45519	:douta	=	16'h	cdb4;
45520	:douta	=	16'h	cd94;
45521	:douta	=	16'h	c574;
45522	:douta	=	16'h	b513;
45523	:douta	=	16'h	b514;
45524	:douta	=	16'h	acf4;
45525	:douta	=	16'h	a4f4;
45526	:douta	=	16'h	9cd3;
45527	:douta	=	16'h	94b4;
45528	:douta	=	16'h	9494;
45529	:douta	=	16'h	8c93;
45530	:douta	=	16'h	8432;
45531	:douta	=	16'h	8412;
45532	:douta	=	16'h	7bf2;
45533	:douta	=	16'h	73b1;
45534	:douta	=	16'h	7391;
45535	:douta	=	16'h	73d1;
45536	:douta	=	16'h	73b1;
45537	:douta	=	16'h	6b90;
45538	:douta	=	16'h	6b91;
45539	:douta	=	16'h	632d;
45540	:douta	=	16'h	18c4;
45541	:douta	=	16'h	18a3;
45542	:douta	=	16'h	5aab;
45543	:douta	=	16'h	732e;
45544	:douta	=	16'h	2147;
45545	:douta	=	16'h	29c9;
45546	:douta	=	16'h	2127;
45547	:douta	=	16'h	18e5;
45548	:douta	=	16'h	1906;
45549	:douta	=	16'h	61e6;
45550	:douta	=	16'h	51e6;
45551	:douta	=	16'h	59e6;
45552	:douta	=	16'h	51e6;
45553	:douta	=	16'h	51c6;
45554	:douta	=	16'h	51c6;
45555	:douta	=	16'h	49a6;
45556	:douta	=	16'h	49a6;
45557	:douta	=	16'h	49a5;
45558	:douta	=	16'h	4986;
45559	:douta	=	16'h	4185;
45560	:douta	=	16'h	41a6;
45561	:douta	=	16'h	4185;
45562	:douta	=	16'h	4166;
45563	:douta	=	16'h	4186;
45564	:douta	=	16'h	4166;
45565	:douta	=	16'h	3966;
45566	:douta	=	16'h	4186;
45567	:douta	=	16'h	3966;
45568	:douta	=	16'h	ff9c;
45569	:douta	=	16'h	ffbd;
45570	:douta	=	16'h	ffbd;
45571	:douta	=	16'h	f71a;
45572	:douta	=	16'h	e698;
45573	:douta	=	16'h	ee98;
45574	:douta	=	16'h	bd96;
45575	:douta	=	16'h	a4b4;
45576	:douta	=	16'h	b535;
45577	:douta	=	16'h	bd76;
45578	:douta	=	16'h	b514;
45579	:douta	=	16'h	cdb5;
45580	:douta	=	16'h	c5b6;
45581	:douta	=	16'h	bd76;
45582	:douta	=	16'h	94b4;
45583	:douta	=	16'h	8433;
45584	:douta	=	16'h	8c74;
45585	:douta	=	16'h	8454;
45586	:douta	=	16'h	8474;
45587	:douta	=	16'h	8454;
45588	:douta	=	16'h	8474;
45589	:douta	=	16'h	8434;
45590	:douta	=	16'h	7413;
45591	:douta	=	16'h	7c13;
45592	:douta	=	16'h	9d17;
45593	:douta	=	16'h	7412;
45594	:douta	=	16'h	18a2;
45595	:douta	=	16'h	20a2;
45596	:douta	=	16'h	18c3;
45597	:douta	=	16'h	20a2;
45598	:douta	=	16'h	1882;
45599	:douta	=	16'h	18a3;
45600	:douta	=	16'h	1883;
45601	:douta	=	16'h	18a2;
45602	:douta	=	16'h	1861;
45603	:douta	=	16'h	1882;
45604	:douta	=	16'h	1881;
45605	:douta	=	16'h	1881;
45606	:douta	=	16'h	1881;
45607	:douta	=	16'h	2082;
45608	:douta	=	16'h	2082;
45609	:douta	=	16'h	20a2;
45610	:douta	=	16'h	20a2;
45611	:douta	=	16'h	20a2;
45612	:douta	=	16'h	20a2;
45613	:douta	=	16'h	28e2;
45614	:douta	=	16'h	28c2;
45615	:douta	=	16'h	28c2;
45616	:douta	=	16'h	28e2;
45617	:douta	=	16'h	30e2;
45618	:douta	=	16'h	2903;
45619	:douta	=	16'h	2988;
45620	:douta	=	16'h	1905;
45621	:douta	=	16'h	3103;
45622	:douta	=	16'h	4143;
45623	:douta	=	16'h	4143;
45624	:douta	=	16'h	4143;
45625	:douta	=	16'h	4963;
45626	:douta	=	16'h	4964;
45627	:douta	=	16'h	5184;
45628	:douta	=	16'h	51a4;
45629	:douta	=	16'h	51a4;
45630	:douta	=	16'h	5163;
45631	:douta	=	16'h	8c91;
45632	:douta	=	16'h	61c4;
45633	:douta	=	16'h	69e4;
45634	:douta	=	16'h	51a4;
45635	:douta	=	16'h	6a04;
45636	:douta	=	16'h	69e4;
45637	:douta	=	16'h	6a04;
45638	:douta	=	16'h	6a04;
45639	:douta	=	16'h	7224;
45640	:douta	=	16'h	7244;
45641	:douta	=	16'h	7a44;
45642	:douta	=	16'h	7224;
45643	:douta	=	16'h	7224;
45644	:douta	=	16'h	7a44;
45645	:douta	=	16'h	7a44;
45646	:douta	=	16'h	7a64;
45647	:douta	=	16'h	8285;
45648	:douta	=	16'h	82a4;
45649	:douta	=	16'h	8ac5;
45650	:douta	=	16'h	8ac5;
45651	:douta	=	16'h	8ae4;
45652	:douta	=	16'h	9304;
45653	:douta	=	16'h	9305;
45654	:douta	=	16'h	9b05;
45655	:douta	=	16'h	9b25;
45656	:douta	=	16'h	a345;
45657	:douta	=	16'h	a345;
45658	:douta	=	16'h	ab45;
45659	:douta	=	16'h	ab65;
45660	:douta	=	16'h	ab65;
45661	:douta	=	16'h	b385;
45662	:douta	=	16'h	b385;
45663	:douta	=	16'h	b3a5;
45664	:douta	=	16'h	b3a5;
45665	:douta	=	16'h	b3c6;
45666	:douta	=	16'h	bbc5;
45667	:douta	=	16'h	bbc5;
45668	:douta	=	16'h	bbc6;
45669	:douta	=	16'h	bbe5;
45670	:douta	=	16'h	bbe5;
45671	:douta	=	16'h	bc06;
45672	:douta	=	16'h	bc06;
45673	:douta	=	16'h	c3e5;
45674	:douta	=	16'h	c405;
45675	:douta	=	16'h	c406;
45676	:douta	=	16'h	c426;
45677	:douta	=	16'h	c405;
45678	:douta	=	16'h	c405;
45679	:douta	=	16'h	c425;
45680	:douta	=	16'h	c425;
45681	:douta	=	16'h	c425;
45682	:douta	=	16'h	cc26;
45683	:douta	=	16'h	cc26;
45684	:douta	=	16'h	cc25;
45685	:douta	=	16'h	cc26;
45686	:douta	=	16'h	cc46;
45687	:douta	=	16'h	cc46;
45688	:douta	=	16'h	cc46;
45689	:douta	=	16'h	cc46;
45690	:douta	=	16'h	cc47;
45691	:douta	=	16'h	cc46;
45692	:douta	=	16'h	cc46;
45693	:douta	=	16'h	cc46;
45694	:douta	=	16'h	cc46;
45695	:douta	=	16'h	cc46;
45696	:douta	=	16'h	cc47;
45697	:douta	=	16'h	cc47;
45698	:douta	=	16'h	d467;
45699	:douta	=	16'h	cc47;
45700	:douta	=	16'h	d467;
45701	:douta	=	16'h	cc66;
45702	:douta	=	16'h	cc66;
45703	:douta	=	16'h	d467;
45704	:douta	=	16'h	d467;
45705	:douta	=	16'h	d467;
45706	:douta	=	16'h	cc47;
45707	:douta	=	16'h	d466;
45708	:douta	=	16'h	cc66;
45709	:douta	=	16'h	d466;
45710	:douta	=	16'h	d467;
45711	:douta	=	16'h	d467;
45712	:douta	=	16'h	d467;
45713	:douta	=	16'h	d468;
45714	:douta	=	16'h	d467;
45715	:douta	=	16'h	d467;
45716	:douta	=	16'h	d467;
45717	:douta	=	16'h	d467;
45718	:douta	=	16'h	d487;
45719	:douta	=	16'h	d467;
45720	:douta	=	16'h	d467;
45721	:douta	=	16'h	d467;
45722	:douta	=	16'h	d467;
45723	:douta	=	16'h	d467;
45724	:douta	=	16'h	d467;
45725	:douta	=	16'h	d467;
45726	:douta	=	16'h	d487;
45727	:douta	=	16'h	d468;
45728	:douta	=	16'h	d488;
45729	:douta	=	16'h	d467;
45730	:douta	=	16'h	d468;
45731	:douta	=	16'h	bd0e;
45732	:douta	=	16'h	c614;
45733	:douta	=	16'h	940f;
45734	:douta	=	16'h	9430;
45735	:douta	=	16'h	9451;
45736	:douta	=	16'h	9452;
45737	:douta	=	16'h	8c32;
45738	:douta	=	16'h	7bb0;
45739	:douta	=	16'h	7bd0;
45740	:douta	=	16'h	736f;
45741	:douta	=	16'h	83f1;
45742	:douta	=	16'h	6b4e;
45743	:douta	=	16'h	630e;
45744	:douta	=	16'h	632e;
45745	:douta	=	16'h	630d;
45746	:douta	=	16'h	41a6;
45747	:douta	=	16'h	3124;
45748	:douta	=	16'h	940e;
45749	:douta	=	16'h	a4b0;
45750	:douta	=	16'h	732a;
45751	:douta	=	16'h	9c4f;
45752	:douta	=	16'h	acaf;
45753	:douta	=	16'h	bd51;
45754	:douta	=	16'h	bd72;
45755	:douta	=	16'h	b531;
45756	:douta	=	16'h	c593;
45757	:douta	=	16'h	de15;
45758	:douta	=	16'h	d5f4;
45759	:douta	=	16'h	cdd3;
45760	:douta	=	16'h	d5f3;
45761	:douta	=	16'h	de15;
45762	:douta	=	16'h	d5f4;
45763	:douta	=	16'h	de15;
45764	:douta	=	16'h	de36;
45765	:douta	=	16'h	e676;
45766	:douta	=	16'h	b513;
45767	:douta	=	16'h	c5b4;
45768	:douta	=	16'h	e657;
45769	:douta	=	16'h	c575;
45770	:douta	=	16'h	bd34;
45771	:douta	=	16'h	b534;
45772	:douta	=	16'h	c575;
45773	:douta	=	16'h	cdd5;
45774	:douta	=	16'h	c574;
45775	:douta	=	16'h	b534;
45776	:douta	=	16'h	bd54;
45777	:douta	=	16'h	bd34;
45778	:douta	=	16'h	acf4;
45779	:douta	=	16'h	a4d4;
45780	:douta	=	16'h	9cb4;
45781	:douta	=	16'h	9cb4;
45782	:douta	=	16'h	9494;
45783	:douta	=	16'h	8c73;
45784	:douta	=	16'h	8c53;
45785	:douta	=	16'h	8c53;
45786	:douta	=	16'h	7bf2;
45787	:douta	=	16'h	73b1;
45788	:douta	=	16'h	73b1;
45789	:douta	=	16'h	738f;
45790	:douta	=	16'h	62cc;
45791	:douta	=	16'h	41c6;
45792	:douta	=	16'h	3144;
45793	:douta	=	16'h	3965;
45794	:douta	=	16'h	3985;
45795	:douta	=	16'h	8369;
45796	:douta	=	16'h	4208;
45797	:douta	=	16'h	2147;
45798	:douta	=	16'h	426c;
45799	:douta	=	16'h	734e;
45800	:douta	=	16'h	18e5;
45801	:douta	=	16'h	29ca;
45802	:douta	=	16'h	2189;
45803	:douta	=	16'h	18e5;
45804	:douta	=	16'h	1907;
45805	:douta	=	16'h	6206;
45806	:douta	=	16'h	51e5;
45807	:douta	=	16'h	59e6;
45808	:douta	=	16'h	51c5;
45809	:douta	=	16'h	49c6;
45810	:douta	=	16'h	49c6;
45811	:douta	=	16'h	49a6;
45812	:douta	=	16'h	49a6;
45813	:douta	=	16'h	49a5;
45814	:douta	=	16'h	4185;
45815	:douta	=	16'h	49a6;
45816	:douta	=	16'h	4185;
45817	:douta	=	16'h	4185;
45818	:douta	=	16'h	4166;
45819	:douta	=	16'h	4166;
45820	:douta	=	16'h	4166;
45821	:douta	=	16'h	3966;
45822	:douta	=	16'h	3966;
45823	:douta	=	16'h	3966;
45824	:douta	=	16'h	ffbd;
45825	:douta	=	16'h	ffbd;
45826	:douta	=	16'h	ffdd;
45827	:douta	=	16'h	de77;
45828	:douta	=	16'h	e677;
45829	:douta	=	16'h	e697;
45830	:douta	=	16'h	ad14;
45831	:douta	=	16'h	a4b4;
45832	:douta	=	16'h	b554;
45833	:douta	=	16'h	b535;
45834	:douta	=	16'h	c595;
45835	:douta	=	16'h	c595;
45836	:douta	=	16'h	bd76;
45837	:douta	=	16'h	bd76;
45838	:douta	=	16'h	8453;
45839	:douta	=	16'h	8c74;
45840	:douta	=	16'h	8c94;
45841	:douta	=	16'h	8c74;
45842	:douta	=	16'h	8474;
45843	:douta	=	16'h	8454;
45844	:douta	=	16'h	8474;
45845	:douta	=	16'h	73f3;
45846	:douta	=	16'h	7c13;
45847	:douta	=	16'h	8454;
45848	:douta	=	16'h	8cb6;
45849	:douta	=	16'h	2145;
45850	:douta	=	16'h	20e3;
45851	:douta	=	16'h	18c3;
45852	:douta	=	16'h	18c3;
45853	:douta	=	16'h	18a3;
45854	:douta	=	16'h	20c3;
45855	:douta	=	16'h	1082;
45856	:douta	=	16'h	1882;
45857	:douta	=	16'h	1882;
45858	:douta	=	16'h	1882;
45859	:douta	=	16'h	1882;
45860	:douta	=	16'h	1881;
45861	:douta	=	16'h	1881;
45862	:douta	=	16'h	20a2;
45863	:douta	=	16'h	20a2;
45864	:douta	=	16'h	20a2;
45865	:douta	=	16'h	20a2;
45866	:douta	=	16'h	2082;
45867	:douta	=	16'h	20a2;
45868	:douta	=	16'h	20c2;
45869	:douta	=	16'h	20c2;
45870	:douta	=	16'h	28e3;
45871	:douta	=	16'h	28e2;
45872	:douta	=	16'h	30e3;
45873	:douta	=	16'h	30e2;
45874	:douta	=	16'h	3125;
45875	:douta	=	16'h	2988;
45876	:douta	=	16'h	18e5;
45877	:douta	=	16'h	4123;
45878	:douta	=	16'h	4143;
45879	:douta	=	16'h	4143;
45880	:douta	=	16'h	4963;
45881	:douta	=	16'h	4963;
45882	:douta	=	16'h	4963;
45883	:douta	=	16'h	51a4;
45884	:douta	=	16'h	51a4;
45885	:douta	=	16'h	59a4;
45886	:douta	=	16'h	5183;
45887	:douta	=	16'h	9d13;
45888	:douta	=	16'h	5983;
45889	:douta	=	16'h	6a04;
45890	:douta	=	16'h	4964;
45891	:douta	=	16'h	7224;
45892	:douta	=	16'h	7204;
45893	:douta	=	16'h	7224;
45894	:douta	=	16'h	7224;
45895	:douta	=	16'h	7244;
45896	:douta	=	16'h	7244;
45897	:douta	=	16'h	7244;
45898	:douta	=	16'h	7224;
45899	:douta	=	16'h	7224;
45900	:douta	=	16'h	7244;
45901	:douta	=	16'h	7a44;
45902	:douta	=	16'h	8284;
45903	:douta	=	16'h	8284;
45904	:douta	=	16'h	8283;
45905	:douta	=	16'h	8ac5;
45906	:douta	=	16'h	8ac5;
45907	:douta	=	16'h	92c4;
45908	:douta	=	16'h	9305;
45909	:douta	=	16'h	9304;
45910	:douta	=	16'h	9b05;
45911	:douta	=	16'h	a325;
45912	:douta	=	16'h	a325;
45913	:douta	=	16'h	a345;
45914	:douta	=	16'h	ab45;
45915	:douta	=	16'h	ab85;
45916	:douta	=	16'h	ab65;
45917	:douta	=	16'h	b385;
45918	:douta	=	16'h	b385;
45919	:douta	=	16'h	b385;
45920	:douta	=	16'h	b3c5;
45921	:douta	=	16'h	b3c5;
45922	:douta	=	16'h	bbe6;
45923	:douta	=	16'h	bbe5;
45924	:douta	=	16'h	bbe5;
45925	:douta	=	16'h	bbe5;
45926	:douta	=	16'h	bbe5;
45927	:douta	=	16'h	bc06;
45928	:douta	=	16'h	bbe5;
45929	:douta	=	16'h	c406;
45930	:douta	=	16'h	c405;
45931	:douta	=	16'h	c426;
45932	:douta	=	16'h	c426;
45933	:douta	=	16'h	c426;
45934	:douta	=	16'h	c406;
45935	:douta	=	16'h	c425;
45936	:douta	=	16'h	c425;
45937	:douta	=	16'h	c425;
45938	:douta	=	16'h	c425;
45939	:douta	=	16'h	c425;
45940	:douta	=	16'h	cc26;
45941	:douta	=	16'h	cc46;
45942	:douta	=	16'h	cc46;
45943	:douta	=	16'h	cc46;
45944	:douta	=	16'h	cc46;
45945	:douta	=	16'h	cc46;
45946	:douta	=	16'h	cc46;
45947	:douta	=	16'h	cc47;
45948	:douta	=	16'h	cc46;
45949	:douta	=	16'h	d467;
45950	:douta	=	16'h	cc66;
45951	:douta	=	16'h	d466;
45952	:douta	=	16'h	cc46;
45953	:douta	=	16'h	cc46;
45954	:douta	=	16'h	d467;
45955	:douta	=	16'h	d467;
45956	:douta	=	16'h	d467;
45957	:douta	=	16'h	cc66;
45958	:douta	=	16'h	cc66;
45959	:douta	=	16'h	d467;
45960	:douta	=	16'h	d467;
45961	:douta	=	16'h	d467;
45962	:douta	=	16'h	d467;
45963	:douta	=	16'h	d466;
45964	:douta	=	16'h	d467;
45965	:douta	=	16'h	d467;
45966	:douta	=	16'h	d467;
45967	:douta	=	16'h	d467;
45968	:douta	=	16'h	d467;
45969	:douta	=	16'h	d488;
45970	:douta	=	16'h	d467;
45971	:douta	=	16'h	d467;
45972	:douta	=	16'h	d467;
45973	:douta	=	16'h	d467;
45974	:douta	=	16'h	d467;
45975	:douta	=	16'h	d467;
45976	:douta	=	16'h	d467;
45977	:douta	=	16'h	d468;
45978	:douta	=	16'h	d468;
45979	:douta	=	16'h	d467;
45980	:douta	=	16'h	d467;
45981	:douta	=	16'h	d467;
45982	:douta	=	16'h	d467;
45983	:douta	=	16'h	d487;
45984	:douta	=	16'h	d467;
45985	:douta	=	16'h	d487;
45986	:douta	=	16'h	d468;
45987	:douta	=	16'h	bccd;
45988	:douta	=	16'h	ce56;
45989	:douta	=	16'h	b44b;
45990	:douta	=	16'h	9430;
45991	:douta	=	16'h	9410;
45992	:douta	=	16'h	8bd0;
45993	:douta	=	16'h	83b0;
45994	:douta	=	16'h	734e;
45995	:douta	=	16'h	734e;
45996	:douta	=	16'h	6b4e;
45997	:douta	=	16'h	62cd;
45998	:douta	=	16'h	62cc;
45999	:douta	=	16'h	49e6;
46000	:douta	=	16'h	41a5;
46001	:douta	=	16'h	5a8a;
46002	:douta	=	16'h	8c0e;
46003	:douta	=	16'h	d614;
46004	:douta	=	16'h	734b;
46005	:douta	=	16'h	8bed;
46006	:douta	=	16'h	acaf;
46007	:douta	=	16'h	bd30;
46008	:douta	=	16'h	c571;
46009	:douta	=	16'h	cdb4;
46010	:douta	=	16'h	cdb3;
46011	:douta	=	16'h	bd52;
46012	:douta	=	16'h	e676;
46013	:douta	=	16'h	de35;
46014	:douta	=	16'h	d614;
46015	:douta	=	16'h	e676;
46016	:douta	=	16'h	de15;
46017	:douta	=	16'h	de15;
46018	:douta	=	16'h	de15;
46019	:douta	=	16'h	de35;
46020	:douta	=	16'h	d5f4;
46021	:douta	=	16'h	d615;
46022	:douta	=	16'h	b513;
46023	:douta	=	16'h	a4d3;
46024	:douta	=	16'h	c596;
46025	:douta	=	16'h	c595;
46026	:douta	=	16'h	9c93;
46027	:douta	=	16'h	b534;
46028	:douta	=	16'h	acf4;
46029	:douta	=	16'h	acf4;
46030	:douta	=	16'h	b515;
46031	:douta	=	16'h	b514;
46032	:douta	=	16'h	a4f4;
46033	:douta	=	16'h	9cb4;
46034	:douta	=	16'h	8c74;
46035	:douta	=	16'h	8432;
46036	:douta	=	16'h	7bd1;
46037	:douta	=	16'h	7bb1;
46038	:douta	=	16'h	7bd1;
46039	:douta	=	16'h	73b1;
46040	:douta	=	16'h	7bd1;
46041	:douta	=	16'h	736f;
46042	:douta	=	16'h	6b0c;
46043	:douta	=	16'h	5a69;
46044	:douta	=	16'h	2903;
46045	:douta	=	16'h	2903;
46046	:douta	=	16'h	41a6;
46047	:douta	=	16'h	62ca;
46048	:douta	=	16'h	5a68;
46049	:douta	=	16'h	5269;
46050	:douta	=	16'h	528b;
46051	:douta	=	16'h	5b50;
46052	:douta	=	16'h	4aef;
46053	:douta	=	16'h	4aef;
46054	:douta	=	16'h	29a9;
46055	:douta	=	16'h	736f;
46056	:douta	=	16'h	31eb;
46057	:douta	=	16'h	1083;
46058	:douta	=	16'h	18e5;
46059	:douta	=	16'h	2126;
46060	:douta	=	16'h	1905;
46061	:douta	=	16'h	4186;
46062	:douta	=	16'h	59e6;
46063	:douta	=	16'h	51e6;
46064	:douta	=	16'h	51c6;
46065	:douta	=	16'h	49c5;
46066	:douta	=	16'h	49c6;
46067	:douta	=	16'h	49a6;
46068	:douta	=	16'h	49a5;
46069	:douta	=	16'h	4186;
46070	:douta	=	16'h	49a6;
46071	:douta	=	16'h	4186;
46072	:douta	=	16'h	4185;
46073	:douta	=	16'h	4185;
46074	:douta	=	16'h	4186;
46075	:douta	=	16'h	3966;
46076	:douta	=	16'h	3966;
46077	:douta	=	16'h	4166;
46078	:douta	=	16'h	3965;
46079	:douta	=	16'h	4166;
46080	:douta	=	16'h	ffbc;
46081	:douta	=	16'h	ffbd;
46082	:douta	=	16'h	fffd;
46083	:douta	=	16'h	de16;
46084	:douta	=	16'h	ee77;
46085	:douta	=	16'h	e677;
46086	:douta	=	16'h	a4f5;
46087	:douta	=	16'h	a493;
46088	:douta	=	16'h	bd55;
46089	:douta	=	16'h	b535;
46090	:douta	=	16'h	cdd6;
46091	:douta	=	16'h	bd75;
46092	:douta	=	16'h	bd55;
46093	:douta	=	16'h	bd76;
46094	:douta	=	16'h	8c53;
46095	:douta	=	16'h	9494;
46096	:douta	=	16'h	8c94;
46097	:douta	=	16'h	8474;
46098	:douta	=	16'h	8474;
46099	:douta	=	16'h	8434;
46100	:douta	=	16'h	8454;
46101	:douta	=	16'h	7c13;
46102	:douta	=	16'h	8475;
46103	:douta	=	16'h	8c74;
46104	:douta	=	16'h	6bb1;
46105	:douta	=	16'h	0841;
46106	:douta	=	16'h	18c3;
46107	:douta	=	16'h	18a2;
46108	:douta	=	16'h	18a3;
46109	:douta	=	16'h	18c3;
46110	:douta	=	16'h	20c3;
46111	:douta	=	16'h	1082;
46112	:douta	=	16'h	1882;
46113	:douta	=	16'h	1861;
46114	:douta	=	16'h	1882;
46115	:douta	=	16'h	1882;
46116	:douta	=	16'h	1881;
46117	:douta	=	16'h	1881;
46118	:douta	=	16'h	18a2;
46119	:douta	=	16'h	2082;
46120	:douta	=	16'h	20a2;
46121	:douta	=	16'h	2082;
46122	:douta	=	16'h	20a2;
46123	:douta	=	16'h	28c2;
46124	:douta	=	16'h	20c2;
46125	:douta	=	16'h	28e3;
46126	:douta	=	16'h	28c2;
46127	:douta	=	16'h	28e2;
46128	:douta	=	16'h	28e2;
46129	:douta	=	16'h	30e3;
46130	:douta	=	16'h	3146;
46131	:douta	=	16'h	2967;
46132	:douta	=	16'h	18a5;
46133	:douta	=	16'h	4123;
46134	:douta	=	16'h	4143;
46135	:douta	=	16'h	4143;
46136	:douta	=	16'h	4964;
46137	:douta	=	16'h	4963;
46138	:douta	=	16'h	4984;
46139	:douta	=	16'h	5184;
46140	:douta	=	16'h	51a4;
46141	:douta	=	16'h	5184;
46142	:douta	=	16'h	5183;
46143	:douta	=	16'h	9d13;
46144	:douta	=	16'h	5983;
46145	:douta	=	16'h	6a04;
46146	:douta	=	16'h	4964;
46147	:douta	=	16'h	7224;
46148	:douta	=	16'h	6a04;
46149	:douta	=	16'h	7224;
46150	:douta	=	16'h	7224;
46151	:douta	=	16'h	7224;
46152	:douta	=	16'h	7244;
46153	:douta	=	16'h	7244;
46154	:douta	=	16'h	7224;
46155	:douta	=	16'h	7224;
46156	:douta	=	16'h	7a44;
46157	:douta	=	16'h	7a44;
46158	:douta	=	16'h	8285;
46159	:douta	=	16'h	8284;
46160	:douta	=	16'h	8aa4;
46161	:douta	=	16'h	8aa4;
46162	:douta	=	16'h	8ac4;
46163	:douta	=	16'h	92e4;
46164	:douta	=	16'h	9304;
46165	:douta	=	16'h	9304;
46166	:douta	=	16'h	9b05;
46167	:douta	=	16'h	9b25;
46168	:douta	=	16'h	a325;
46169	:douta	=	16'h	a345;
46170	:douta	=	16'h	ab64;
46171	:douta	=	16'h	ab65;
46172	:douta	=	16'h	ab85;
46173	:douta	=	16'h	b385;
46174	:douta	=	16'h	b385;
46175	:douta	=	16'h	b3a5;
46176	:douta	=	16'h	b3c5;
46177	:douta	=	16'h	b3c5;
46178	:douta	=	16'h	bbe6;
46179	:douta	=	16'h	bbe5;
46180	:douta	=	16'h	bbe5;
46181	:douta	=	16'h	bbe5;
46182	:douta	=	16'h	bbe5;
46183	:douta	=	16'h	bc06;
46184	:douta	=	16'h	bbe5;
46185	:douta	=	16'h	c406;
46186	:douta	=	16'h	c405;
46187	:douta	=	16'h	c426;
46188	:douta	=	16'h	c426;
46189	:douta	=	16'h	c426;
46190	:douta	=	16'h	c426;
46191	:douta	=	16'h	c425;
46192	:douta	=	16'h	c425;
46193	:douta	=	16'h	c425;
46194	:douta	=	16'h	c405;
46195	:douta	=	16'h	c425;
46196	:douta	=	16'h	cc26;
46197	:douta	=	16'h	cc26;
46198	:douta	=	16'h	cc26;
46199	:douta	=	16'h	cc26;
46200	:douta	=	16'h	cc46;
46201	:douta	=	16'h	cc46;
46202	:douta	=	16'h	cc46;
46203	:douta	=	16'h	cc46;
46204	:douta	=	16'h	cc46;
46205	:douta	=	16'h	cc46;
46206	:douta	=	16'h	cc46;
46207	:douta	=	16'h	cc46;
46208	:douta	=	16'h	d467;
46209	:douta	=	16'h	d467;
46210	:douta	=	16'h	d467;
46211	:douta	=	16'h	d467;
46212	:douta	=	16'h	d467;
46213	:douta	=	16'h	cc66;
46214	:douta	=	16'h	d466;
46215	:douta	=	16'h	cc47;
46216	:douta	=	16'h	d467;
46217	:douta	=	16'h	d467;
46218	:douta	=	16'h	cc66;
46219	:douta	=	16'h	d466;
46220	:douta	=	16'h	d467;
46221	:douta	=	16'h	d467;
46222	:douta	=	16'h	d467;
46223	:douta	=	16'h	d467;
46224	:douta	=	16'h	d468;
46225	:douta	=	16'h	d468;
46226	:douta	=	16'h	d467;
46227	:douta	=	16'h	d467;
46228	:douta	=	16'h	d467;
46229	:douta	=	16'h	d467;
46230	:douta	=	16'h	d467;
46231	:douta	=	16'h	d467;
46232	:douta	=	16'h	d467;
46233	:douta	=	16'h	d467;
46234	:douta	=	16'h	d467;
46235	:douta	=	16'h	d467;
46236	:douta	=	16'h	d467;
46237	:douta	=	16'h	d467;
46238	:douta	=	16'h	d467;
46239	:douta	=	16'h	d467;
46240	:douta	=	16'h	d467;
46241	:douta	=	16'h	d467;
46242	:douta	=	16'h	d468;
46243	:douta	=	16'h	b4ad;
46244	:douta	=	16'h	ce56;
46245	:douta	=	16'h	dc65;
46246	:douta	=	16'h	8c31;
46247	:douta	=	16'h	8bef;
46248	:douta	=	16'h	838f;
46249	:douta	=	16'h	83af;
46250	:douta	=	16'h	6b4e;
46251	:douta	=	16'h	734e;
46252	:douta	=	16'h	6b4d;
46253	:douta	=	16'h	41c8;
46254	:douta	=	16'h	41c6;
46255	:douta	=	16'h	5248;
46256	:douta	=	16'h	6b2c;
46257	:douta	=	16'h	7b6d;
46258	:douta	=	16'h	d615;
46259	:douta	=	16'h	de14;
46260	:douta	=	16'h	8bac;
46261	:douta	=	16'h	bd51;
46262	:douta	=	16'h	bd11;
46263	:douta	=	16'h	cd71;
46264	:douta	=	16'h	cdb2;
46265	:douta	=	16'h	d5d4;
46266	:douta	=	16'h	c5b3;
46267	:douta	=	16'h	cdd4;
46268	:douta	=	16'h	e697;
46269	:douta	=	16'h	de56;
46270	:douta	=	16'h	cdb3;
46271	:douta	=	16'h	e676;
46272	:douta	=	16'h	de15;
46273	:douta	=	16'h	d5d4;
46274	:douta	=	16'h	de15;
46275	:douta	=	16'h	d5d4;
46276	:douta	=	16'h	bd74;
46277	:douta	=	16'h	cd94;
46278	:douta	=	16'h	c574;
46279	:douta	=	16'h	a4b3;
46280	:douta	=	16'h	bd75;
46281	:douta	=	16'h	bd55;
46282	:douta	=	16'h	94b3;
46283	:douta	=	16'h	a4b4;
46284	:douta	=	16'h	9cb4;
46285	:douta	=	16'h	a4b4;
46286	:douta	=	16'h	a4d5;
46287	:douta	=	16'h	a4d5;
46288	:douta	=	16'h	9cb4;
46289	:douta	=	16'h	9cb4;
46290	:douta	=	16'h	8c52;
46291	:douta	=	16'h	8412;
46292	:douta	=	16'h	73b0;
46293	:douta	=	16'h	7370;
46294	:douta	=	16'h	6b6f;
46295	:douta	=	16'h	732e;
46296	:douta	=	16'h	6b2d;
46297	:douta	=	16'h	6b0c;
46298	:douta	=	16'h	2903;
46299	:douta	=	16'h	2103;
46300	:douta	=	16'h	49e6;
46301	:douta	=	16'h	5a68;
46302	:douta	=	16'h	62ea;
46303	:douta	=	16'h	736c;
46304	:douta	=	16'h	83ad;
46305	:douta	=	16'h	7bae;
46306	:douta	=	16'h	6b6f;
46307	:douta	=	16'h	5b30;
46308	:douta	=	16'h	52ef;
46309	:douta	=	16'h	4af0;
46310	:douta	=	16'h	2989;
46311	:douta	=	16'h	6b2e;
46312	:douta	=	16'h	530f;
46313	:douta	=	16'h	1906;
46314	:douta	=	16'h	10a3;
46315	:douta	=	16'h	1925;
46316	:douta	=	16'h	1906;
46317	:douta	=	16'h	59e6;
46318	:douta	=	16'h	51e6;
46319	:douta	=	16'h	51c6;
46320	:douta	=	16'h	51c5;
46321	:douta	=	16'h	49c6;
46322	:douta	=	16'h	49c6;
46323	:douta	=	16'h	49a6;
46324	:douta	=	16'h	49a5;
46325	:douta	=	16'h	4185;
46326	:douta	=	16'h	49a6;
46327	:douta	=	16'h	4185;
46328	:douta	=	16'h	4185;
46329	:douta	=	16'h	41a6;
46330	:douta	=	16'h	4165;
46331	:douta	=	16'h	4186;
46332	:douta	=	16'h	4165;
46333	:douta	=	16'h	4186;
46334	:douta	=	16'h	4165;
46335	:douta	=	16'h	3966;
46336	:douta	=	16'h	ffbd;
46337	:douta	=	16'h	ffdd;
46338	:douta	=	16'h	ffdd;
46339	:douta	=	16'h	de16;
46340	:douta	=	16'h	e677;
46341	:douta	=	16'h	d5f6;
46342	:douta	=	16'h	a4d4;
46343	:douta	=	16'h	9c93;
46344	:douta	=	16'h	bd96;
46345	:douta	=	16'h	c595;
46346	:douta	=	16'h	cdb5;
46347	:douta	=	16'h	bd55;
46348	:douta	=	16'h	bd75;
46349	:douta	=	16'h	9cd5;
46350	:douta	=	16'h	9494;
46351	:douta	=	16'h	94b5;
46352	:douta	=	16'h	8c74;
46353	:douta	=	16'h	8c74;
46354	:douta	=	16'h	8474;
46355	:douta	=	16'h	8454;
46356	:douta	=	16'h	7c33;
46357	:douta	=	16'h	8454;
46358	:douta	=	16'h	8454;
46359	:douta	=	16'h	94f7;
46360	:douta	=	16'h	2925;
46361	:douta	=	16'h	1861;
46362	:douta	=	16'h	20e3;
46363	:douta	=	16'h	20c2;
46364	:douta	=	16'h	18e2;
46365	:douta	=	16'h	18a3;
46366	:douta	=	16'h	18c3;
46367	:douta	=	16'h	1082;
46368	:douta	=	16'h	1882;
46369	:douta	=	16'h	1882;
46370	:douta	=	16'h	1882;
46371	:douta	=	16'h	1882;
46372	:douta	=	16'h	1881;
46373	:douta	=	16'h	2082;
46374	:douta	=	16'h	20a2;
46375	:douta	=	16'h	1881;
46376	:douta	=	16'h	2082;
46377	:douta	=	16'h	20a2;
46378	:douta	=	16'h	20a2;
46379	:douta	=	16'h	20a2;
46380	:douta	=	16'h	28e3;
46381	:douta	=	16'h	28c2;
46382	:douta	=	16'h	28e2;
46383	:douta	=	16'h	28e2;
46384	:douta	=	16'h	3103;
46385	:douta	=	16'h	3103;
46386	:douta	=	16'h	39c8;
46387	:douta	=	16'h	2126;
46388	:douta	=	16'h	18c4;
46389	:douta	=	16'h	4163;
46390	:douta	=	16'h	4143;
46391	:douta	=	16'h	4163;
46392	:douta	=	16'h	4963;
46393	:douta	=	16'h	4984;
46394	:douta	=	16'h	5184;
46395	:douta	=	16'h	51a4;
46396	:douta	=	16'h	59a4;
46397	:douta	=	16'h	5163;
46398	:douta	=	16'h	5a05;
46399	:douta	=	16'h	9cd1;
46400	:douta	=	16'h	61c4;
46401	:douta	=	16'h	6204;
46402	:douta	=	16'h	4963;
46403	:douta	=	16'h	61c4;
46404	:douta	=	16'h	7224;
46405	:douta	=	16'h	7224;
46406	:douta	=	16'h	7224;
46407	:douta	=	16'h	7244;
46408	:douta	=	16'h	7244;
46409	:douta	=	16'h	7a65;
46410	:douta	=	16'h	7a44;
46411	:douta	=	16'h	7244;
46412	:douta	=	16'h	7a64;
46413	:douta	=	16'h	7a64;
46414	:douta	=	16'h	8264;
46415	:douta	=	16'h	82a4;
46416	:douta	=	16'h	82a4;
46417	:douta	=	16'h	8ac4;
46418	:douta	=	16'h	8ac4;
46419	:douta	=	16'h	9304;
46420	:douta	=	16'h	9b25;
46421	:douta	=	16'h	9305;
46422	:douta	=	16'h	9b45;
46423	:douta	=	16'h	9b25;
46424	:douta	=	16'h	a345;
46425	:douta	=	16'h	a345;
46426	:douta	=	16'h	ab64;
46427	:douta	=	16'h	ab85;
46428	:douta	=	16'h	b385;
46429	:douta	=	16'h	b385;
46430	:douta	=	16'h	b385;
46431	:douta	=	16'h	b3a5;
46432	:douta	=	16'h	bbc5;
46433	:douta	=	16'h	bbc5;
46434	:douta	=	16'h	bbe6;
46435	:douta	=	16'h	bbe6;
46436	:douta	=	16'h	bbe5;
46437	:douta	=	16'h	bbe5;
46438	:douta	=	16'h	bbe5;
46439	:douta	=	16'h	bc06;
46440	:douta	=	16'h	bc06;
46441	:douta	=	16'h	c406;
46442	:douta	=	16'h	c406;
46443	:douta	=	16'h	c405;
46444	:douta	=	16'h	c426;
46445	:douta	=	16'h	cc26;
46446	:douta	=	16'h	c426;
46447	:douta	=	16'h	c425;
46448	:douta	=	16'h	cc26;
46449	:douta	=	16'h	c425;
46450	:douta	=	16'h	cc26;
46451	:douta	=	16'h	c425;
46452	:douta	=	16'h	cc46;
46453	:douta	=	16'h	cc26;
46454	:douta	=	16'h	cc46;
46455	:douta	=	16'h	cc46;
46456	:douta	=	16'h	cc46;
46457	:douta	=	16'h	cc47;
46458	:douta	=	16'h	cc47;
46459	:douta	=	16'h	cc46;
46460	:douta	=	16'h	cc46;
46461	:douta	=	16'h	cc46;
46462	:douta	=	16'h	cc47;
46463	:douta	=	16'h	cc67;
46464	:douta	=	16'h	cc47;
46465	:douta	=	16'h	d467;
46466	:douta	=	16'h	d467;
46467	:douta	=	16'h	d467;
46468	:douta	=	16'h	d467;
46469	:douta	=	16'h	d467;
46470	:douta	=	16'h	cc66;
46471	:douta	=	16'h	d467;
46472	:douta	=	16'h	d467;
46473	:douta	=	16'h	cc47;
46474	:douta	=	16'h	d467;
46475	:douta	=	16'h	d467;
46476	:douta	=	16'h	d467;
46477	:douta	=	16'h	d467;
46478	:douta	=	16'h	d467;
46479	:douta	=	16'h	d468;
46480	:douta	=	16'h	d468;
46481	:douta	=	16'h	d467;
46482	:douta	=	16'h	d467;
46483	:douta	=	16'h	d487;
46484	:douta	=	16'h	d467;
46485	:douta	=	16'h	d467;
46486	:douta	=	16'h	d467;
46487	:douta	=	16'h	d467;
46488	:douta	=	16'h	d467;
46489	:douta	=	16'h	d467;
46490	:douta	=	16'h	d467;
46491	:douta	=	16'h	d467;
46492	:douta	=	16'h	d487;
46493	:douta	=	16'h	d487;
46494	:douta	=	16'h	d467;
46495	:douta	=	16'h	d468;
46496	:douta	=	16'h	d488;
46497	:douta	=	16'h	d467;
46498	:douta	=	16'h	d468;
46499	:douta	=	16'h	b4cd;
46500	:douta	=	16'h	ce56;
46501	:douta	=	16'h	cc46;
46502	:douta	=	16'h	dca6;
46503	:douta	=	16'h	a44e;
46504	:douta	=	16'h	83af;
46505	:douta	=	16'h	62ec;
46506	:douta	=	16'h	3986;
46507	:douta	=	16'h	4a28;
46508	:douta	=	16'h	5247;
46509	:douta	=	16'h	9c4f;
46510	:douta	=	16'h	736b;
46511	:douta	=	16'h	a490;
46512	:douta	=	16'h	9cb0;
46513	:douta	=	16'h	d614;
46514	:douta	=	16'h	b532;
46515	:douta	=	16'h	8bee;
46516	:douta	=	16'h	d5d3;
46517	:douta	=	16'h	d5f3;
46518	:douta	=	16'h	de14;
46519	:douta	=	16'h	d5d3;
46520	:douta	=	16'h	ddf4;
46521	:douta	=	16'h	d5d4;
46522	:douta	=	16'h	cdb3;
46523	:douta	=	16'h	e677;
46524	:douta	=	16'h	de56;
46525	:douta	=	16'h	d5d4;
46526	:douta	=	16'h	bd33;
46527	:douta	=	16'h	bd74;
46528	:douta	=	16'h	d5d5;
46529	:douta	=	16'h	c574;
46530	:douta	=	16'h	bd54;
46531	:douta	=	16'h	b554;
46532	:douta	=	16'h	ad14;
46533	:douta	=	16'h	a4d4;
46534	:douta	=	16'h	acf4;
46535	:douta	=	16'h	ad14;
46536	:douta	=	16'h	a4f4;
46537	:douta	=	16'h	9cd5;
46538	:douta	=	16'h	9494;
46539	:douta	=	16'h	8c53;
46540	:douta	=	16'h	8452;
46541	:douta	=	16'h	8432;
46542	:douta	=	16'h	8432;
46543	:douta	=	16'h	8c33;
46544	:douta	=	16'h	8432;
46545	:douta	=	16'h	7bf1;
46546	:douta	=	16'h	8432;
46547	:douta	=	16'h	7bf1;
46548	:douta	=	16'h	62ed;
46549	:douta	=	16'h	5248;
46550	:douta	=	16'h	3944;
46551	:douta	=	16'h	3944;
46552	:douta	=	16'h	49e5;
46553	:douta	=	16'h	5a88;
46554	:douta	=	16'h	5268;
46555	:douta	=	16'h	5a89;
46556	:douta	=	16'h	6aea;
46557	:douta	=	16'h	734b;
46558	:douta	=	16'h	7b8c;
46559	:douta	=	16'h	83ad;
46560	:douta	=	16'h	940e;
46561	:douta	=	16'h	524a;
46562	:douta	=	16'h	18e6;
46563	:douta	=	16'h	2126;
46564	:douta	=	16'h	2146;
46565	:douta	=	16'h	2146;
46566	:douta	=	16'h	2147;
46567	:douta	=	16'h	5249;
46568	:douta	=	16'h	2106;
46569	:douta	=	16'h	3a2b;
46570	:douta	=	16'h	3a2b;
46571	:douta	=	16'h	18e5;
46572	:douta	=	16'h	10e6;
46573	:douta	=	16'h	5a06;
46574	:douta	=	16'h	59e6;
46575	:douta	=	16'h	51c6;
46576	:douta	=	16'h	51c6;
46577	:douta	=	16'h	49c6;
46578	:douta	=	16'h	49c6;
46579	:douta	=	16'h	49a6;
46580	:douta	=	16'h	49c6;
46581	:douta	=	16'h	49a6;
46582	:douta	=	16'h	4186;
46583	:douta	=	16'h	4186;
46584	:douta	=	16'h	41a6;
46585	:douta	=	16'h	4185;
46586	:douta	=	16'h	4185;
46587	:douta	=	16'h	4185;
46588	:douta	=	16'h	4186;
46589	:douta	=	16'h	4166;
46590	:douta	=	16'h	4166;
46591	:douta	=	16'h	4166;
46592	:douta	=	16'h	ffbd;
46593	:douta	=	16'h	ffde;
46594	:douta	=	16'h	ff7c;
46595	:douta	=	16'h	de36;
46596	:douta	=	16'h	e677;
46597	:douta	=	16'h	c5b5;
46598	:douta	=	16'h	a4b4;
46599	:douta	=	16'h	9c93;
46600	:douta	=	16'h	ad35;
46601	:douta	=	16'h	cdd6;
46602	:douta	=	16'h	c5b5;
46603	:douta	=	16'h	bd55;
46604	:douta	=	16'h	bd75;
46605	:douta	=	16'h	9474;
46606	:douta	=	16'h	94b5;
46607	:douta	=	16'h	94b5;
46608	:douta	=	16'h	8c94;
46609	:douta	=	16'h	8c75;
46610	:douta	=	16'h	8454;
46611	:douta	=	16'h	8454;
46612	:douta	=	16'h	7c13;
46613	:douta	=	16'h	8454;
46614	:douta	=	16'h	8474;
46615	:douta	=	16'h	9d58;
46616	:douta	=	16'h	0800;
46617	:douta	=	16'h	20c2;
46618	:douta	=	16'h	20c3;
46619	:douta	=	16'h	18a3;
46620	:douta	=	16'h	18c3;
46621	:douta	=	16'h	18c3;
46622	:douta	=	16'h	20e3;
46623	:douta	=	16'h	1861;
46624	:douta	=	16'h	1882;
46625	:douta	=	16'h	1882;
46626	:douta	=	16'h	1882;
46627	:douta	=	16'h	1881;
46628	:douta	=	16'h	18a2;
46629	:douta	=	16'h	20a2;
46630	:douta	=	16'h	2082;
46631	:douta	=	16'h	1881;
46632	:douta	=	16'h	2082;
46633	:douta	=	16'h	2082;
46634	:douta	=	16'h	20a2;
46635	:douta	=	16'h	20a2;
46636	:douta	=	16'h	28c2;
46637	:douta	=	16'h	28c2;
46638	:douta	=	16'h	30e2;
46639	:douta	=	16'h	30e3;
46640	:douta	=	16'h	30e2;
46641	:douta	=	16'h	3144;
46642	:douta	=	16'h	39e9;
46643	:douta	=	16'h	2126;
46644	:douta	=	16'h	18c4;
46645	:douta	=	16'h	4143;
46646	:douta	=	16'h	4143;
46647	:douta	=	16'h	4963;
46648	:douta	=	16'h	4963;
46649	:douta	=	16'h	4963;
46650	:douta	=	16'h	5184;
46651	:douta	=	16'h	51a4;
46652	:douta	=	16'h	51a4;
46653	:douta	=	16'h	5163;
46654	:douta	=	16'h	6267;
46655	:douta	=	16'h	9c6f;
46656	:douta	=	16'h	69e4;
46657	:douta	=	16'h	6a04;
46658	:douta	=	16'h	4984;
46659	:douta	=	16'h	61c4;
46660	:douta	=	16'h	7224;
46661	:douta	=	16'h	6a24;
46662	:douta	=	16'h	7224;
46663	:douta	=	16'h	7a44;
46664	:douta	=	16'h	7244;
46665	:douta	=	16'h	7244;
46666	:douta	=	16'h	7a44;
46667	:douta	=	16'h	7244;
46668	:douta	=	16'h	7a64;
46669	:douta	=	16'h	7a64;
46670	:douta	=	16'h	8284;
46671	:douta	=	16'h	82a4;
46672	:douta	=	16'h	8aa4;
46673	:douta	=	16'h	8ac4;
46674	:douta	=	16'h	8ac5;
46675	:douta	=	16'h	92e4;
46676	:douta	=	16'h	9305;
46677	:douta	=	16'h	9b25;
46678	:douta	=	16'h	9b05;
46679	:douta	=	16'h	9b25;
46680	:douta	=	16'h	a345;
46681	:douta	=	16'h	a345;
46682	:douta	=	16'h	ab64;
46683	:douta	=	16'h	ab85;
46684	:douta	=	16'h	b385;
46685	:douta	=	16'h	b385;
46686	:douta	=	16'h	b385;
46687	:douta	=	16'h	b3a5;
46688	:douta	=	16'h	bbc6;
46689	:douta	=	16'h	bbc5;
46690	:douta	=	16'h	bbe6;
46691	:douta	=	16'h	bbe6;
46692	:douta	=	16'h	bbe5;
46693	:douta	=	16'h	bbe5;
46694	:douta	=	16'h	bbe5;
46695	:douta	=	16'h	bc06;
46696	:douta	=	16'h	c406;
46697	:douta	=	16'h	c406;
46698	:douta	=	16'h	c406;
46699	:douta	=	16'h	c426;
46700	:douta	=	16'h	c426;
46701	:douta	=	16'h	c426;
46702	:douta	=	16'h	cc26;
46703	:douta	=	16'h	c426;
46704	:douta	=	16'h	cc26;
46705	:douta	=	16'h	cc26;
46706	:douta	=	16'h	cc26;
46707	:douta	=	16'h	cc26;
46708	:douta	=	16'h	cc46;
46709	:douta	=	16'h	cc46;
46710	:douta	=	16'h	cc46;
46711	:douta	=	16'h	cc26;
46712	:douta	=	16'h	cc46;
46713	:douta	=	16'h	cc46;
46714	:douta	=	16'h	cc46;
46715	:douta	=	16'h	cc46;
46716	:douta	=	16'h	cc46;
46717	:douta	=	16'h	cc46;
46718	:douta	=	16'h	cc46;
46719	:douta	=	16'h	cc47;
46720	:douta	=	16'h	d467;
46721	:douta	=	16'h	cc47;
46722	:douta	=	16'h	d467;
46723	:douta	=	16'h	d467;
46724	:douta	=	16'h	d467;
46725	:douta	=	16'h	d467;
46726	:douta	=	16'h	cc66;
46727	:douta	=	16'h	d467;
46728	:douta	=	16'h	cc47;
46729	:douta	=	16'h	d467;
46730	:douta	=	16'h	d467;
46731	:douta	=	16'h	cc67;
46732	:douta	=	16'h	d466;
46733	:douta	=	16'h	d467;
46734	:douta	=	16'h	d467;
46735	:douta	=	16'h	d487;
46736	:douta	=	16'h	d467;
46737	:douta	=	16'h	d467;
46738	:douta	=	16'h	d488;
46739	:douta	=	16'h	d467;
46740	:douta	=	16'h	d467;
46741	:douta	=	16'h	d487;
46742	:douta	=	16'h	d467;
46743	:douta	=	16'h	d467;
46744	:douta	=	16'h	cc67;
46745	:douta	=	16'h	d487;
46746	:douta	=	16'h	d487;
46747	:douta	=	16'h	d487;
46748	:douta	=	16'h	d487;
46749	:douta	=	16'h	d467;
46750	:douta	=	16'h	d467;
46751	:douta	=	16'h	d468;
46752	:douta	=	16'h	d488;
46753	:douta	=	16'h	d487;
46754	:douta	=	16'h	d468;
46755	:douta	=	16'h	bccd;
46756	:douta	=	16'h	ce56;
46757	:douta	=	16'h	cc46;
46758	:douta	=	16'h	dc86;
46759	:douta	=	16'h	cc89;
46760	:douta	=	16'h	6b2d;
46761	:douta	=	16'h	62ca;
46762	:douta	=	16'h	6aeb;
46763	:douta	=	16'h	7b8d;
46764	:douta	=	16'h	b4f2;
46765	:douta	=	16'h	6aea;
46766	:douta	=	16'h	8c2e;
46767	:douta	=	16'h	acd2;
46768	:douta	=	16'h	acf2;
46769	:douta	=	16'h	de56;
46770	:douta	=	16'h	a490;
46771	:douta	=	16'h	a48f;
46772	:douta	=	16'h	de15;
46773	:douta	=	16'h	de15;
46774	:douta	=	16'h	d5f5;
46775	:douta	=	16'h	d614;
46776	:douta	=	16'h	de15;
46777	:douta	=	16'h	d5f4;
46778	:douta	=	16'h	d5f4;
46779	:douta	=	16'h	de36;
46780	:douta	=	16'h	de16;
46781	:douta	=	16'h	d5f5;
46782	:douta	=	16'h	bd33;
46783	:douta	=	16'h	acf3;
46784	:douta	=	16'h	c594;
46785	:douta	=	16'h	bd54;
46786	:douta	=	16'h	b535;
46787	:douta	=	16'h	a4f5;
46788	:douta	=	16'h	9cb4;
46789	:douta	=	16'h	a4d5;
46790	:douta	=	16'h	9cb4;
46791	:douta	=	16'h	9cb4;
46792	:douta	=	16'h	94b4;
46793	:douta	=	16'h	a4d5;
46794	:douta	=	16'h	7c12;
46795	:douta	=	16'h	8433;
46796	:douta	=	16'h	8452;
46797	:douta	=	16'h	9493;
46798	:douta	=	16'h	8432;
46799	:douta	=	16'h	8412;
46800	:douta	=	16'h	7bf1;
46801	:douta	=	16'h	7bd0;
46802	:douta	=	16'h	7baf;
46803	:douta	=	16'h	5aaa;
46804	:douta	=	16'h	41a5;
46805	:douta	=	16'h	0000;
46806	:douta	=	16'h	0000;
46807	:douta	=	16'h	5aa8;
46808	:douta	=	16'h	5aa8;
46809	:douta	=	16'h	8c0e;
46810	:douta	=	16'h	6aeb;
46811	:douta	=	16'h	6acb;
46812	:douta	=	16'h	732b;
46813	:douta	=	16'h	7b8c;
46814	:douta	=	16'h	838d;
46815	:douta	=	16'h	8bce;
46816	:douta	=	16'h	9c90;
46817	:douta	=	16'h	524a;
46818	:douta	=	16'h	2127;
46819	:douta	=	16'h	18e5;
46820	:douta	=	16'h	10c4;
46821	:douta	=	16'h	10a4;
46822	:douta	=	16'h	10a4;
46823	:douta	=	16'h	39a6;
46824	:douta	=	16'h	08a3;
46825	:douta	=	16'h	2126;
46826	:douta	=	16'h	2167;
46827	:douta	=	16'h	2167;
46828	:douta	=	16'h	08a4;
46829	:douta	=	16'h	6247;
46830	:douta	=	16'h	51e6;
46831	:douta	=	16'h	51c6;
46832	:douta	=	16'h	49c6;
46833	:douta	=	16'h	49c6;
46834	:douta	=	16'h	49c6;
46835	:douta	=	16'h	49a6;
46836	:douta	=	16'h	49a6;
46837	:douta	=	16'h	49a6;
46838	:douta	=	16'h	4186;
46839	:douta	=	16'h	49a6;
46840	:douta	=	16'h	4185;
46841	:douta	=	16'h	4185;
46842	:douta	=	16'h	4185;
46843	:douta	=	16'h	4185;
46844	:douta	=	16'h	4186;
46845	:douta	=	16'h	4186;
46846	:douta	=	16'h	4186;
46847	:douta	=	16'h	4186;
46848	:douta	=	16'h	ffbd;
46849	:douta	=	16'h	ffbc;
46850	:douta	=	16'h	de16;
46851	:douta	=	16'h	e698;
46852	:douta	=	16'h	d5f6;
46853	:douta	=	16'h	a4f4;
46854	:douta	=	16'h	9c93;
46855	:douta	=	16'h	ad15;
46856	:douta	=	16'h	b515;
46857	:douta	=	16'h	cdb5;
46858	:douta	=	16'h	c595;
46859	:douta	=	16'h	bd55;
46860	:douta	=	16'h	b576;
46861	:douta	=	16'h	8c53;
46862	:douta	=	16'h	94b5;
46863	:douta	=	16'h	9494;
46864	:douta	=	16'h	8c74;
46865	:douta	=	16'h	8c74;
46866	:douta	=	16'h	8454;
46867	:douta	=	16'h	8434;
46868	:douta	=	16'h	8454;
46869	:douta	=	16'h	8454;
46870	:douta	=	16'h	8c74;
46871	:douta	=	16'h	73f2;
46872	:douta	=	16'h	20a2;
46873	:douta	=	16'h	20e3;
46874	:douta	=	16'h	20a3;
46875	:douta	=	16'h	20c3;
46876	:douta	=	16'h	18a3;
46877	:douta	=	16'h	20e3;
46878	:douta	=	16'h	18c3;
46879	:douta	=	16'h	1882;
46880	:douta	=	16'h	1882;
46881	:douta	=	16'h	1882;
46882	:douta	=	16'h	1882;
46883	:douta	=	16'h	18a2;
46884	:douta	=	16'h	2082;
46885	:douta	=	16'h	1881;
46886	:douta	=	16'h	20a2;
46887	:douta	=	16'h	20a2;
46888	:douta	=	16'h	20a2;
46889	:douta	=	16'h	20a2;
46890	:douta	=	16'h	20a2;
46891	:douta	=	16'h	20c2;
46892	:douta	=	16'h	28e2;
46893	:douta	=	16'h	28e2;
46894	:douta	=	16'h	28e2;
46895	:douta	=	16'h	28e2;
46896	:douta	=	16'h	3103;
46897	:douta	=	16'h	3146;
46898	:douta	=	16'h	31c9;
46899	:douta	=	16'h	18e5;
46900	:douta	=	16'h	28e3;
46901	:douta	=	16'h	4143;
46902	:douta	=	16'h	4163;
46903	:douta	=	16'h	4963;
46904	:douta	=	16'h	4984;
46905	:douta	=	16'h	5184;
46906	:douta	=	16'h	5184;
46907	:douta	=	16'h	59a4;
46908	:douta	=	16'h	51a4;
46909	:douta	=	16'h	5183;
46910	:douta	=	16'h	6aeb;
46911	:douta	=	16'h	8bec;
46912	:douta	=	16'h	6a04;
46913	:douta	=	16'h	6204;
46914	:douta	=	16'h	4984;
46915	:douta	=	16'h	59a4;
46916	:douta	=	16'h	7224;
46917	:douta	=	16'h	7224;
46918	:douta	=	16'h	7244;
46919	:douta	=	16'h	7a64;
46920	:douta	=	16'h	7a64;
46921	:douta	=	16'h	7a44;
46922	:douta	=	16'h	7244;
46923	:douta	=	16'h	7a44;
46924	:douta	=	16'h	7a64;
46925	:douta	=	16'h	7a64;
46926	:douta	=	16'h	8285;
46927	:douta	=	16'h	82a5;
46928	:douta	=	16'h	8aa4;
46929	:douta	=	16'h	8ac4;
46930	:douta	=	16'h	8ae4;
46931	:douta	=	16'h	9304;
46932	:douta	=	16'h	9b05;
46933	:douta	=	16'h	9b05;
46934	:douta	=	16'h	9b25;
46935	:douta	=	16'h	a325;
46936	:douta	=	16'h	a345;
46937	:douta	=	16'h	a365;
46938	:douta	=	16'h	ab65;
46939	:douta	=	16'h	ab85;
46940	:douta	=	16'h	ab85;
46941	:douta	=	16'h	b3a5;
46942	:douta	=	16'h	b3a5;
46943	:douta	=	16'h	b3a6;
46944	:douta	=	16'h	b3a6;
46945	:douta	=	16'h	bbe6;
46946	:douta	=	16'h	bbe6;
46947	:douta	=	16'h	bbe6;
46948	:douta	=	16'h	bbe5;
46949	:douta	=	16'h	c406;
46950	:douta	=	16'h	c406;
46951	:douta	=	16'h	bc06;
46952	:douta	=	16'h	bc06;
46953	:douta	=	16'h	c406;
46954	:douta	=	16'h	c405;
46955	:douta	=	16'h	c406;
46956	:douta	=	16'h	c426;
46957	:douta	=	16'h	c426;
46958	:douta	=	16'h	c426;
46959	:douta	=	16'h	cc47;
46960	:douta	=	16'h	cc46;
46961	:douta	=	16'h	c426;
46962	:douta	=	16'h	c426;
46963	:douta	=	16'h	cc46;
46964	:douta	=	16'h	cc46;
46965	:douta	=	16'h	cc46;
46966	:douta	=	16'h	cc47;
46967	:douta	=	16'h	cc47;
46968	:douta	=	16'h	cc46;
46969	:douta	=	16'h	cc46;
46970	:douta	=	16'h	cc46;
46971	:douta	=	16'h	cc46;
46972	:douta	=	16'h	cc46;
46973	:douta	=	16'h	cc46;
46974	:douta	=	16'h	cc47;
46975	:douta	=	16'h	cc46;
46976	:douta	=	16'h	cc47;
46977	:douta	=	16'h	cc47;
46978	:douta	=	16'h	d467;
46979	:douta	=	16'h	d467;
46980	:douta	=	16'h	d467;
46981	:douta	=	16'h	d467;
46982	:douta	=	16'h	d467;
46983	:douta	=	16'h	cc67;
46984	:douta	=	16'h	d467;
46985	:douta	=	16'h	d467;
46986	:douta	=	16'h	d467;
46987	:douta	=	16'h	d467;
46988	:douta	=	16'h	cc67;
46989	:douta	=	16'h	d467;
46990	:douta	=	16'h	cc67;
46991	:douta	=	16'h	d467;
46992	:douta	=	16'h	d467;
46993	:douta	=	16'h	d467;
46994	:douta	=	16'h	d467;
46995	:douta	=	16'h	d467;
46996	:douta	=	16'h	d487;
46997	:douta	=	16'h	d467;
46998	:douta	=	16'h	d487;
46999	:douta	=	16'h	d487;
47000	:douta	=	16'h	d487;
47001	:douta	=	16'h	d467;
47002	:douta	=	16'h	d467;
47003	:douta	=	16'h	d467;
47004	:douta	=	16'h	d488;
47005	:douta	=	16'h	d487;
47006	:douta	=	16'h	d467;
47007	:douta	=	16'h	d487;
47008	:douta	=	16'h	d468;
47009	:douta	=	16'h	d467;
47010	:douta	=	16'h	d468;
47011	:douta	=	16'h	bcce;
47012	:douta	=	16'h	ce77;
47013	:douta	=	16'h	cc46;
47014	:douta	=	16'h	cc87;
47015	:douta	=	16'h	d486;
47016	:douta	=	16'h	9430;
47017	:douta	=	16'h	940f;
47018	:douta	=	16'h	7b6c;
47019	:douta	=	16'h	9c2e;
47020	:douta	=	16'h	734a;
47021	:douta	=	16'h	c571;
47022	:douta	=	16'h	bd52;
47023	:douta	=	16'h	bd73;
47024	:douta	=	16'h	cdf5;
47025	:douta	=	16'h	cdd5;
47026	:douta	=	16'h	9c8f;
47027	:douta	=	16'h	cdd6;
47028	:douta	=	16'h	d615;
47029	:douta	=	16'h	de56;
47030	:douta	=	16'h	d5d4;
47031	:douta	=	16'h	d5f4;
47032	:douta	=	16'h	d5f4;
47033	:douta	=	16'h	d5d3;
47034	:douta	=	16'h	cdd3;
47035	:douta	=	16'h	bd33;
47036	:douta	=	16'h	b514;
47037	:douta	=	16'h	b513;
47038	:douta	=	16'h	b533;
47039	:douta	=	16'h	b513;
47040	:douta	=	16'h	a4d3;
47041	:douta	=	16'h	acf4;
47042	:douta	=	16'h	9cd4;
47043	:douta	=	16'h	9cb4;
47044	:douta	=	16'h	8c53;
47045	:douta	=	16'h	9cb4;
47046	:douta	=	16'h	8c73;
47047	:douta	=	16'h	8c73;
47048	:douta	=	16'h	8412;
47049	:douta	=	16'h	7c32;
47050	:douta	=	16'h	8c53;
47051	:douta	=	16'h	7bb0;
47052	:douta	=	16'h	83d1;
47053	:douta	=	16'h	7b8f;
47054	:douta	=	16'h	736d;
47055	:douta	=	16'h	51e6;
47056	:douta	=	16'h	49c4;
47057	:douta	=	16'h	41a5;
47058	:douta	=	16'h	41a5;
47059	:douta	=	16'h	5226;
47060	:douta	=	16'h	5a89;
47061	:douta	=	16'h	732c;
47062	:douta	=	16'h	734b;
47063	:douta	=	16'h	62c9;
47064	:douta	=	16'h	6b0b;
47065	:douta	=	16'h	6b0a;
47066	:douta	=	16'h	83cd;
47067	:douta	=	16'h	83cd;
47068	:douta	=	16'h	8bee;
47069	:douta	=	16'h	942e;
47070	:douta	=	16'h	944f;
47071	:douta	=	16'h	9c4f;
47072	:douta	=	16'h	acf2;
47073	:douta	=	16'h	7b8e;
47074	:douta	=	16'h	5acc;
47075	:douta	=	16'h	2967;
47076	:douta	=	16'h	1104;
47077	:douta	=	16'h	10e3;
47078	:douta	=	16'h	10c3;
47079	:douta	=	16'h	0883;
47080	:douta	=	16'h	39a7;
47081	:douta	=	16'h	0042;
47082	:douta	=	16'h	1084;
47083	:douta	=	16'h	2126;
47084	:douta	=	16'h	2947;
47085	:douta	=	16'h	5249;
47086	:douta	=	16'h	51a5;
47087	:douta	=	16'h	51c6;
47088	:douta	=	16'h	49a6;
47089	:douta	=	16'h	49a6;
47090	:douta	=	16'h	49a6;
47091	:douta	=	16'h	4986;
47092	:douta	=	16'h	4986;
47093	:douta	=	16'h	49a6;
47094	:douta	=	16'h	49a6;
47095	:douta	=	16'h	4185;
47096	:douta	=	16'h	4185;
47097	:douta	=	16'h	4185;
47098	:douta	=	16'h	4185;
47099	:douta	=	16'h	4186;
47100	:douta	=	16'h	4166;
47101	:douta	=	16'h	4186;
47102	:douta	=	16'h	4165;
47103	:douta	=	16'h	4186;
47104	:douta	=	16'h	ffbd;
47105	:douta	=	16'h	f75a;
47106	:douta	=	16'h	d5b5;
47107	:douta	=	16'h	e678;
47108	:douta	=	16'h	c5b6;
47109	:douta	=	16'h	a4b4;
47110	:douta	=	16'h	a4b3;
47111	:douta	=	16'h	b535;
47112	:douta	=	16'h	b535;
47113	:douta	=	16'h	c595;
47114	:douta	=	16'h	bd75;
47115	:douta	=	16'h	bd55;
47116	:douta	=	16'h	ad56;
47117	:douta	=	16'h	9493;
47118	:douta	=	16'h	94b5;
47119	:douta	=	16'h	8c74;
47120	:douta	=	16'h	8c95;
47121	:douta	=	16'h	8c74;
47122	:douta	=	16'h	8474;
47123	:douta	=	16'h	8454;
47124	:douta	=	16'h	8474;
47125	:douta	=	16'h	8454;
47126	:douta	=	16'h	8c75;
47127	:douta	=	16'h	4acd;
47128	:douta	=	16'h	20a3;
47129	:douta	=	16'h	20c3;
47130	:douta	=	16'h	20c3;
47131	:douta	=	16'h	20a3;
47132	:douta	=	16'h	20c2;
47133	:douta	=	16'h	20e3;
47134	:douta	=	16'h	18a2;
47135	:douta	=	16'h	1882;
47136	:douta	=	16'h	1882;
47137	:douta	=	16'h	1882;
47138	:douta	=	16'h	1882;
47139	:douta	=	16'h	1881;
47140	:douta	=	16'h	2082;
47141	:douta	=	16'h	1881;
47142	:douta	=	16'h	20a2;
47143	:douta	=	16'h	20a2;
47144	:douta	=	16'h	2082;
47145	:douta	=	16'h	20c2;
47146	:douta	=	16'h	20a2;
47147	:douta	=	16'h	28c2;
47148	:douta	=	16'h	28e2;
47149	:douta	=	16'h	28e2;
47150	:douta	=	16'h	30e3;
47151	:douta	=	16'h	28e2;
47152	:douta	=	16'h	30e2;
47153	:douta	=	16'h	3166;
47154	:douta	=	16'h	31c9;
47155	:douta	=	16'h	18c5;
47156	:douta	=	16'h	28e3;
47157	:douta	=	16'h	4143;
47158	:douta	=	16'h	4963;
47159	:douta	=	16'h	4963;
47160	:douta	=	16'h	4964;
47161	:douta	=	16'h	4983;
47162	:douta	=	16'h	51a4;
47163	:douta	=	16'h	51a4;
47164	:douta	=	16'h	59c4;
47165	:douta	=	16'h	59a4;
47166	:douta	=	16'h	734d;
47167	:douta	=	16'h	836a;
47168	:douta	=	16'h	6a04;
47169	:douta	=	16'h	61e4;
47170	:douta	=	16'h	4984;
47171	:douta	=	16'h	59c4;
47172	:douta	=	16'h	7224;
47173	:douta	=	16'h	7224;
47174	:douta	=	16'h	7224;
47175	:douta	=	16'h	7244;
47176	:douta	=	16'h	7244;
47177	:douta	=	16'h	7a44;
47178	:douta	=	16'h	7a44;
47179	:douta	=	16'h	7a44;
47180	:douta	=	16'h	7a64;
47181	:douta	=	16'h	7a64;
47182	:douta	=	16'h	8284;
47183	:douta	=	16'h	82a5;
47184	:douta	=	16'h	8aa4;
47185	:douta	=	16'h	8ac4;
47186	:douta	=	16'h	8ac5;
47187	:douta	=	16'h	9305;
47188	:douta	=	16'h	9b05;
47189	:douta	=	16'h	9b05;
47190	:douta	=	16'h	9b45;
47191	:douta	=	16'h	9b25;
47192	:douta	=	16'h	a365;
47193	:douta	=	16'h	ab85;
47194	:douta	=	16'h	ab65;
47195	:douta	=	16'h	ab85;
47196	:douta	=	16'h	aba5;
47197	:douta	=	16'h	b3a5;
47198	:douta	=	16'h	b385;
47199	:douta	=	16'h	b3a5;
47200	:douta	=	16'h	bbc6;
47201	:douta	=	16'h	bbc5;
47202	:douta	=	16'h	bbe6;
47203	:douta	=	16'h	bbe6;
47204	:douta	=	16'h	bbe6;
47205	:douta	=	16'h	bc06;
47206	:douta	=	16'h	bbe5;
47207	:douta	=	16'h	c406;
47208	:douta	=	16'h	c406;
47209	:douta	=	16'h	c406;
47210	:douta	=	16'h	c426;
47211	:douta	=	16'h	c406;
47212	:douta	=	16'h	c426;
47213	:douta	=	16'h	c426;
47214	:douta	=	16'h	c426;
47215	:douta	=	16'h	cc26;
47216	:douta	=	16'h	c426;
47217	:douta	=	16'h	cc26;
47218	:douta	=	16'h	cc26;
47219	:douta	=	16'h	cc26;
47220	:douta	=	16'h	cc46;
47221	:douta	=	16'h	c426;
47222	:douta	=	16'h	cc47;
47223	:douta	=	16'h	cc47;
47224	:douta	=	16'h	cc46;
47225	:douta	=	16'h	cc46;
47226	:douta	=	16'h	cc46;
47227	:douta	=	16'h	cc46;
47228	:douta	=	16'h	cc47;
47229	:douta	=	16'h	cc46;
47230	:douta	=	16'h	cc47;
47231	:douta	=	16'h	cc47;
47232	:douta	=	16'h	cc46;
47233	:douta	=	16'h	d467;
47234	:douta	=	16'h	cc47;
47235	:douta	=	16'h	cc47;
47236	:douta	=	16'h	cc67;
47237	:douta	=	16'h	cc67;
47238	:douta	=	16'h	d467;
47239	:douta	=	16'h	cc47;
47240	:douta	=	16'h	d467;
47241	:douta	=	16'h	d467;
47242	:douta	=	16'h	d467;
47243	:douta	=	16'h	d467;
47244	:douta	=	16'h	cc67;
47245	:douta	=	16'h	d467;
47246	:douta	=	16'h	d467;
47247	:douta	=	16'h	d467;
47248	:douta	=	16'h	d468;
47249	:douta	=	16'h	d467;
47250	:douta	=	16'h	d487;
47251	:douta	=	16'h	d487;
47252	:douta	=	16'h	d467;
47253	:douta	=	16'h	d467;
47254	:douta	=	16'h	d467;
47255	:douta	=	16'h	d487;
47256	:douta	=	16'h	d487;
47257	:douta	=	16'h	d467;
47258	:douta	=	16'h	d467;
47259	:douta	=	16'h	d467;
47260	:douta	=	16'h	d488;
47261	:douta	=	16'h	d487;
47262	:douta	=	16'h	d467;
47263	:douta	=	16'h	d487;
47264	:douta	=	16'h	d488;
47265	:douta	=	16'h	d467;
47266	:douta	=	16'h	d468;
47267	:douta	=	16'h	bcce;
47268	:douta	=	16'h	ce77;
47269	:douta	=	16'h	cc45;
47270	:douta	=	16'h	d487;
47271	:douta	=	16'h	d489;
47272	:douta	=	16'h	ac2b;
47273	:douta	=	16'h	a4d3;
47274	:douta	=	16'h	836d;
47275	:douta	=	16'h	bd53;
47276	:douta	=	16'h	838d;
47277	:douta	=	16'h	cdb3;
47278	:douta	=	16'h	bd72;
47279	:douta	=	16'h	cdb4;
47280	:douta	=	16'h	de36;
47281	:douta	=	16'h	c594;
47282	:douta	=	16'h	ad11;
47283	:douta	=	16'h	e636;
47284	:douta	=	16'h	d5f5;
47285	:douta	=	16'h	de56;
47286	:douta	=	16'h	d5d5;
47287	:douta	=	16'h	cd73;
47288	:douta	=	16'h	d5d4;
47289	:douta	=	16'h	cd73;
47290	:douta	=	16'h	c533;
47291	:douta	=	16'h	acf3;
47292	:douta	=	16'h	acd3;
47293	:douta	=	16'h	a4d3;
47294	:douta	=	16'h	acd3;
47295	:douta	=	16'h	acf3;
47296	:douta	=	16'h	a4d3;
47297	:douta	=	16'h	a4d3;
47298	:douta	=	16'h	8c74;
47299	:douta	=	16'h	8c73;
47300	:douta	=	16'h	7c12;
47301	:douta	=	16'h	9494;
47302	:douta	=	16'h	83f2;
47303	:douta	=	16'h	8412;
47304	:douta	=	16'h	8412;
47305	:douta	=	16'h	73b1;
47306	:douta	=	16'h	8411;
47307	:douta	=	16'h	6aeb;
47308	:douta	=	16'h	6b0c;
47309	:douta	=	16'h	49c5;
47310	:douta	=	16'h	3984;
47311	:douta	=	16'h	28e2;
47312	:douta	=	16'h	5a87;
47313	:douta	=	16'h	5a88;
47314	:douta	=	16'h	62a9;
47315	:douta	=	16'h	628a;
47316	:douta	=	16'h	62ca;
47317	:douta	=	16'h	7bcd;
47318	:douta	=	16'h	7b8c;
47319	:douta	=	16'h	736c;
47320	:douta	=	16'h	7b8c;
47321	:douta	=	16'h	7b8d;
47322	:douta	=	16'h	940e;
47323	:douta	=	16'h	9c4e;
47324	:douta	=	16'h	942f;
47325	:douta	=	16'h	9c6f;
47326	:douta	=	16'h	a490;
47327	:douta	=	16'h	a490;
47328	:douta	=	16'h	acd1;
47329	:douta	=	16'h	8bf0;
47330	:douta	=	16'h	6b2e;
47331	:douta	=	16'h	4a8b;
47332	:douta	=	16'h	2127;
47333	:douta	=	16'h	2126;
47334	:douta	=	16'h	1905;
47335	:douta	=	16'h	10e3;
47336	:douta	=	16'h	18c4;
47337	:douta	=	16'h	10c4;
47338	:douta	=	16'h	18c4;
47339	:douta	=	16'h	0882;
47340	:douta	=	16'h	18e5;
47341	:douta	=	16'h	41e9;
47342	:douta	=	16'h	4965;
47343	:douta	=	16'h	51c6;
47344	:douta	=	16'h	49a6;
47345	:douta	=	16'h	49a6;
47346	:douta	=	16'h	49a5;
47347	:douta	=	16'h	49a6;
47348	:douta	=	16'h	49a6;
47349	:douta	=	16'h	49a6;
47350	:douta	=	16'h	49a6;
47351	:douta	=	16'h	4186;
47352	:douta	=	16'h	4186;
47353	:douta	=	16'h	4185;
47354	:douta	=	16'h	4165;
47355	:douta	=	16'h	4165;
47356	:douta	=	16'h	4145;
47357	:douta	=	16'h	3924;
47358	:douta	=	16'h	3903;
47359	:douta	=	16'h	30e3;
47360	:douta	=	16'h	fffd;
47361	:douta	=	16'h	d5d5;
47362	:douta	=	16'h	d5d5;
47363	:douta	=	16'h	e677;
47364	:douta	=	16'h	acf4;
47365	:douta	=	16'h	a4b3;
47366	:douta	=	16'h	ad14;
47367	:douta	=	16'h	b556;
47368	:douta	=	16'h	cdb6;
47369	:douta	=	16'h	c595;
47370	:douta	=	16'h	bd75;
47371	:douta	=	16'h	b556;
47372	:douta	=	16'h	9cb4;
47373	:douta	=	16'h	9494;
47374	:douta	=	16'h	9495;
47375	:douta	=	16'h	94b5;
47376	:douta	=	16'h	8c94;
47377	:douta	=	16'h	8c74;
47378	:douta	=	16'h	8454;
47379	:douta	=	16'h	8454;
47380	:douta	=	16'h	8c95;
47381	:douta	=	16'h	8454;
47382	:douta	=	16'h	9d58;
47383	:douta	=	16'h	1020;
47384	:douta	=	16'h	20e3;
47385	:douta	=	16'h	20c3;
47386	:douta	=	16'h	20c3;
47387	:douta	=	16'h	20a3;
47388	:douta	=	16'h	18c3;
47389	:douta	=	16'h	20e3;
47390	:douta	=	16'h	1882;
47391	:douta	=	16'h	1882;
47392	:douta	=	16'h	1882;
47393	:douta	=	16'h	1882;
47394	:douta	=	16'h	2082;
47395	:douta	=	16'h	20a2;
47396	:douta	=	16'h	1881;
47397	:douta	=	16'h	1881;
47398	:douta	=	16'h	20a2;
47399	:douta	=	16'h	20a2;
47400	:douta	=	16'h	20a2;
47401	:douta	=	16'h	20a2;
47402	:douta	=	16'h	20a2;
47403	:douta	=	16'h	28e2;
47404	:douta	=	16'h	28e2;
47405	:douta	=	16'h	28e2;
47406	:douta	=	16'h	30e2;
47407	:douta	=	16'h	30e2;
47408	:douta	=	16'h	3103;
47409	:douta	=	16'h	39a8;
47410	:douta	=	16'h	31a8;
47411	:douta	=	16'h	18c5;
47412	:douta	=	16'h	3903;
47413	:douta	=	16'h	4143;
47414	:douta	=	16'h	4963;
47415	:douta	=	16'h	4963;
47416	:douta	=	16'h	5184;
47417	:douta	=	16'h	5184;
47418	:douta	=	16'h	5184;
47419	:douta	=	16'h	59c4;
47420	:douta	=	16'h	59c4;
47421	:douta	=	16'h	6206;
47422	:douta	=	16'h	8430;
47423	:douta	=	16'h	72a7;
47424	:douta	=	16'h	6a04;
47425	:douta	=	16'h	6a24;
47426	:douta	=	16'h	4163;
47427	:douta	=	16'h	59a4;
47428	:douta	=	16'h	7244;
47429	:douta	=	16'h	7244;
47430	:douta	=	16'h	7244;
47431	:douta	=	16'h	7a64;
47432	:douta	=	16'h	7a64;
47433	:douta	=	16'h	7a64;
47434	:douta	=	16'h	7a44;
47435	:douta	=	16'h	7a44;
47436	:douta	=	16'h	7a64;
47437	:douta	=	16'h	7a84;
47438	:douta	=	16'h	8284;
47439	:douta	=	16'h	82a4;
47440	:douta	=	16'h	8aa4;
47441	:douta	=	16'h	8ae5;
47442	:douta	=	16'h	92e5;
47443	:douta	=	16'h	9304;
47444	:douta	=	16'h	9b05;
47445	:douta	=	16'h	9b05;
47446	:douta	=	16'h	a345;
47447	:douta	=	16'h	a345;
47448	:douta	=	16'h	a345;
47449	:douta	=	16'h	ab65;
47450	:douta	=	16'h	ab65;
47451	:douta	=	16'h	b385;
47452	:douta	=	16'h	b385;
47453	:douta	=	16'h	b3a5;
47454	:douta	=	16'h	bbc6;
47455	:douta	=	16'h	bbc6;
47456	:douta	=	16'h	bbc6;
47457	:douta	=	16'h	bbe6;
47458	:douta	=	16'h	bbe6;
47459	:douta	=	16'h	bbe6;
47460	:douta	=	16'h	bbe6;
47461	:douta	=	16'h	c406;
47462	:douta	=	16'h	bbe5;
47463	:douta	=	16'h	c406;
47464	:douta	=	16'h	c406;
47465	:douta	=	16'h	c406;
47466	:douta	=	16'h	c426;
47467	:douta	=	16'h	c426;
47468	:douta	=	16'h	c426;
47469	:douta	=	16'h	c426;
47470	:douta	=	16'h	c426;
47471	:douta	=	16'h	c426;
47472	:douta	=	16'h	c426;
47473	:douta	=	16'h	cc26;
47474	:douta	=	16'h	cc26;
47475	:douta	=	16'h	cc47;
47476	:douta	=	16'h	cc46;
47477	:douta	=	16'h	cc47;
47478	:douta	=	16'h	cc47;
47479	:douta	=	16'h	cc47;
47480	:douta	=	16'h	cc46;
47481	:douta	=	16'h	cc46;
47482	:douta	=	16'h	cc46;
47483	:douta	=	16'h	cc46;
47484	:douta	=	16'h	cc46;
47485	:douta	=	16'h	cc46;
47486	:douta	=	16'h	cc47;
47487	:douta	=	16'h	cc46;
47488	:douta	=	16'h	cc47;
47489	:douta	=	16'h	d467;
47490	:douta	=	16'h	cc46;
47491	:douta	=	16'h	cc47;
47492	:douta	=	16'h	cc47;
47493	:douta	=	16'h	cc67;
47494	:douta	=	16'h	d467;
47495	:douta	=	16'h	d467;
47496	:douta	=	16'h	d467;
47497	:douta	=	16'h	d467;
47498	:douta	=	16'h	d467;
47499	:douta	=	16'h	d467;
47500	:douta	=	16'h	d467;
47501	:douta	=	16'h	d467;
47502	:douta	=	16'h	d467;
47503	:douta	=	16'h	d467;
47504	:douta	=	16'h	d467;
47505	:douta	=	16'h	d467;
47506	:douta	=	16'h	d467;
47507	:douta	=	16'h	d467;
47508	:douta	=	16'h	d467;
47509	:douta	=	16'h	d467;
47510	:douta	=	16'h	d467;
47511	:douta	=	16'h	d467;
47512	:douta	=	16'h	d487;
47513	:douta	=	16'h	d487;
47514	:douta	=	16'h	d487;
47515	:douta	=	16'h	d467;
47516	:douta	=	16'h	d487;
47517	:douta	=	16'h	d487;
47518	:douta	=	16'h	d488;
47519	:douta	=	16'h	d468;
47520	:douta	=	16'h	d468;
47521	:douta	=	16'h	d488;
47522	:douta	=	16'h	d467;
47523	:douta	=	16'h	b4ce;
47524	:douta	=	16'h	ce76;
47525	:douta	=	16'h	cc45;
47526	:douta	=	16'h	d488;
47527	:douta	=	16'h	d487;
47528	:douta	=	16'h	dc87;
47529	:douta	=	16'h	abec;
47530	:douta	=	16'h	b512;
47531	:douta	=	16'h	acd0;
47532	:douta	=	16'h	b512;
47533	:douta	=	16'h	cdd4;
47534	:douta	=	16'h	c593;
47535	:douta	=	16'h	d615;
47536	:douta	=	16'h	de57;
47537	:douta	=	16'h	b513;
47538	:douta	=	16'h	de57;
47539	:douta	=	16'h	de36;
47540	:douta	=	16'h	cdb5;
47541	:douta	=	16'h	cdb5;
47542	:douta	=	16'h	d616;
47543	:douta	=	16'h	acf3;
47544	:douta	=	16'h	b514;
47545	:douta	=	16'h	a4b2;
47546	:douta	=	16'h	9c93;
47547	:douta	=	16'h	9c93;
47548	:douta	=	16'h	9c73;
47549	:douta	=	16'h	9c94;
47550	:douta	=	16'h	8c32;
47551	:douta	=	16'h	8c11;
47552	:douta	=	16'h	9473;
47553	:douta	=	16'h	9452;
47554	:douta	=	16'h	7bd0;
47555	:douta	=	16'h	8412;
47556	:douta	=	16'h	7bf2;
47557	:douta	=	16'h	7390;
47558	:douta	=	16'h	83d0;
47559	:douta	=	16'h	62aa;
47560	:douta	=	16'h	3965;
47561	:douta	=	16'h	3944;
47562	:douta	=	16'h	3103;
47563	:douta	=	16'h	41a5;
47564	:douta	=	16'h	49e6;
47565	:douta	=	16'h	6ac9;
47566	:douta	=	16'h	62a9;
47567	:douta	=	16'h	5a88;
47568	:douta	=	16'h	6ae9;
47569	:douta	=	16'h	732a;
47570	:douta	=	16'h	7b8c;
47571	:douta	=	16'h	7b8c;
47572	:douta	=	16'h	83cd;
47573	:douta	=	16'h	9c6f;
47574	:douta	=	16'h	a490;
47575	:douta	=	16'h	acf0;
47576	:douta	=	16'h	b511;
47577	:douta	=	16'h	b4f0;
47578	:douta	=	16'h	b4f0;
47579	:douta	=	16'h	b511;
47580	:douta	=	16'h	b511;
47581	:douta	=	16'h	b511;
47582	:douta	=	16'h	bd31;
47583	:douta	=	16'h	acd1;
47584	:douta	=	16'h	acd1;
47585	:douta	=	16'h	8c30;
47586	:douta	=	16'h	7bd0;
47587	:douta	=	16'h	6b6f;
47588	:douta	=	16'h	52ed;
47589	:douta	=	16'h	424b;
47590	:douta	=	16'h	2968;
47591	:douta	=	16'h	2967;
47592	:douta	=	16'h	1906;
47593	:douta	=	16'h	31c9;
47594	:douta	=	16'h	18e5;
47595	:douta	=	16'h	2988;
47596	:douta	=	16'h	10c5;
47597	:douta	=	16'h	0863;
47598	:douta	=	16'h	72a9;
47599	:douta	=	16'h	51a5;
47600	:douta	=	16'h	4985;
47601	:douta	=	16'h	4965;
47602	:douta	=	16'h	4124;
47603	:douta	=	16'h	4124;
47604	:douta	=	16'h	3944;
47605	:douta	=	16'h	4165;
47606	:douta	=	16'h	41a6;
47607	:douta	=	16'h	5208;
47608	:douta	=	16'h	5aab;
47609	:douta	=	16'h	630c;
47610	:douta	=	16'h	6b8f;
47611	:douta	=	16'h	73d1;
47612	:douta	=	16'h	7c53;
47613	:douta	=	16'h	84b5;
47614	:douta	=	16'h	84b4;
47615	:douta	=	16'h	84b4;
47616	:douta	=	16'h	ffdd;
47617	:douta	=	16'h	d5b5;
47618	:douta	=	16'h	d5f6;
47619	:douta	=	16'h	e677;
47620	:douta	=	16'h	9cb3;
47621	:douta	=	16'h	a4b3;
47622	:douta	=	16'h	b535;
47623	:douta	=	16'h	ad15;
47624	:douta	=	16'h	cdf6;
47625	:douta	=	16'h	bd95;
47626	:douta	=	16'h	b555;
47627	:douta	=	16'h	ad35;
47628	:douta	=	16'h	9494;
47629	:douta	=	16'h	8c74;
47630	:douta	=	16'h	8c94;
47631	:douta	=	16'h	94b5;
47632	:douta	=	16'h	8c95;
47633	:douta	=	16'h	8c74;
47634	:douta	=	16'h	8454;
47635	:douta	=	16'h	8c74;
47636	:douta	=	16'h	8c74;
47637	:douta	=	16'h	8c95;
47638	:douta	=	16'h	9517;
47639	:douta	=	16'h	1040;
47640	:douta	=	16'h	20c3;
47641	:douta	=	16'h	20c3;
47642	:douta	=	16'h	20a3;
47643	:douta	=	16'h	20a3;
47644	:douta	=	16'h	18c3;
47645	:douta	=	16'h	18c3;
47646	:douta	=	16'h	1882;
47647	:douta	=	16'h	1882;
47648	:douta	=	16'h	18a2;
47649	:douta	=	16'h	1882;
47650	:douta	=	16'h	1882;
47651	:douta	=	16'h	1882;
47652	:douta	=	16'h	20a2;
47653	:douta	=	16'h	1881;
47654	:douta	=	16'h	20a2;
47655	:douta	=	16'h	20a2;
47656	:douta	=	16'h	20a2;
47657	:douta	=	16'h	28e2;
47658	:douta	=	16'h	20a2;
47659	:douta	=	16'h	28e3;
47660	:douta	=	16'h	28e2;
47661	:douta	=	16'h	28e2;
47662	:douta	=	16'h	30e2;
47663	:douta	=	16'h	30e3;
47664	:douta	=	16'h	30e2;
47665	:douta	=	16'h	39c9;
47666	:douta	=	16'h	31a8;
47667	:douta	=	16'h	18a4;
47668	:douta	=	16'h	4123;
47669	:douta	=	16'h	4143;
47670	:douta	=	16'h	4963;
47671	:douta	=	16'h	4984;
47672	:douta	=	16'h	4963;
47673	:douta	=	16'h	5184;
47674	:douta	=	16'h	59a4;
47675	:douta	=	16'h	59c4;
47676	:douta	=	16'h	59c4;
47677	:douta	=	16'h	6267;
47678	:douta	=	16'h	94b2;
47679	:douta	=	16'h	6a44;
47680	:douta	=	16'h	6a04;
47681	:douta	=	16'h	6a24;
47682	:douta	=	16'h	4143;
47683	:douta	=	16'h	61c4;
47684	:douta	=	16'h	7224;
47685	:douta	=	16'h	7244;
47686	:douta	=	16'h	7a44;
47687	:douta	=	16'h	7a64;
47688	:douta	=	16'h	7a84;
47689	:douta	=	16'h	7a64;
47690	:douta	=	16'h	7a64;
47691	:douta	=	16'h	7a44;
47692	:douta	=	16'h	7a64;
47693	:douta	=	16'h	8284;
47694	:douta	=	16'h	82a4;
47695	:douta	=	16'h	82a4;
47696	:douta	=	16'h	8aa4;
47697	:douta	=	16'h	8ae4;
47698	:douta	=	16'h	92e5;
47699	:douta	=	16'h	9304;
47700	:douta	=	16'h	9b05;
47701	:douta	=	16'h	9b25;
47702	:douta	=	16'h	9b45;
47703	:douta	=	16'h	a345;
47704	:douta	=	16'h	a365;
47705	:douta	=	16'h	ab85;
47706	:douta	=	16'h	ab85;
47707	:douta	=	16'h	b385;
47708	:douta	=	16'h	b385;
47709	:douta	=	16'h	b3a5;
47710	:douta	=	16'h	b3a5;
47711	:douta	=	16'h	bbc6;
47712	:douta	=	16'h	bbc6;
47713	:douta	=	16'h	bbe6;
47714	:douta	=	16'h	bbe6;
47715	:douta	=	16'h	bbc6;
47716	:douta	=	16'h	bbe6;
47717	:douta	=	16'h	c406;
47718	:douta	=	16'h	bc06;
47719	:douta	=	16'h	c406;
47720	:douta	=	16'h	c406;
47721	:douta	=	16'h	c406;
47722	:douta	=	16'h	c426;
47723	:douta	=	16'h	c426;
47724	:douta	=	16'h	c426;
47725	:douta	=	16'h	c426;
47726	:douta	=	16'h	c426;
47727	:douta	=	16'h	cc26;
47728	:douta	=	16'h	cc46;
47729	:douta	=	16'h	cc46;
47730	:douta	=	16'h	cc47;
47731	:douta	=	16'h	cc47;
47732	:douta	=	16'h	c426;
47733	:douta	=	16'h	cc47;
47734	:douta	=	16'h	cc47;
47735	:douta	=	16'h	cc46;
47736	:douta	=	16'h	cc46;
47737	:douta	=	16'h	cc46;
47738	:douta	=	16'h	cc46;
47739	:douta	=	16'h	cc46;
47740	:douta	=	16'h	cc46;
47741	:douta	=	16'h	cc46;
47742	:douta	=	16'h	cc46;
47743	:douta	=	16'h	cc46;
47744	:douta	=	16'h	cc47;
47745	:douta	=	16'h	cc47;
47746	:douta	=	16'h	cc46;
47747	:douta	=	16'h	cc47;
47748	:douta	=	16'h	cc46;
47749	:douta	=	16'h	cc67;
47750	:douta	=	16'h	d467;
47751	:douta	=	16'h	d467;
47752	:douta	=	16'h	d467;
47753	:douta	=	16'h	d467;
47754	:douta	=	16'h	d467;
47755	:douta	=	16'h	d467;
47756	:douta	=	16'h	d467;
47757	:douta	=	16'h	d467;
47758	:douta	=	16'h	d467;
47759	:douta	=	16'h	cc67;
47760	:douta	=	16'h	d467;
47761	:douta	=	16'h	d487;
47762	:douta	=	16'h	d487;
47763	:douta	=	16'h	d487;
47764	:douta	=	16'h	d487;
47765	:douta	=	16'h	cc67;
47766	:douta	=	16'h	d467;
47767	:douta	=	16'h	d467;
47768	:douta	=	16'h	d467;
47769	:douta	=	16'h	d487;
47770	:douta	=	16'h	d487;
47771	:douta	=	16'h	d467;
47772	:douta	=	16'h	d487;
47773	:douta	=	16'h	d467;
47774	:douta	=	16'h	d468;
47775	:douta	=	16'h	d488;
47776	:douta	=	16'h	d488;
47777	:douta	=	16'h	d487;
47778	:douta	=	16'h	d466;
47779	:douta	=	16'h	b4ce;
47780	:douta	=	16'h	ce76;
47781	:douta	=	16'h	cc45;
47782	:douta	=	16'h	d468;
47783	:douta	=	16'h	cc87;
47784	:douta	=	16'h	e486;
47785	:douta	=	16'h	abcb;
47786	:douta	=	16'h	acd1;
47787	:douta	=	16'h	acd1;
47788	:douta	=	16'h	b511;
47789	:douta	=	16'h	cdd4;
47790	:douta	=	16'h	c573;
47791	:douta	=	16'h	de37;
47792	:douta	=	16'h	d616;
47793	:douta	=	16'h	b513;
47794	:douta	=	16'h	de57;
47795	:douta	=	16'h	cdd5;
47796	:douta	=	16'h	c596;
47797	:douta	=	16'h	bd75;
47798	:douta	=	16'h	bd75;
47799	:douta	=	16'h	acf3;
47800	:douta	=	16'h	9c93;
47801	:douta	=	16'h	9c93;
47802	:douta	=	16'h	9452;
47803	:douta	=	16'h	9473;
47804	:douta	=	16'h	9473;
47805	:douta	=	16'h	9473;
47806	:douta	=	16'h	8c12;
47807	:douta	=	16'h	83f1;
47808	:douta	=	16'h	7bb0;
47809	:douta	=	16'h	8c33;
47810	:douta	=	16'h	7390;
47811	:douta	=	16'h	7bd0;
47812	:douta	=	16'h	738e;
47813	:douta	=	16'h	39a6;
47814	:douta	=	16'h	41a6;
47815	:douta	=	16'h	49a5;
47816	:douta	=	16'h	3944;
47817	:douta	=	16'h	3984;
47818	:douta	=	16'h	5227;
47819	:douta	=	16'h	5a88;
47820	:douta	=	16'h	6288;
47821	:douta	=	16'h	7b6b;
47822	:douta	=	16'h	7b6b;
47823	:douta	=	16'h	6aea;
47824	:douta	=	16'h	732a;
47825	:douta	=	16'h	7b6c;
47826	:douta	=	16'h	83cd;
47827	:douta	=	16'h	8c0d;
47828	:douta	=	16'h	9c4f;
47829	:douta	=	16'h	a4af;
47830	:douta	=	16'h	acf0;
47831	:douta	=	16'h	bd31;
47832	:douta	=	16'h	bd31;
47833	:douta	=	16'h	c551;
47834	:douta	=	16'h	c551;
47835	:douta	=	16'h	c572;
47836	:douta	=	16'h	c572;
47837	:douta	=	16'h	c552;
47838	:douta	=	16'h	bd52;
47839	:douta	=	16'h	b4d1;
47840	:douta	=	16'h	a4b1;
47841	:douta	=	16'h	8c30;
47842	:douta	=	16'h	83f0;
47843	:douta	=	16'h	6b6f;
47844	:douta	=	16'h	5b0e;
47845	:douta	=	16'h	52ac;
47846	:douta	=	16'h	39e9;
47847	:douta	=	16'h	31a8;
47848	:douta	=	16'h	2126;
47849	:douta	=	16'h	31c8;
47850	:douta	=	16'h	2106;
47851	:douta	=	16'h	2968;
47852	:douta	=	16'h	2988;
47853	:douta	=	16'h	0883;
47854	:douta	=	16'h	832c;
47855	:douta	=	16'h	51a5;
47856	:douta	=	16'h	4a07;
47857	:douta	=	16'h	5228;
47858	:douta	=	16'h	5aab;
47859	:douta	=	16'h	6b4e;
47860	:douta	=	16'h	6b6f;
47861	:douta	=	16'h	73f1;
47862	:douta	=	16'h	7432;
47863	:douta	=	16'h	7c73;
47864	:douta	=	16'h	7c73;
47865	:douta	=	16'h	7c94;
47866	:douta	=	16'h	7c73;
47867	:douta	=	16'h	7452;
47868	:douta	=	16'h	6bd0;
47869	:douta	=	16'h	636e;
47870	:douta	=	16'h	5b2d;
47871	:douta	=	16'h	52cb;
47872	:douta	=	16'h	f6f9;
47873	:douta	=	16'h	cdb5;
47874	:douta	=	16'h	de37;
47875	:douta	=	16'h	de37;
47876	:douta	=	16'h	a4b3;
47877	:douta	=	16'h	a4d3;
47878	:douta	=	16'h	acf5;
47879	:douta	=	16'h	b514;
47880	:douta	=	16'h	cdb5;
47881	:douta	=	16'h	b535;
47882	:douta	=	16'h	b555;
47883	:douta	=	16'h	9494;
47884	:douta	=	16'h	9cb4;
47885	:douta	=	16'h	9474;
47886	:douta	=	16'h	8c94;
47887	:douta	=	16'h	94b5;
47888	:douta	=	16'h	8c95;
47889	:douta	=	16'h	8c74;
47890	:douta	=	16'h	8433;
47891	:douta	=	16'h	8c95;
47892	:douta	=	16'h	8475;
47893	:douta	=	16'h	9d38;
47894	:douta	=	16'h	3a4a;
47895	:douta	=	16'h	20c3;
47896	:douta	=	16'h	20c3;
47897	:douta	=	16'h	20c3;
47898	:douta	=	16'h	20c3;
47899	:douta	=	16'h	20c3;
47900	:douta	=	16'h	18a3;
47901	:douta	=	16'h	18c3;
47902	:douta	=	16'h	1882;
47903	:douta	=	16'h	1882;
47904	:douta	=	16'h	1882;
47905	:douta	=	16'h	1882;
47906	:douta	=	16'h	2082;
47907	:douta	=	16'h	2082;
47908	:douta	=	16'h	20a2;
47909	:douta	=	16'h	20a2;
47910	:douta	=	16'h	20a2;
47911	:douta	=	16'h	2082;
47912	:douta	=	16'h	20a2;
47913	:douta	=	16'h	20c2;
47914	:douta	=	16'h	28c2;
47915	:douta	=	16'h	28e2;
47916	:douta	=	16'h	28c2;
47917	:douta	=	16'h	28c2;
47918	:douta	=	16'h	30e3;
47919	:douta	=	16'h	30e3;
47920	:douta	=	16'h	30e2;
47921	:douta	=	16'h	39e9;
47922	:douta	=	16'h	2967;
47923	:douta	=	16'h	28e4;
47924	:douta	=	16'h	4943;
47925	:douta	=	16'h	4143;
47926	:douta	=	16'h	4963;
47927	:douta	=	16'h	4963;
47928	:douta	=	16'h	5184;
47929	:douta	=	16'h	5184;
47930	:douta	=	16'h	51a3;
47931	:douta	=	16'h	59a4;
47932	:douta	=	16'h	61c4;
47933	:douta	=	16'h	6b0a;
47934	:douta	=	16'h	a555;
47935	:douta	=	16'h	61a3;
47936	:douta	=	16'h	6a24;
47937	:douta	=	16'h	6a24;
47938	:douta	=	16'h	4164;
47939	:douta	=	16'h	51a4;
47940	:douta	=	16'h	7244;
47941	:douta	=	16'h	7a64;
47942	:douta	=	16'h	7a44;
47943	:douta	=	16'h	7a64;
47944	:douta	=	16'h	7a64;
47945	:douta	=	16'h	7a44;
47946	:douta	=	16'h	7a64;
47947	:douta	=	16'h	7a84;
47948	:douta	=	16'h	7a64;
47949	:douta	=	16'h	8284;
47950	:douta	=	16'h	82a4;
47951	:douta	=	16'h	8ac5;
47952	:douta	=	16'h	8ac4;
47953	:douta	=	16'h	8ae4;
47954	:douta	=	16'h	92e5;
47955	:douta	=	16'h	9305;
47956	:douta	=	16'h	9b25;
47957	:douta	=	16'h	9b26;
47958	:douta	=	16'h	a346;
47959	:douta	=	16'h	a345;
47960	:douta	=	16'h	a365;
47961	:douta	=	16'h	ab65;
47962	:douta	=	16'h	ab65;
47963	:douta	=	16'h	b3a5;
47964	:douta	=	16'h	b3a5;
47965	:douta	=	16'h	b3a5;
47966	:douta	=	16'h	b3a5;
47967	:douta	=	16'h	bbc5;
47968	:douta	=	16'h	bbc5;
47969	:douta	=	16'h	bbe6;
47970	:douta	=	16'h	bbc6;
47971	:douta	=	16'h	bbe6;
47972	:douta	=	16'h	bc06;
47973	:douta	=	16'h	c406;
47974	:douta	=	16'h	c406;
47975	:douta	=	16'h	c406;
47976	:douta	=	16'h	c406;
47977	:douta	=	16'h	c426;
47978	:douta	=	16'h	c426;
47979	:douta	=	16'h	c426;
47980	:douta	=	16'h	c426;
47981	:douta	=	16'h	c426;
47982	:douta	=	16'h	c426;
47983	:douta	=	16'h	cc26;
47984	:douta	=	16'h	cc46;
47985	:douta	=	16'h	c426;
47986	:douta	=	16'h	cc26;
47987	:douta	=	16'h	cc46;
47988	:douta	=	16'h	cc46;
47989	:douta	=	16'h	cc46;
47990	:douta	=	16'h	cc26;
47991	:douta	=	16'h	cc46;
47992	:douta	=	16'h	cc46;
47993	:douta	=	16'h	cc46;
47994	:douta	=	16'h	cc46;
47995	:douta	=	16'h	cc46;
47996	:douta	=	16'h	cc46;
47997	:douta	=	16'h	cc67;
47998	:douta	=	16'h	cc46;
47999	:douta	=	16'h	cc47;
48000	:douta	=	16'h	cc46;
48001	:douta	=	16'h	cc67;
48002	:douta	=	16'h	cc47;
48003	:douta	=	16'h	cc46;
48004	:douta	=	16'h	cc47;
48005	:douta	=	16'h	d467;
48006	:douta	=	16'h	d467;
48007	:douta	=	16'h	d467;
48008	:douta	=	16'h	d467;
48009	:douta	=	16'h	d467;
48010	:douta	=	16'h	d467;
48011	:douta	=	16'h	cc67;
48012	:douta	=	16'h	d467;
48013	:douta	=	16'h	d467;
48014	:douta	=	16'h	cc47;
48015	:douta	=	16'h	d468;
48016	:douta	=	16'h	d468;
48017	:douta	=	16'h	d487;
48018	:douta	=	16'h	d487;
48019	:douta	=	16'h	d467;
48020	:douta	=	16'h	d487;
48021	:douta	=	16'h	d487;
48022	:douta	=	16'h	d467;
48023	:douta	=	16'h	d467;
48024	:douta	=	16'h	d487;
48025	:douta	=	16'h	d467;
48026	:douta	=	16'h	d487;
48027	:douta	=	16'h	d487;
48028	:douta	=	16'h	d467;
48029	:douta	=	16'h	d467;
48030	:douta	=	16'h	d487;
48031	:douta	=	16'h	d488;
48032	:douta	=	16'h	d488;
48033	:douta	=	16'h	d487;
48034	:douta	=	16'h	d467;
48035	:douta	=	16'h	b4ce;
48036	:douta	=	16'h	ce76;
48037	:douta	=	16'h	cc45;
48038	:douta	=	16'h	d488;
48039	:douta	=	16'h	d487;
48040	:douta	=	16'h	d467;
48041	:douta	=	16'h	cc87;
48042	:douta	=	16'h	944f;
48043	:douta	=	16'h	a4b1;
48044	:douta	=	16'h	acd1;
48045	:douta	=	16'h	c553;
48046	:douta	=	16'h	c594;
48047	:douta	=	16'h	cdf5;
48048	:douta	=	16'h	c5b5;
48049	:douta	=	16'h	bd54;
48050	:douta	=	16'h	c5b6;
48051	:douta	=	16'h	bd96;
48052	:douta	=	16'h	b556;
48053	:douta	=	16'h	b556;
48054	:douta	=	16'h	a4f5;
48055	:douta	=	16'h	9493;
48056	:douta	=	16'h	9c94;
48057	:douta	=	16'h	8411;
48058	:douta	=	16'h	7bf1;
48059	:douta	=	16'h	83f1;
48060	:douta	=	16'h	83f0;
48061	:douta	=	16'h	7bb0;
48062	:douta	=	16'h	7bd0;
48063	:douta	=	16'h	83f0;
48064	:douta	=	16'h	734d;
48065	:douta	=	16'h	5248;
48066	:douta	=	16'h	4a27;
48067	:douta	=	16'h	2903;
48068	:douta	=	16'h	3123;
48069	:douta	=	16'h	6aea;
48070	:douta	=	16'h	732b;
48071	:douta	=	16'h	62ca;
48072	:douta	=	16'h	6aea;
48073	:douta	=	16'h	732a;
48074	:douta	=	16'h	730a;
48075	:douta	=	16'h	730a;
48076	:douta	=	16'h	732a;
48077	:douta	=	16'h	8bcc;
48078	:douta	=	16'h	8bee;
48079	:douta	=	16'h	8c0e;
48080	:douta	=	16'h	942e;
48081	:douta	=	16'h	944f;
48082	:douta	=	16'h	9c8f;
48083	:douta	=	16'h	9c6f;
48084	:douta	=	16'h	a4af;
48085	:douta	=	16'h	b510;
48086	:douta	=	16'h	bd51;
48087	:douta	=	16'h	c572;
48088	:douta	=	16'h	c572;
48089	:douta	=	16'h	cd92;
48090	:douta	=	16'h	cdb3;
48091	:douta	=	16'h	d5d4;
48092	:douta	=	16'h	cdb3;
48093	:douta	=	16'h	cd93;
48094	:douta	=	16'h	c573;
48095	:douta	=	16'h	acd2;
48096	:douta	=	16'h	a4b1;
48097	:douta	=	16'h	8c10;
48098	:douta	=	16'h	8410;
48099	:douta	=	16'h	632e;
48100	:douta	=	16'h	5aec;
48101	:douta	=	16'h	52cd;
48102	:douta	=	16'h	4aad;
48103	:douta	=	16'h	426c;
48104	:douta	=	16'h	31c9;
48105	:douta	=	16'h	2106;
48106	:douta	=	16'h	2126;
48107	:douta	=	16'h	1905;
48108	:douta	=	16'h	2126;
48109	:douta	=	16'h	2127;
48110	:douta	=	16'h	0062;
48111	:douta	=	16'h	10e5;
48112	:douta	=	16'h	52ab;
48113	:douta	=	16'h	8471;
48114	:douta	=	16'h	6b6e;
48115	:douta	=	16'h	632c;
48116	:douta	=	16'h	5acb;
48117	:douta	=	16'h	52aa;
48118	:douta	=	16'h	5289;
48119	:douta	=	16'h	5228;
48120	:douta	=	16'h	49e7;
48121	:douta	=	16'h	49c6;
48122	:douta	=	16'h	49a5;
48123	:douta	=	16'h	4985;
48124	:douta	=	16'h	4965;
48125	:douta	=	16'h	4985;
48126	:douta	=	16'h	4985;
48127	:douta	=	16'h	5185;
48128	:douta	=	16'h	e697;
48129	:douta	=	16'h	d5b5;
48130	:douta	=	16'h	de77;
48131	:douta	=	16'h	cdd6;
48132	:douta	=	16'h	a4d4;
48133	:douta	=	16'h	a4b3;
48134	:douta	=	16'h	acf5;
48135	:douta	=	16'h	c595;
48136	:douta	=	16'h	c595;
48137	:douta	=	16'h	b535;
48138	:douta	=	16'h	b555;
48139	:douta	=	16'h	9453;
48140	:douta	=	16'h	9cd5;
48141	:douta	=	16'h	9494;
48142	:douta	=	16'h	8c74;
48143	:douta	=	16'h	94b5;
48144	:douta	=	16'h	8c74;
48145	:douta	=	16'h	8c74;
48146	:douta	=	16'h	8433;
48147	:douta	=	16'h	8475;
48148	:douta	=	16'h	8c74;
48149	:douta	=	16'h	7c33;
48150	:douta	=	16'h	18a2;
48151	:douta	=	16'h	20c3;
48152	:douta	=	16'h	20c3;
48153	:douta	=	16'h	20a2;
48154	:douta	=	16'h	20c3;
48155	:douta	=	16'h	20c3;
48156	:douta	=	16'h	18a3;
48157	:douta	=	16'h	18a3;
48158	:douta	=	16'h	1882;
48159	:douta	=	16'h	1882;
48160	:douta	=	16'h	1882;
48161	:douta	=	16'h	1882;
48162	:douta	=	16'h	2082;
48163	:douta	=	16'h	2082;
48164	:douta	=	16'h	20a2;
48165	:douta	=	16'h	2082;
48166	:douta	=	16'h	20a2;
48167	:douta	=	16'h	20a2;
48168	:douta	=	16'h	20c2;
48169	:douta	=	16'h	28c2;
48170	:douta	=	16'h	20c2;
48171	:douta	=	16'h	20c2;
48172	:douta	=	16'h	28e2;
48173	:douta	=	16'h	30e2;
48174	:douta	=	16'h	30e3;
48175	:douta	=	16'h	3103;
48176	:douta	=	16'h	3103;
48177	:douta	=	16'h	31c9;
48178	:douta	=	16'h	2947;
48179	:douta	=	16'h	3103;
48180	:douta	=	16'h	4963;
48181	:douta	=	16'h	4963;
48182	:douta	=	16'h	4963;
48183	:douta	=	16'h	4963;
48184	:douta	=	16'h	5184;
48185	:douta	=	16'h	59a4;
48186	:douta	=	16'h	51a4;
48187	:douta	=	16'h	59c4;
48188	:douta	=	16'h	61c4;
48189	:douta	=	16'h	734c;
48190	:douta	=	16'h	ad74;
48191	:douta	=	16'h	61a3;
48192	:douta	=	16'h	6a04;
48193	:douta	=	16'h	6a24;
48194	:douta	=	16'h	4964;
48195	:douta	=	16'h	5184;
48196	:douta	=	16'h	7224;
48197	:douta	=	16'h	7a64;
48198	:douta	=	16'h	7a44;
48199	:douta	=	16'h	7a64;
48200	:douta	=	16'h	7a85;
48201	:douta	=	16'h	7a64;
48202	:douta	=	16'h	7a44;
48203	:douta	=	16'h	7a64;
48204	:douta	=	16'h	7a64;
48205	:douta	=	16'h	8284;
48206	:douta	=	16'h	82a4;
48207	:douta	=	16'h	8ac4;
48208	:douta	=	16'h	8ac4;
48209	:douta	=	16'h	8ae4;
48210	:douta	=	16'h	92e5;
48211	:douta	=	16'h	9305;
48212	:douta	=	16'h	9b26;
48213	:douta	=	16'h	9b26;
48214	:douta	=	16'h	a346;
48215	:douta	=	16'h	a345;
48216	:douta	=	16'h	ab65;
48217	:douta	=	16'h	ab65;
48218	:douta	=	16'h	ab85;
48219	:douta	=	16'h	b3a5;
48220	:douta	=	16'h	b3a5;
48221	:douta	=	16'h	b3a6;
48222	:douta	=	16'h	b3a6;
48223	:douta	=	16'h	bbc5;
48224	:douta	=	16'h	bbc5;
48225	:douta	=	16'h	bbe6;
48226	:douta	=	16'h	bbe6;
48227	:douta	=	16'h	bbe6;
48228	:douta	=	16'h	bbe5;
48229	:douta	=	16'h	c406;
48230	:douta	=	16'h	c406;
48231	:douta	=	16'h	c406;
48232	:douta	=	16'h	c406;
48233	:douta	=	16'h	c426;
48234	:douta	=	16'h	c426;
48235	:douta	=	16'h	c426;
48236	:douta	=	16'h	c426;
48237	:douta	=	16'h	c426;
48238	:douta	=	16'h	cc26;
48239	:douta	=	16'h	cc26;
48240	:douta	=	16'h	cc46;
48241	:douta	=	16'h	cc46;
48242	:douta	=	16'h	cc26;
48243	:douta	=	16'h	cc47;
48244	:douta	=	16'h	cc26;
48245	:douta	=	16'h	cc46;
48246	:douta	=	16'h	cc46;
48247	:douta	=	16'h	cc46;
48248	:douta	=	16'h	cc46;
48249	:douta	=	16'h	cc46;
48250	:douta	=	16'h	cc46;
48251	:douta	=	16'h	cc46;
48252	:douta	=	16'h	cc46;
48253	:douta	=	16'h	cc46;
48254	:douta	=	16'h	cc46;
48255	:douta	=	16'h	cc46;
48256	:douta	=	16'h	cc67;
48257	:douta	=	16'h	cc47;
48258	:douta	=	16'h	cc47;
48259	:douta	=	16'h	cc47;
48260	:douta	=	16'h	cc67;
48261	:douta	=	16'h	d467;
48262	:douta	=	16'h	d467;
48263	:douta	=	16'h	d467;
48264	:douta	=	16'h	d467;
48265	:douta	=	16'h	d467;
48266	:douta	=	16'h	d467;
48267	:douta	=	16'h	d467;
48268	:douta	=	16'h	cc67;
48269	:douta	=	16'h	d487;
48270	:douta	=	16'h	d467;
48271	:douta	=	16'h	d468;
48272	:douta	=	16'h	d488;
48273	:douta	=	16'h	d467;
48274	:douta	=	16'h	d487;
48275	:douta	=	16'h	d467;
48276	:douta	=	16'h	d467;
48277	:douta	=	16'h	d467;
48278	:douta	=	16'h	d467;
48279	:douta	=	16'h	d487;
48280	:douta	=	16'h	d487;
48281	:douta	=	16'h	d468;
48282	:douta	=	16'h	d467;
48283	:douta	=	16'h	d487;
48284	:douta	=	16'h	d467;
48285	:douta	=	16'h	d487;
48286	:douta	=	16'h	d468;
48287	:douta	=	16'h	d488;
48288	:douta	=	16'h	d488;
48289	:douta	=	16'h	d467;
48290	:douta	=	16'h	d467;
48291	:douta	=	16'h	b4ce;
48292	:douta	=	16'h	ce56;
48293	:douta	=	16'h	cc25;
48294	:douta	=	16'h	d488;
48295	:douta	=	16'h	d487;
48296	:douta	=	16'h	d487;
48297	:douta	=	16'h	d485;
48298	:douta	=	16'h	9430;
48299	:douta	=	16'h	a491;
48300	:douta	=	16'h	a472;
48301	:douta	=	16'h	b4f3;
48302	:douta	=	16'h	c553;
48303	:douta	=	16'h	c5b5;
48304	:douta	=	16'h	c595;
48305	:douta	=	16'h	bd54;
48306	:douta	=	16'h	b575;
48307	:douta	=	16'h	ad36;
48308	:douta	=	16'h	ad56;
48309	:douta	=	16'h	9cf5;
48310	:douta	=	16'h	9cd4;
48311	:douta	=	16'h	8433;
48312	:douta	=	16'h	8433;
48313	:douta	=	16'h	7bd1;
48314	:douta	=	16'h	7b90;
48315	:douta	=	16'h	83d0;
48316	:douta	=	16'h	7b8f;
48317	:douta	=	16'h	7b8f;
48318	:douta	=	16'h	7b6e;
48319	:douta	=	16'h	6aeb;
48320	:douta	=	16'h	49e5;
48321	:douta	=	16'h	3944;
48322	:douta	=	16'h	4185;
48323	:douta	=	16'h	5247;
48324	:douta	=	16'h	5a88;
48325	:douta	=	16'h	6288;
48326	:douta	=	16'h	9c6f;
48327	:douta	=	16'h	838c;
48328	:douta	=	16'h	730b;
48329	:douta	=	16'h	7b4b;
48330	:douta	=	16'h	7b4b;
48331	:douta	=	16'h	836b;
48332	:douta	=	16'h	834b;
48333	:douta	=	16'h	8bac;
48334	:douta	=	16'h	940e;
48335	:douta	=	16'h	9c6f;
48336	:douta	=	16'h	acd0;
48337	:douta	=	16'h	acd0;
48338	:douta	=	16'h	acd0;
48339	:douta	=	16'h	acaf;
48340	:douta	=	16'h	b510;
48341	:douta	=	16'h	cd92;
48342	:douta	=	16'h	cdb3;
48343	:douta	=	16'h	cdb3;
48344	:douta	=	16'h	cdb3;
48345	:douta	=	16'h	d5d4;
48346	:douta	=	16'h	cdb4;
48347	:douta	=	16'h	cdd4;
48348	:douta	=	16'h	cdb3;
48349	:douta	=	16'h	c573;
48350	:douta	=	16'h	cd93;
48351	:douta	=	16'h	b512;
48352	:douta	=	16'h	acd2;
48353	:douta	=	16'h	9431;
48354	:douta	=	16'h	8c30;
48355	:douta	=	16'h	6b6f;
48356	:douta	=	16'h	5b0d;
48357	:douta	=	16'h	5aed;
48358	:douta	=	16'h	52cd;
48359	:douta	=	16'h	4a8d;
48360	:douta	=	16'h	3a4c;
48361	:douta	=	16'h	2126;
48362	:douta	=	16'h	2967;
48363	:douta	=	16'h	10a4;
48364	:douta	=	16'h	1905;
48365	:douta	=	16'h	2147;
48366	:douta	=	16'h	1083;
48367	:douta	=	16'h	18e5;
48368	:douta	=	16'h	2925;
48369	:douta	=	16'h	5a89;
48370	:douta	=	16'h	5226;
48371	:douta	=	16'h	49c6;
48372	:douta	=	16'h	49a5;
48373	:douta	=	16'h	49a5;
48374	:douta	=	16'h	4985;
48375	:douta	=	16'h	4985;
48376	:douta	=	16'h	4985;
48377	:douta	=	16'h	4985;
48378	:douta	=	16'h	4985;
48379	:douta	=	16'h	49a5;
48380	:douta	=	16'h	51a5;
48381	:douta	=	16'h	51a5;
48382	:douta	=	16'h	51c5;
48383	:douta	=	16'h	49a5;
48384	:douta	=	16'h	d615;
48385	:douta	=	16'h	de37;
48386	:douta	=	16'h	ee98;
48387	:douta	=	16'h	ad14;
48388	:douta	=	16'h	a4b3;
48389	:douta	=	16'h	acf4;
48390	:douta	=	16'h	bd54;
48391	:douta	=	16'h	d5f6;
48392	:douta	=	16'h	bd75;
48393	:douta	=	16'h	b555;
48394	:douta	=	16'h	ad16;
48395	:douta	=	16'h	9c73;
48396	:douta	=	16'h	9cb5;
48397	:douta	=	16'h	94b5;
48398	:douta	=	16'h	8c94;
48399	:douta	=	16'h	94b5;
48400	:douta	=	16'h	9495;
48401	:douta	=	16'h	8454;
48402	:douta	=	16'h	8454;
48403	:douta	=	16'h	8c95;
48404	:douta	=	16'h	94f7;
48405	:douta	=	16'h	2124;
48406	:douta	=	16'h	1861;
48407	:douta	=	16'h	20a3;
48408	:douta	=	16'h	20c3;
48409	:douta	=	16'h	20c3;
48410	:douta	=	16'h	20a3;
48411	:douta	=	16'h	20c3;
48412	:douta	=	16'h	20c3;
48413	:douta	=	16'h	1882;
48414	:douta	=	16'h	1882;
48415	:douta	=	16'h	1882;
48416	:douta	=	16'h	1882;
48417	:douta	=	16'h	1861;
48418	:douta	=	16'h	20a2;
48419	:douta	=	16'h	20a2;
48420	:douta	=	16'h	20a2;
48421	:douta	=	16'h	20a2;
48422	:douta	=	16'h	20a2;
48423	:douta	=	16'h	20a2;
48424	:douta	=	16'h	20c2;
48425	:douta	=	16'h	20c2;
48426	:douta	=	16'h	28c2;
48427	:douta	=	16'h	28e2;
48428	:douta	=	16'h	3103;
48429	:douta	=	16'h	30e2;
48430	:douta	=	16'h	3103;
48431	:douta	=	16'h	3103;
48432	:douta	=	16'h	3944;
48433	:douta	=	16'h	31a8;
48434	:douta	=	16'h	1906;
48435	:douta	=	16'h	3944;
48436	:douta	=	16'h	4963;
48437	:douta	=	16'h	4963;
48438	:douta	=	16'h	4963;
48439	:douta	=	16'h	4984;
48440	:douta	=	16'h	5184;
48441	:douta	=	16'h	5184;
48442	:douta	=	16'h	59a4;
48443	:douta	=	16'h	61c4;
48444	:douta	=	16'h	59a3;
48445	:douta	=	16'h	8c50;
48446	:douta	=	16'h	ad12;
48447	:douta	=	16'h	69e3;
48448	:douta	=	16'h	6a24;
48449	:douta	=	16'h	6a24;
48450	:douta	=	16'h	6a24;
48451	:douta	=	16'h	4164;
48452	:douta	=	16'h	7a64;
48453	:douta	=	16'h	7244;
48454	:douta	=	16'h	7a64;
48455	:douta	=	16'h	7a84;
48456	:douta	=	16'h	7a84;
48457	:douta	=	16'h	7a64;
48458	:douta	=	16'h	7a84;
48459	:douta	=	16'h	7a64;
48460	:douta	=	16'h	8284;
48461	:douta	=	16'h	8285;
48462	:douta	=	16'h	82a4;
48463	:douta	=	16'h	8aa4;
48464	:douta	=	16'h	8ac5;
48465	:douta	=	16'h	8ae4;
48466	:douta	=	16'h	92e5;
48467	:douta	=	16'h	9b25;
48468	:douta	=	16'h	a326;
48469	:douta	=	16'h	a346;
48470	:douta	=	16'h	a346;
48471	:douta	=	16'h	a345;
48472	:douta	=	16'h	ab65;
48473	:douta	=	16'h	ab85;
48474	:douta	=	16'h	b385;
48475	:douta	=	16'h	b3a5;
48476	:douta	=	16'h	b3a6;
48477	:douta	=	16'h	b3a6;
48478	:douta	=	16'h	b3a6;
48479	:douta	=	16'h	bbc5;
48480	:douta	=	16'h	bbe6;
48481	:douta	=	16'h	bbe6;
48482	:douta	=	16'h	bbe6;
48483	:douta	=	16'h	bbe6;
48484	:douta	=	16'h	bbe6;
48485	:douta	=	16'h	c406;
48486	:douta	=	16'h	bc06;
48487	:douta	=	16'h	c406;
48488	:douta	=	16'h	c406;
48489	:douta	=	16'h	c405;
48490	:douta	=	16'h	c426;
48491	:douta	=	16'h	c426;
48492	:douta	=	16'h	c426;
48493	:douta	=	16'h	c426;
48494	:douta	=	16'h	c425;
48495	:douta	=	16'h	c426;
48496	:douta	=	16'h	cc26;
48497	:douta	=	16'h	cc26;
48498	:douta	=	16'h	c425;
48499	:douta	=	16'h	cc47;
48500	:douta	=	16'h	cc46;
48501	:douta	=	16'h	cc46;
48502	:douta	=	16'h	cc46;
48503	:douta	=	16'h	cc45;
48504	:douta	=	16'h	cc46;
48505	:douta	=	16'h	cc46;
48506	:douta	=	16'h	cc46;
48507	:douta	=	16'h	cc47;
48508	:douta	=	16'h	cc46;
48509	:douta	=	16'h	cc47;
48510	:douta	=	16'h	cc67;
48511	:douta	=	16'h	cc67;
48512	:douta	=	16'h	cc46;
48513	:douta	=	16'h	cc47;
48514	:douta	=	16'h	cc47;
48515	:douta	=	16'h	d467;
48516	:douta	=	16'h	cc67;
48517	:douta	=	16'h	d467;
48518	:douta	=	16'h	d467;
48519	:douta	=	16'h	d467;
48520	:douta	=	16'h	d467;
48521	:douta	=	16'h	d467;
48522	:douta	=	16'h	d467;
48523	:douta	=	16'h	cc67;
48524	:douta	=	16'h	d467;
48525	:douta	=	16'h	d467;
48526	:douta	=	16'h	d467;
48527	:douta	=	16'h	d468;
48528	:douta	=	16'h	d488;
48529	:douta	=	16'h	d467;
48530	:douta	=	16'h	d467;
48531	:douta	=	16'h	d467;
48532	:douta	=	16'h	d467;
48533	:douta	=	16'h	d467;
48534	:douta	=	16'h	d467;
48535	:douta	=	16'h	d467;
48536	:douta	=	16'h	d467;
48537	:douta	=	16'h	d488;
48538	:douta	=	16'h	d488;
48539	:douta	=	16'h	d488;
48540	:douta	=	16'h	d488;
48541	:douta	=	16'h	d488;
48542	:douta	=	16'h	d488;
48543	:douta	=	16'h	d467;
48544	:douta	=	16'h	cc87;
48545	:douta	=	16'h	d488;
48546	:douta	=	16'h	d487;
48547	:douta	=	16'h	b4ee;
48548	:douta	=	16'h	ce77;
48549	:douta	=	16'h	cc25;
48550	:douta	=	16'h	d467;
48551	:douta	=	16'h	d488;
48552	:douta	=	16'h	cc87;
48553	:douta	=	16'h	d487;
48554	:douta	=	16'h	ac4d;
48555	:douta	=	16'h	9430;
48556	:douta	=	16'h	a4b2;
48557	:douta	=	16'h	9c92;
48558	:douta	=	16'h	9c93;
48559	:douta	=	16'h	ad15;
48560	:douta	=	16'h	b535;
48561	:douta	=	16'h	b515;
48562	:douta	=	16'h	9494;
48563	:douta	=	16'h	9493;
48564	:douta	=	16'h	8c73;
48565	:douta	=	16'h	8c53;
48566	:douta	=	16'h	7bd1;
48567	:douta	=	16'h	73b0;
48568	:douta	=	16'h	73b0;
48569	:douta	=	16'h	736f;
48570	:douta	=	16'h	8412;
48571	:douta	=	16'h	6acc;
48572	:douta	=	16'h	49c5;
48573	:douta	=	16'h	3964;
48574	:douta	=	16'h	4185;
48575	:douta	=	16'h	62a9;
48576	:douta	=	16'h	62c9;
48577	:douta	=	16'h	62c9;
48578	:douta	=	16'h	6b0a;
48579	:douta	=	16'h	6b2a;
48580	:douta	=	16'h	6b4a;
48581	:douta	=	16'h	5a68;
48582	:douta	=	16'h	acd0;
48583	:douta	=	16'h	a4b0;
48584	:douta	=	16'h	9c2e;
48585	:douta	=	16'h	940e;
48586	:douta	=	16'h	940e;
48587	:douta	=	16'h	93ed;
48588	:douta	=	16'h	940e;
48589	:douta	=	16'h	9c4e;
48590	:douta	=	16'h	a48e;
48591	:douta	=	16'h	b4f0;
48592	:douta	=	16'h	c551;
48593	:douta	=	16'h	c551;
48594	:douta	=	16'h	c572;
48595	:douta	=	16'h	cd93;
48596	:douta	=	16'h	d5d4;
48597	:douta	=	16'h	d5f4;
48598	:douta	=	16'h	d5f4;
48599	:douta	=	16'h	d5d4;
48600	:douta	=	16'h	d5f5;
48601	:douta	=	16'h	d5f4;
48602	:douta	=	16'h	cdd4;
48603	:douta	=	16'h	cdd4;
48604	:douta	=	16'h	cdb4;
48605	:douta	=	16'h	cd93;
48606	:douta	=	16'h	c573;
48607	:douta	=	16'h	bd53;
48608	:douta	=	16'h	b513;
48609	:douta	=	16'h	9c51;
48610	:douta	=	16'h	8c31;
48611	:douta	=	16'h	83f0;
48612	:douta	=	16'h	630e;
48613	:douta	=	16'h	52ed;
48614	:douta	=	16'h	5b2f;
48615	:douta	=	16'h	52ee;
48616	:douta	=	16'h	4ace;
48617	:douta	=	16'h	31c9;
48618	:douta	=	16'h	528b;
48619	:douta	=	16'h	10c3;
48620	:douta	=	16'h	20e5;
48621	:douta	=	16'h	2126;
48622	:douta	=	16'h	2126;
48623	:douta	=	16'h	08a4;
48624	:douta	=	16'h	10e5;
48625	:douta	=	16'h	2904;
48626	:douta	=	16'h	51c5;
48627	:douta	=	16'h	51a6;
48628	:douta	=	16'h	51c5;
48629	:douta	=	16'h	49a5;
48630	:douta	=	16'h	49a5;
48631	:douta	=	16'h	49a5;
48632	:douta	=	16'h	51c6;
48633	:douta	=	16'h	51c6;
48634	:douta	=	16'h	49a5;
48635	:douta	=	16'h	51c6;
48636	:douta	=	16'h	51c6;
48637	:douta	=	16'h	59c6;
48638	:douta	=	16'h	51c6;
48639	:douta	=	16'h	51c5;
48640	:douta	=	16'h	cdb5;
48641	:douta	=	16'h	e677;
48642	:douta	=	16'h	e677;
48643	:douta	=	16'h	acd4;
48644	:douta	=	16'h	a4b3;
48645	:douta	=	16'h	ad15;
48646	:douta	=	16'h	cdd5;
48647	:douta	=	16'h	d5d6;
48648	:douta	=	16'h	b555;
48649	:douta	=	16'h	b536;
48650	:douta	=	16'h	a4f5;
48651	:douta	=	16'h	9c94;
48652	:douta	=	16'h	9493;
48653	:douta	=	16'h	94b5;
48654	:douta	=	16'h	8c94;
48655	:douta	=	16'h	9495;
48656	:douta	=	16'h	8c94;
48657	:douta	=	16'h	8434;
48658	:douta	=	16'h	8454;
48659	:douta	=	16'h	8c95;
48660	:douta	=	16'h	a558;
48661	:douta	=	16'h	1020;
48662	:douta	=	16'h	20c3;
48663	:douta	=	16'h	20a3;
48664	:douta	=	16'h	20c3;
48665	:douta	=	16'h	20a3;
48666	:douta	=	16'h	20c3;
48667	:douta	=	16'h	18c3;
48668	:douta	=	16'h	20c3;
48669	:douta	=	16'h	1882;
48670	:douta	=	16'h	1882;
48671	:douta	=	16'h	1881;
48672	:douta	=	16'h	1881;
48673	:douta	=	16'h	1882;
48674	:douta	=	16'h	20a2;
48675	:douta	=	16'h	20a2;
48676	:douta	=	16'h	20a2;
48677	:douta	=	16'h	20a2;
48678	:douta	=	16'h	20a2;
48679	:douta	=	16'h	20c2;
48680	:douta	=	16'h	20a2;
48681	:douta	=	16'h	28c2;
48682	:douta	=	16'h	28c2;
48683	:douta	=	16'h	28e2;
48684	:douta	=	16'h	30e3;
48685	:douta	=	16'h	3103;
48686	:douta	=	16'h	3103;
48687	:douta	=	16'h	3903;
48688	:douta	=	16'h	3144;
48689	:douta	=	16'h	3188;
48690	:douta	=	16'h	1905;
48691	:douta	=	16'h	4143;
48692	:douta	=	16'h	4963;
48693	:douta	=	16'h	4964;
48694	:douta	=	16'h	4983;
48695	:douta	=	16'h	51a4;
48696	:douta	=	16'h	5184;
48697	:douta	=	16'h	59a4;
48698	:douta	=	16'h	51a4;
48699	:douta	=	16'h	59c4;
48700	:douta	=	16'h	5983;
48701	:douta	=	16'h	94d3;
48702	:douta	=	16'h	9cb0;
48703	:douta	=	16'h	6a03;
48704	:douta	=	16'h	6a24;
48705	:douta	=	16'h	6a24;
48706	:douta	=	16'h	7264;
48707	:douta	=	16'h	49a4;
48708	:douta	=	16'h	7a83;
48709	:douta	=	16'h	7a44;
48710	:douta	=	16'h	7a64;
48711	:douta	=	16'h	7a64;
48712	:douta	=	16'h	7a84;
48713	:douta	=	16'h	7a64;
48714	:douta	=	16'h	7a84;
48715	:douta	=	16'h	7a64;
48716	:douta	=	16'h	8284;
48717	:douta	=	16'h	8284;
48718	:douta	=	16'h	8284;
48719	:douta	=	16'h	8aa4;
48720	:douta	=	16'h	8ac5;
48721	:douta	=	16'h	8ac4;
48722	:douta	=	16'h	92e4;
48723	:douta	=	16'h	9325;
48724	:douta	=	16'h	9b45;
48725	:douta	=	16'h	9b45;
48726	:douta	=	16'h	a366;
48727	:douta	=	16'h	a345;
48728	:douta	=	16'h	ab65;
48729	:douta	=	16'h	ab65;
48730	:douta	=	16'h	b385;
48731	:douta	=	16'h	b3a6;
48732	:douta	=	16'h	b3a5;
48733	:douta	=	16'h	bbc6;
48734	:douta	=	16'h	b3a6;
48735	:douta	=	16'h	bbc5;
48736	:douta	=	16'h	bbe6;
48737	:douta	=	16'h	bbe6;
48738	:douta	=	16'h	bbe6;
48739	:douta	=	16'h	bbe6;
48740	:douta	=	16'h	bbe5;
48741	:douta	=	16'h	c406;
48742	:douta	=	16'h	c406;
48743	:douta	=	16'h	c407;
48744	:douta	=	16'h	c407;
48745	:douta	=	16'h	c405;
48746	:douta	=	16'h	c406;
48747	:douta	=	16'h	c426;
48748	:douta	=	16'h	c426;
48749	:douta	=	16'h	c446;
48750	:douta	=	16'h	c426;
48751	:douta	=	16'h	c426;
48752	:douta	=	16'h	c426;
48753	:douta	=	16'h	cc46;
48754	:douta	=	16'h	cc46;
48755	:douta	=	16'h	cc26;
48756	:douta	=	16'h	cc26;
48757	:douta	=	16'h	cc46;
48758	:douta	=	16'h	cc46;
48759	:douta	=	16'h	cc46;
48760	:douta	=	16'h	cc46;
48761	:douta	=	16'h	cc46;
48762	:douta	=	16'h	cc46;
48763	:douta	=	16'h	cc47;
48764	:douta	=	16'h	cc47;
48765	:douta	=	16'h	cc47;
48766	:douta	=	16'h	cc47;
48767	:douta	=	16'h	cc67;
48768	:douta	=	16'h	cc46;
48769	:douta	=	16'h	cc47;
48770	:douta	=	16'h	cc47;
48771	:douta	=	16'h	d467;
48772	:douta	=	16'h	cc47;
48773	:douta	=	16'h	d467;
48774	:douta	=	16'h	d467;
48775	:douta	=	16'h	cc67;
48776	:douta	=	16'h	d467;
48777	:douta	=	16'h	cc67;
48778	:douta	=	16'h	d468;
48779	:douta	=	16'h	d467;
48780	:douta	=	16'h	cc67;
48781	:douta	=	16'h	d488;
48782	:douta	=	16'h	d468;
48783	:douta	=	16'h	d487;
48784	:douta	=	16'h	d487;
48785	:douta	=	16'h	d468;
48786	:douta	=	16'h	d467;
48787	:douta	=	16'h	d487;
48788	:douta	=	16'h	d467;
48789	:douta	=	16'h	d467;
48790	:douta	=	16'h	d487;
48791	:douta	=	16'h	d467;
48792	:douta	=	16'h	d468;
48793	:douta	=	16'h	d468;
48794	:douta	=	16'h	d488;
48795	:douta	=	16'h	d488;
48796	:douta	=	16'h	d467;
48797	:douta	=	16'h	d467;
48798	:douta	=	16'h	d488;
48799	:douta	=	16'h	cc68;
48800	:douta	=	16'h	d468;
48801	:douta	=	16'h	d487;
48802	:douta	=	16'h	d487;
48803	:douta	=	16'h	b4ce;
48804	:douta	=	16'h	ce76;
48805	:douta	=	16'h	cc25;
48806	:douta	=	16'h	d468;
48807	:douta	=	16'h	d488;
48808	:douta	=	16'h	cc87;
48809	:douta	=	16'h	cc88;
48810	:douta	=	16'h	cc69;
48811	:douta	=	16'h	942f;
48812	:douta	=	16'h	9c92;
48813	:douta	=	16'h	9c72;
48814	:douta	=	16'h	9c93;
48815	:douta	=	16'h	9473;
48816	:douta	=	16'h	9c93;
48817	:douta	=	16'h	a4d4;
48818	:douta	=	16'h	8432;
48819	:douta	=	16'h	8c53;
48820	:douta	=	16'h	8c32;
48821	:douta	=	16'h	8411;
48822	:douta	=	16'h	7bd2;
48823	:douta	=	16'h	736e;
48824	:douta	=	16'h	736f;
48825	:douta	=	16'h	6aeb;
48826	:douta	=	16'h	6aeb;
48827	:douta	=	16'h	3984;
48828	:douta	=	16'h	3944;
48829	:douta	=	16'h	3984;
48830	:douta	=	16'h	734c;
48831	:douta	=	16'h	734b;
48832	:douta	=	16'h	6b0a;
48833	:douta	=	16'h	730a;
48834	:douta	=	16'h	732b;
48835	:douta	=	16'h	736b;
48836	:douta	=	16'h	7b8b;
48837	:douta	=	16'h	5ac9;
48838	:douta	=	16'h	8bed;
48839	:douta	=	16'h	acb0;
48840	:douta	=	16'h	a490;
48841	:douta	=	16'h	acaf;
48842	:douta	=	16'h	a48f;
48843	:douta	=	16'h	9c4e;
48844	:douta	=	16'h	a46e;
48845	:douta	=	16'h	ac8e;
48846	:douta	=	16'h	accf;
48847	:douta	=	16'h	bd31;
48848	:douta	=	16'h	c572;
48849	:douta	=	16'h	c552;
48850	:douta	=	16'h	cdb4;
48851	:douta	=	16'h	d5d4;
48852	:douta	=	16'h	d5f4;
48853	:douta	=	16'h	de35;
48854	:douta	=	16'h	de15;
48855	:douta	=	16'h	ddf4;
48856	:douta	=	16'h	d5d4;
48857	:douta	=	16'h	d5d4;
48858	:douta	=	16'h	c593;
48859	:douta	=	16'h	cd94;
48860	:douta	=	16'h	c573;
48861	:douta	=	16'h	c573;
48862	:douta	=	16'h	bd33;
48863	:douta	=	16'h	bd53;
48864	:douta	=	16'h	b513;
48865	:douta	=	16'h	9cb2;
48866	:douta	=	16'h	9472;
48867	:douta	=	16'h	8431;
48868	:douta	=	16'h	634e;
48869	:douta	=	16'h	52ac;
48870	:douta	=	16'h	4a6b;
48871	:douta	=	16'h	426b;
48872	:douta	=	16'h	3a4c;
48873	:douta	=	16'h	3a4c;
48874	:douta	=	16'h	62ec;
48875	:douta	=	16'h	0883;
48876	:douta	=	16'h	18c5;
48877	:douta	=	16'h	1905;
48878	:douta	=	16'h	2147;
48879	:douta	=	16'h	18e5;
48880	:douta	=	16'h	1946;
48881	:douta	=	16'h	18e5;
48882	:douta	=	16'h	59e6;
48883	:douta	=	16'h	51c6;
48884	:douta	=	16'h	51c5;
48885	:douta	=	16'h	51a5;
48886	:douta	=	16'h	51c6;
48887	:douta	=	16'h	51c6;
48888	:douta	=	16'h	51c6;
48889	:douta	=	16'h	51c6;
48890	:douta	=	16'h	51c5;
48891	:douta	=	16'h	51a6;
48892	:douta	=	16'h	51c6;
48893	:douta	=	16'h	51c6;
48894	:douta	=	16'h	51c6;
48895	:douta	=	16'h	59e6;
48896	:douta	=	16'h	bd12;
48897	:douta	=	16'h	e698;
48898	:douta	=	16'h	cdd6;
48899	:douta	=	16'h	b535;
48900	:douta	=	16'h	ad14;
48901	:douta	=	16'h	ad15;
48902	:douta	=	16'h	d616;
48903	:douta	=	16'h	c595;
48904	:douta	=	16'h	b554;
48905	:douta	=	16'h	a536;
48906	:douta	=	16'h	9494;
48907	:douta	=	16'h	9474;
48908	:douta	=	16'h	94b4;
48909	:douta	=	16'h	9494;
48910	:douta	=	16'h	94b5;
48911	:douta	=	16'h	9495;
48912	:douta	=	16'h	8474;
48913	:douta	=	16'h	8433;
48914	:douta	=	16'h	8c94;
48915	:douta	=	16'h	9d59;
48916	:douta	=	16'h	6b90;
48917	:douta	=	16'h	20a3;
48918	:douta	=	16'h	20c3;
48919	:douta	=	16'h	20a3;
48920	:douta	=	16'h	20c3;
48921	:douta	=	16'h	20c3;
48922	:douta	=	16'h	20c3;
48923	:douta	=	16'h	20c3;
48924	:douta	=	16'h	20e3;
48925	:douta	=	16'h	18a2;
48926	:douta	=	16'h	1881;
48927	:douta	=	16'h	20a2;
48928	:douta	=	16'h	18a2;
48929	:douta	=	16'h	20a2;
48930	:douta	=	16'h	20a2;
48931	:douta	=	16'h	20a2;
48932	:douta	=	16'h	20a2;
48933	:douta	=	16'h	20a2;
48934	:douta	=	16'h	2082;
48935	:douta	=	16'h	20c2;
48936	:douta	=	16'h	28e2;
48937	:douta	=	16'h	28c2;
48938	:douta	=	16'h	28c2;
48939	:douta	=	16'h	28e3;
48940	:douta	=	16'h	28e2;
48941	:douta	=	16'h	3103;
48942	:douta	=	16'h	3103;
48943	:douta	=	16'h	3103;
48944	:douta	=	16'h	3986;
48945	:douta	=	16'h	2967;
48946	:douta	=	16'h	10c5;
48947	:douta	=	16'h	4963;
48948	:douta	=	16'h	4963;
48949	:douta	=	16'h	4984;
48950	:douta	=	16'h	5184;
48951	:douta	=	16'h	5184;
48952	:douta	=	16'h	59a4;
48953	:douta	=	16'h	59a4;
48954	:douta	=	16'h	59c4;
48955	:douta	=	16'h	61e4;
48956	:douta	=	16'h	59a3;
48957	:douta	=	16'h	a573;
48958	:douta	=	16'h	940c;
48959	:douta	=	16'h	6a24;
48960	:douta	=	16'h	6a24;
48961	:douta	=	16'h	7224;
48962	:douta	=	16'h	7a64;
48963	:douta	=	16'h	6204;
48964	:douta	=	16'h	7a64;
48965	:douta	=	16'h	7a64;
48966	:douta	=	16'h	7a84;
48967	:douta	=	16'h	7a84;
48968	:douta	=	16'h	7a84;
48969	:douta	=	16'h	7a84;
48970	:douta	=	16'h	7a64;
48971	:douta	=	16'h	8285;
48972	:douta	=	16'h	7a64;
48973	:douta	=	16'h	82a4;
48974	:douta	=	16'h	82a5;
48975	:douta	=	16'h	8ac4;
48976	:douta	=	16'h	8ac5;
48977	:douta	=	16'h	8ac4;
48978	:douta	=	16'h	9305;
48979	:douta	=	16'h	9325;
48980	:douta	=	16'h	9b45;
48981	:douta	=	16'h	a325;
48982	:douta	=	16'h	a345;
48983	:douta	=	16'h	a345;
48984	:douta	=	16'h	ab65;
48985	:douta	=	16'h	ab85;
48986	:douta	=	16'h	b385;
48987	:douta	=	16'h	b3a6;
48988	:douta	=	16'h	b3a6;
48989	:douta	=	16'h	b3a6;
48990	:douta	=	16'h	bbc6;
48991	:douta	=	16'h	bbc6;
48992	:douta	=	16'h	bbe6;
48993	:douta	=	16'h	bc06;
48994	:douta	=	16'h	bbe6;
48995	:douta	=	16'h	bbe5;
48996	:douta	=	16'h	bc06;
48997	:douta	=	16'h	c406;
48998	:douta	=	16'h	c406;
48999	:douta	=	16'h	c405;
49000	:douta	=	16'h	c426;
49001	:douta	=	16'h	c426;
49002	:douta	=	16'h	c426;
49003	:douta	=	16'h	c426;
49004	:douta	=	16'h	c426;
49005	:douta	=	16'h	c426;
49006	:douta	=	16'h	c426;
49007	:douta	=	16'h	cc46;
49008	:douta	=	16'h	cc46;
49009	:douta	=	16'h	cc26;
49010	:douta	=	16'h	cc26;
49011	:douta	=	16'h	cc46;
49012	:douta	=	16'h	cc47;
49013	:douta	=	16'h	cc47;
49014	:douta	=	16'h	cc47;
49015	:douta	=	16'h	cc47;
49016	:douta	=	16'h	cc47;
49017	:douta	=	16'h	cc46;
49018	:douta	=	16'h	cc47;
49019	:douta	=	16'h	cc46;
49020	:douta	=	16'h	cc46;
49021	:douta	=	16'h	cc47;
49022	:douta	=	16'h	cc67;
49023	:douta	=	16'h	cc67;
49024	:douta	=	16'h	cc47;
49025	:douta	=	16'h	cc46;
49026	:douta	=	16'h	cc46;
49027	:douta	=	16'h	d467;
49028	:douta	=	16'h	d467;
49029	:douta	=	16'h	d467;
49030	:douta	=	16'h	d468;
49031	:douta	=	16'h	d467;
49032	:douta	=	16'h	d467;
49033	:douta	=	16'h	cc67;
49034	:douta	=	16'h	cc67;
49035	:douta	=	16'h	d467;
49036	:douta	=	16'h	d467;
49037	:douta	=	16'h	d468;
49038	:douta	=	16'h	cc67;
49039	:douta	=	16'h	d487;
49040	:douta	=	16'h	d467;
49041	:douta	=	16'h	d467;
49042	:douta	=	16'h	d487;
49043	:douta	=	16'h	d467;
49044	:douta	=	16'h	d467;
49045	:douta	=	16'h	d467;
49046	:douta	=	16'h	d467;
49047	:douta	=	16'h	d467;
49048	:douta	=	16'h	d487;
49049	:douta	=	16'h	d487;
49050	:douta	=	16'h	d487;
49051	:douta	=	16'h	d487;
49052	:douta	=	16'h	d488;
49053	:douta	=	16'h	d488;
49054	:douta	=	16'h	d488;
49055	:douta	=	16'h	d488;
49056	:douta	=	16'h	d487;
49057	:douta	=	16'h	cc68;
49058	:douta	=	16'h	d467;
49059	:douta	=	16'h	accd;
49060	:douta	=	16'h	d677;
49061	:douta	=	16'h	cc25;
49062	:douta	=	16'h	d467;
49063	:douta	=	16'h	cc68;
49064	:douta	=	16'h	d468;
49065	:douta	=	16'h	cc88;
49066	:douta	=	16'h	d485;
49067	:douta	=	16'h	c468;
49068	:douta	=	16'h	9430;
49069	:douta	=	16'h	9431;
49070	:douta	=	16'h	8bf1;
49071	:douta	=	16'h	83f1;
49072	:douta	=	16'h	83d1;
49073	:douta	=	16'h	7bb0;
49074	:douta	=	16'h	7bf1;
49075	:douta	=	16'h	738f;
49076	:douta	=	16'h	8c33;
49077	:douta	=	16'h	9432;
49078	:douta	=	16'h	4a26;
49079	:douta	=	16'h	49e6;
49080	:douta	=	16'h	3964;
49081	:douta	=	16'h	39a4;
49082	:douta	=	16'h	4a06;
49083	:douta	=	16'h	5a68;
49084	:douta	=	16'h	62aa;
49085	:douta	=	16'h	7b8d;
49086	:douta	=	16'h	8bcd;
49087	:douta	=	16'h	6b0a;
49088	:douta	=	16'h	838d;
49089	:douta	=	16'h	838c;
49090	:douta	=	16'h	83ad;
49091	:douta	=	16'h	83cd;
49092	:douta	=	16'h	93ee;
49093	:douta	=	16'h	a470;
49094	:douta	=	16'h	5268;
49095	:douta	=	16'h	942f;
49096	:douta	=	16'h	ac8f;
49097	:douta	=	16'h	bd10;
49098	:douta	=	16'h	b4d0;
49099	:douta	=	16'h	b4f0;
49100	:douta	=	16'h	bd51;
49101	:douta	=	16'h	c552;
49102	:douta	=	16'h	cd92;
49103	:douta	=	16'h	d5d3;
49104	:douta	=	16'h	cdb3;
49105	:douta	=	16'h	cdb3;
49106	:douta	=	16'h	cdd3;
49107	:douta	=	16'h	d615;
49108	:douta	=	16'h	d614;
49109	:douta	=	16'h	d5f4;
49110	:douta	=	16'h	d5f4;
49111	:douta	=	16'h	d5b3;
49112	:douta	=	16'h	cd73;
49113	:douta	=	16'h	c533;
49114	:douta	=	16'h	b4f3;
49115	:douta	=	16'h	b4f3;
49116	:douta	=	16'h	acf3;
49117	:douta	=	16'h	acd3;
49118	:douta	=	16'h	acd3;
49119	:douta	=	16'h	a4b3;
49120	:douta	=	16'h	a4d3;
49121	:douta	=	16'h	acf4;
49122	:douta	=	16'h	9cd3;
49123	:douta	=	16'h	8c93;
49124	:douta	=	16'h	7c32;
49125	:douta	=	16'h	7412;
49126	:douta	=	16'h	5b0e;
49127	:douta	=	16'h	422a;
49128	:douta	=	16'h	2987;
49129	:douta	=	16'h	1927;
49130	:douta	=	16'h	52ac;
49131	:douta	=	16'h	1927;
49132	:douta	=	16'h	2127;
49133	:douta	=	16'h	08a3;
49134	:douta	=	16'h	2105;
49135	:douta	=	16'h	18c5;
49136	:douta	=	16'h	2168;
49137	:douta	=	16'h	08c6;
49138	:douta	=	16'h	51c5;
49139	:douta	=	16'h	59e6;
49140	:douta	=	16'h	51c6;
49141	:douta	=	16'h	51c5;
49142	:douta	=	16'h	51c5;
49143	:douta	=	16'h	59e6;
49144	:douta	=	16'h	51c6;
49145	:douta	=	16'h	51c6;
49146	:douta	=	16'h	59e6;
49147	:douta	=	16'h	59e6;
49148	:douta	=	16'h	59c6;
49149	:douta	=	16'h	59e6;
49150	:douta	=	16'h	59e6;
49151	:douta	=	16'h	59e6;
49152	:douta	=	16'h	cd54;
49153	:douta	=	16'h	de77;
49154	:douta	=	16'h	c575;
49155	:douta	=	16'h	b534;
49156	:douta	=	16'h	acf4;
49157	:douta	=	16'h	b535;
49158	:douta	=	16'h	cdb5;
49159	:douta	=	16'h	bd75;
49160	:douta	=	16'h	b555;
49161	:douta	=	16'h	9cf5;
49162	:douta	=	16'h	8c73;
49163	:douta	=	16'h	9474;
49164	:douta	=	16'h	94b4;
49165	:douta	=	16'h	9494;
49166	:douta	=	16'h	94d5;
49167	:douta	=	16'h	8c94;
49168	:douta	=	16'h	8454;
49169	:douta	=	16'h	8433;
49170	:douta	=	16'h	8474;
49171	:douta	=	16'h	9517;
49172	:douta	=	16'h	31c6;
49173	:douta	=	16'h	20c3;
49174	:douta	=	16'h	20c2;
49175	:douta	=	16'h	20a3;
49176	:douta	=	16'h	20c3;
49177	:douta	=	16'h	20c3;
49178	:douta	=	16'h	20a3;
49179	:douta	=	16'h	20a3;
49180	:douta	=	16'h	20c3;
49181	:douta	=	16'h	20a2;
49182	:douta	=	16'h	20a2;
49183	:douta	=	16'h	20a2;
49184	:douta	=	16'h	20a2;
49185	:douta	=	16'h	20a2;
49186	:douta	=	16'h	20c2;
49187	:douta	=	16'h	20a2;
49188	:douta	=	16'h	20a2;
49189	:douta	=	16'h	20a2;
49190	:douta	=	16'h	20a2;
49191	:douta	=	16'h	20a2;
49192	:douta	=	16'h	28c2;
49193	:douta	=	16'h	28c2;
49194	:douta	=	16'h	28c2;
49195	:douta	=	16'h	28e2;
49196	:douta	=	16'h	30e3;
49197	:douta	=	16'h	3103;
49198	:douta	=	16'h	3103;
49199	:douta	=	16'h	3903;
49200	:douta	=	16'h	41c8;
49201	:douta	=	16'h	2947;
49202	:douta	=	16'h	10a4;
49203	:douta	=	16'h	4963;
49204	:douta	=	16'h	4964;
49205	:douta	=	16'h	5163;
49206	:douta	=	16'h	5184;
49207	:douta	=	16'h	5184;
49208	:douta	=	16'h	59a4;
49209	:douta	=	16'h	59a4;
49210	:douta	=	16'h	59c4;
49211	:douta	=	16'h	61c3;
49212	:douta	=	16'h	61c4;
49213	:douta	=	16'h	a573;
49214	:douta	=	16'h	8b8a;
49215	:douta	=	16'h	7244;
49216	:douta	=	16'h	6a04;
49217	:douta	=	16'h	7224;
49218	:douta	=	16'h	7244;
49219	:douta	=	16'h	7224;
49220	:douta	=	16'h	6a04;
49221	:douta	=	16'h	7a64;
49222	:douta	=	16'h	7a64;
49223	:douta	=	16'h	7aa4;
49224	:douta	=	16'h	7a84;
49225	:douta	=	16'h	7a84;
49226	:douta	=	16'h	82a5;
49227	:douta	=	16'h	8285;
49228	:douta	=	16'h	82a4;
49229	:douta	=	16'h	82a4;
49230	:douta	=	16'h	82a4;
49231	:douta	=	16'h	8ac5;
49232	:douta	=	16'h	8ac4;
49233	:douta	=	16'h	92e4;
49234	:douta	=	16'h	9305;
49235	:douta	=	16'h	9325;
49236	:douta	=	16'h	a346;
49237	:douta	=	16'h	a346;
49238	:douta	=	16'h	a345;
49239	:douta	=	16'h	a366;
49240	:douta	=	16'h	ab85;
49241	:douta	=	16'h	ab85;
49242	:douta	=	16'h	b385;
49243	:douta	=	16'h	b3a6;
49244	:douta	=	16'h	b3a5;
49245	:douta	=	16'h	bbc6;
49246	:douta	=	16'h	bbc6;
49247	:douta	=	16'h	bbc6;
49248	:douta	=	16'h	bbe6;
49249	:douta	=	16'h	bbe6;
49250	:douta	=	16'h	bbe5;
49251	:douta	=	16'h	bbe5;
49252	:douta	=	16'h	bbe5;
49253	:douta	=	16'h	c406;
49254	:douta	=	16'h	bc06;
49255	:douta	=	16'h	c426;
49256	:douta	=	16'h	c405;
49257	:douta	=	16'h	c426;
49258	:douta	=	16'h	c426;
49259	:douta	=	16'h	c426;
49260	:douta	=	16'h	c426;
49261	:douta	=	16'h	c426;
49262	:douta	=	16'h	c426;
49263	:douta	=	16'h	cc46;
49264	:douta	=	16'h	cc47;
49265	:douta	=	16'h	c426;
49266	:douta	=	16'h	cc26;
49267	:douta	=	16'h	c446;
49268	:douta	=	16'h	cc47;
49269	:douta	=	16'h	cc47;
49270	:douta	=	16'h	cc46;
49271	:douta	=	16'h	cc46;
49272	:douta	=	16'h	cc47;
49273	:douta	=	16'h	cc47;
49274	:douta	=	16'h	cc67;
49275	:douta	=	16'h	cc47;
49276	:douta	=	16'h	cc67;
49277	:douta	=	16'h	cc47;
49278	:douta	=	16'h	cc67;
49279	:douta	=	16'h	cc67;
49280	:douta	=	16'h	d467;
49281	:douta	=	16'h	cc67;
49282	:douta	=	16'h	cc67;
49283	:douta	=	16'h	d467;
49284	:douta	=	16'h	d467;
49285	:douta	=	16'h	d467;
49286	:douta	=	16'h	cc67;
49287	:douta	=	16'h	cc67;
49288	:douta	=	16'h	cc67;
49289	:douta	=	16'h	d468;
49290	:douta	=	16'h	d467;
49291	:douta	=	16'h	d467;
49292	:douta	=	16'h	d467;
49293	:douta	=	16'h	d468;
49294	:douta	=	16'h	d467;
49295	:douta	=	16'h	d467;
49296	:douta	=	16'h	d487;
49297	:douta	=	16'h	d467;
49298	:douta	=	16'h	d487;
49299	:douta	=	16'h	d467;
49300	:douta	=	16'h	d467;
49301	:douta	=	16'h	d487;
49302	:douta	=	16'h	d467;
49303	:douta	=	16'h	d467;
49304	:douta	=	16'h	d487;
49305	:douta	=	16'h	d488;
49306	:douta	=	16'h	d488;
49307	:douta	=	16'h	d488;
49308	:douta	=	16'h	d488;
49309	:douta	=	16'h	d487;
49310	:douta	=	16'h	d487;
49311	:douta	=	16'h	d487;
49312	:douta	=	16'h	d487;
49313	:douta	=	16'h	d488;
49314	:douta	=	16'h	d468;
49315	:douta	=	16'h	b50e;
49316	:douta	=	16'h	ceb7;
49317	:douta	=	16'h	cc05;
49318	:douta	=	16'h	cc68;
49319	:douta	=	16'h	cc88;
49320	:douta	=	16'h	d487;
49321	:douta	=	16'h	cc68;
49322	:douta	=	16'h	cc68;
49323	:douta	=	16'h	dca5;
49324	:douta	=	16'h	83d1;
49325	:douta	=	16'h	8c10;
49326	:douta	=	16'h	8bf1;
49327	:douta	=	16'h	736f;
49328	:douta	=	16'h	7b90;
49329	:douta	=	16'h	7b90;
49330	:douta	=	16'h	734e;
49331	:douta	=	16'h	734e;
49332	:douta	=	16'h	5a8a;
49333	:douta	=	16'h	5269;
49334	:douta	=	16'h	3965;
49335	:douta	=	16'h	49c5;
49336	:douta	=	16'h	5206;
49337	:douta	=	16'h	62e9;
49338	:douta	=	16'h	6aea;
49339	:douta	=	16'h	62e9;
49340	:douta	=	16'h	7b6c;
49341	:douta	=	16'h	9c6f;
49342	:douta	=	16'h	7b4c;
49343	:douta	=	16'h	732b;
49344	:douta	=	16'h	940e;
49345	:douta	=	16'h	940e;
49346	:douta	=	16'h	940e;
49347	:douta	=	16'h	9c2e;
49348	:douta	=	16'h	a46f;
49349	:douta	=	16'h	b4d1;
49350	:douta	=	16'h	5a69;
49351	:douta	=	16'h	838c;
49352	:douta	=	16'h	a490;
49353	:douta	=	16'h	bd31;
49354	:douta	=	16'h	bd11;
49355	:douta	=	16'h	c551;
49356	:douta	=	16'h	c572;
49357	:douta	=	16'h	cdd4;
49358	:douta	=	16'h	d5d4;
49359	:douta	=	16'h	d5f4;
49360	:douta	=	16'h	de15;
49361	:douta	=	16'h	de15;
49362	:douta	=	16'h	cd93;
49363	:douta	=	16'h	d5b3;
49364	:douta	=	16'h	d5b4;
49365	:douta	=	16'h	c572;
49366	:douta	=	16'h	c553;
49367	:douta	=	16'h	b513;
49368	:douta	=	16'h	b4f3;
49369	:douta	=	16'h	acd3;
49370	:douta	=	16'h	acd3;
49371	:douta	=	16'h	a4d4;
49372	:douta	=	16'h	a4d4;
49373	:douta	=	16'h	a4b4;
49374	:douta	=	16'h	94b5;
49375	:douta	=	16'h	9cb4;
49376	:douta	=	16'h	94b4;
49377	:douta	=	16'h	94b4;
49378	:douta	=	16'h	94d4;
49379	:douta	=	16'h	94b4;
49380	:douta	=	16'h	8453;
49381	:douta	=	16'h	8474;
49382	:douta	=	16'h	7cb6;
49383	:douta	=	16'h	7434;
49384	:douta	=	16'h	4a8d;
49385	:douta	=	16'h	29a9;
49386	:douta	=	16'h	39e8;
49387	:douta	=	16'h	2988;
49388	:douta	=	16'h	2968;
49389	:douta	=	16'h	2127;
49390	:douta	=	16'h	18c4;
49391	:douta	=	16'h	10a4;
49392	:douta	=	16'h	1946;
49393	:douta	=	16'h	2147;
49394	:douta	=	16'h	59e6;
49395	:douta	=	16'h	51e6;
49396	:douta	=	16'h	59e6;
49397	:douta	=	16'h	51c6;
49398	:douta	=	16'h	59e6;
49399	:douta	=	16'h	59e6;
49400	:douta	=	16'h	51c6;
49401	:douta	=	16'h	5a06;
49402	:douta	=	16'h	59e6;
49403	:douta	=	16'h	59e6;
49404	:douta	=	16'h	6206;
49405	:douta	=	16'h	59e6;
49406	:douta	=	16'h	6206;
49407	:douta	=	16'h	6206;
49408	:douta	=	16'h	d5b5;
49409	:douta	=	16'h	cdb5;
49410	:douta	=	16'h	bd34;
49411	:douta	=	16'h	b534;
49412	:douta	=	16'h	ad14;
49413	:douta	=	16'h	cdd5;
49414	:douta	=	16'h	bd95;
49415	:douta	=	16'h	bd55;
49416	:douta	=	16'h	ad35;
49417	:douta	=	16'h	9453;
49418	:douta	=	16'h	9473;
49419	:douta	=	16'h	9cb4;
49420	:douta	=	16'h	94b4;
49421	:douta	=	16'h	94d5;
49422	:douta	=	16'h	94b5;
49423	:douta	=	16'h	8c74;
49424	:douta	=	16'h	7c33;
49425	:douta	=	16'h	8454;
49426	:douta	=	16'h	94d6;
49427	:douta	=	16'h	2945;
49428	:douta	=	16'h	1040;
49429	:douta	=	16'h	20c3;
49430	:douta	=	16'h	20c3;
49431	:douta	=	16'h	20a3;
49432	:douta	=	16'h	20e3;
49433	:douta	=	16'h	20c3;
49434	:douta	=	16'h	20c3;
49435	:douta	=	16'h	20a2;
49436	:douta	=	16'h	20a3;
49437	:douta	=	16'h	18a1;
49438	:douta	=	16'h	18a2;
49439	:douta	=	16'h	1881;
49440	:douta	=	16'h	1881;
49441	:douta	=	16'h	20a2;
49442	:douta	=	16'h	2082;
49443	:douta	=	16'h	20a2;
49444	:douta	=	16'h	20a2;
49445	:douta	=	16'h	20a2;
49446	:douta	=	16'h	20c2;
49447	:douta	=	16'h	20c2;
49448	:douta	=	16'h	28c2;
49449	:douta	=	16'h	28e2;
49450	:douta	=	16'h	28e2;
49451	:douta	=	16'h	30e3;
49452	:douta	=	16'h	30e3;
49453	:douta	=	16'h	30e3;
49454	:douta	=	16'h	3103;
49455	:douta	=	16'h	3903;
49456	:douta	=	16'h	39e8;
49457	:douta	=	16'h	1906;
49458	:douta	=	16'h	18a4;
49459	:douta	=	16'h	4963;
49460	:douta	=	16'h	4963;
49461	:douta	=	16'h	4983;
49462	:douta	=	16'h	5184;
49463	:douta	=	16'h	51a4;
49464	:douta	=	16'h	59a4;
49465	:douta	=	16'h	59a4;
49466	:douta	=	16'h	61c4;
49467	:douta	=	16'h	59c3;
49468	:douta	=	16'h	6225;
49469	:douta	=	16'h	a4f2;
49470	:douta	=	16'h	7266;
49471	:douta	=	16'h	6a24;
49472	:douta	=	16'h	7225;
49473	:douta	=	16'h	7244;
49474	:douta	=	16'h	7244;
49475	:douta	=	16'h	8285;
49476	:douta	=	16'h	51a4;
49477	:douta	=	16'h	7a64;
49478	:douta	=	16'h	7a64;
49479	:douta	=	16'h	8284;
49480	:douta	=	16'h	8284;
49481	:douta	=	16'h	7a64;
49482	:douta	=	16'h	8285;
49483	:douta	=	16'h	7a64;
49484	:douta	=	16'h	8284;
49485	:douta	=	16'h	82a4;
49486	:douta	=	16'h	8ac5;
49487	:douta	=	16'h	8aa4;
49488	:douta	=	16'h	8ac5;
49489	:douta	=	16'h	92c4;
49490	:douta	=	16'h	9304;
49491	:douta	=	16'h	9b26;
49492	:douta	=	16'h	a346;
49493	:douta	=	16'h	a346;
49494	:douta	=	16'h	a366;
49495	:douta	=	16'h	a365;
49496	:douta	=	16'h	ab85;
49497	:douta	=	16'h	ab85;
49498	:douta	=	16'h	b3a5;
49499	:douta	=	16'h	b3a5;
49500	:douta	=	16'h	b3a6;
49501	:douta	=	16'h	b3a6;
49502	:douta	=	16'h	bbc6;
49503	:douta	=	16'h	bbc6;
49504	:douta	=	16'h	bbe6;
49505	:douta	=	16'h	bbe6;
49506	:douta	=	16'h	bc05;
49507	:douta	=	16'h	bbe5;
49508	:douta	=	16'h	c406;
49509	:douta	=	16'h	c406;
49510	:douta	=	16'h	c406;
49511	:douta	=	16'h	c406;
49512	:douta	=	16'h	c406;
49513	:douta	=	16'h	c405;
49514	:douta	=	16'h	c426;
49515	:douta	=	16'h	c426;
49516	:douta	=	16'h	c426;
49517	:douta	=	16'h	c426;
49518	:douta	=	16'h	c446;
49519	:douta	=	16'h	c446;
49520	:douta	=	16'h	c446;
49521	:douta	=	16'h	c446;
49522	:douta	=	16'h	c446;
49523	:douta	=	16'h	c446;
49524	:douta	=	16'h	cc47;
49525	:douta	=	16'h	cc47;
49526	:douta	=	16'h	cc47;
49527	:douta	=	16'h	cc47;
49528	:douta	=	16'h	cc47;
49529	:douta	=	16'h	cc47;
49530	:douta	=	16'h	cc67;
49531	:douta	=	16'h	cc47;
49532	:douta	=	16'h	cc67;
49533	:douta	=	16'h	cc67;
49534	:douta	=	16'h	cc67;
49535	:douta	=	16'h	cc67;
49536	:douta	=	16'h	cc46;
49537	:douta	=	16'h	cc46;
49538	:douta	=	16'h	cc67;
49539	:douta	=	16'h	cc67;
49540	:douta	=	16'h	d467;
49541	:douta	=	16'h	cc67;
49542	:douta	=	16'h	cc47;
49543	:douta	=	16'h	d468;
49544	:douta	=	16'h	d468;
49545	:douta	=	16'h	d468;
49546	:douta	=	16'h	d488;
49547	:douta	=	16'h	d468;
49548	:douta	=	16'h	d467;
49549	:douta	=	16'h	d467;
49550	:douta	=	16'h	cc67;
49551	:douta	=	16'h	d487;
49552	:douta	=	16'h	d467;
49553	:douta	=	16'h	d467;
49554	:douta	=	16'h	d467;
49555	:douta	=	16'h	d487;
49556	:douta	=	16'h	d487;
49557	:douta	=	16'h	d487;
49558	:douta	=	16'h	cc67;
49559	:douta	=	16'h	d488;
49560	:douta	=	16'h	cc68;
49561	:douta	=	16'h	d488;
49562	:douta	=	16'h	d488;
49563	:douta	=	16'h	d488;
49564	:douta	=	16'h	d488;
49565	:douta	=	16'h	d488;
49566	:douta	=	16'h	d488;
49567	:douta	=	16'h	d488;
49568	:douta	=	16'h	d488;
49569	:douta	=	16'h	d488;
49570	:douta	=	16'h	d487;
49571	:douta	=	16'h	acce;
49572	:douta	=	16'h	d677;
49573	:douta	=	16'h	cc03;
49574	:douta	=	16'h	cc66;
49575	:douta	=	16'h	cc46;
49576	:douta	=	16'h	cc24;
49577	:douta	=	16'h	cc04;
49578	:douta	=	16'h	cc25;
49579	:douta	=	16'h	c426;
49580	:douta	=	16'h	bc4a;
49581	:douta	=	16'h	8c30;
49582	:douta	=	16'h	8c31;
49583	:douta	=	16'h	7b8f;
49584	:douta	=	16'h	734d;
49585	:douta	=	16'h	5a48;
49586	:douta	=	16'h	41c5;
49587	:douta	=	16'h	4a06;
49588	:douta	=	16'h	62a9;
49589	:douta	=	16'h	732a;
49590	:douta	=	16'h	6b0a;
49591	:douta	=	16'h	6b0b;
49592	:douta	=	16'h	8bee;
49593	:douta	=	16'h	734b;
49594	:douta	=	16'h	7b8c;
49595	:douta	=	16'h	8bed;
49596	:douta	=	16'h	bd51;
49597	:douta	=	16'h	b511;
49598	:douta	=	16'h	7b8c;
49599	:douta	=	16'h	a48f;
49600	:douta	=	16'h	acd0;
49601	:douta	=	16'h	b510;
49602	:douta	=	16'h	b4d0;
49603	:douta	=	16'h	bd10;
49604	:douta	=	16'h	c531;
49605	:douta	=	16'h	d5d3;
49606	:douta	=	16'h	8bce;
49607	:douta	=	16'h	62aa;
49608	:douta	=	16'h	acd1;
49609	:douta	=	16'h	bd32;
49610	:douta	=	16'h	c573;
49611	:douta	=	16'h	cd93;
49612	:douta	=	16'h	d5b3;
49613	:douta	=	16'h	d5f4;
49614	:douta	=	16'h	d614;
49615	:douta	=	16'h	de15;
49616	:douta	=	16'h	d5b3;
49617	:douta	=	16'h	d5b3;
49618	:douta	=	16'h	acf3;
49619	:douta	=	16'h	acf3;
49620	:douta	=	16'h	acf4;
49621	:douta	=	16'h	9c94;
49622	:douta	=	16'h	9cb5;
49623	:douta	=	16'h	9cb4;
49624	:douta	=	16'h	9cb4;
49625	:douta	=	16'h	9cb4;
49626	:douta	=	16'h	8c74;
49627	:douta	=	16'h	8c53;
49628	:douta	=	16'h	8c73;
49629	:douta	=	16'h	8433;
49630	:douta	=	16'h	7c12;
49631	:douta	=	16'h	7390;
49632	:douta	=	16'h	738f;
49633	:douta	=	16'h	6b2d;
49634	:douta	=	16'h	5269;
49635	:douta	=	16'h	41c7;
49636	:douta	=	16'h	3985;
49637	:douta	=	16'h	3144;
49638	:douta	=	16'h	28e2;
49639	:douta	=	16'h	2903;
49640	:douta	=	16'h	422a;
49641	:douta	=	16'h	31ea;
49642	:douta	=	16'h	2168;
49643	:douta	=	16'h	52ac;
49644	:douta	=	16'h	2168;
49645	:douta	=	16'h	2126;
49646	:douta	=	16'h	2126;
49647	:douta	=	16'h	2127;
49648	:douta	=	16'h	0042;
49649	:douta	=	16'h	5a8a;
49650	:douta	=	16'h	59e6;
49651	:douta	=	16'h	59e6;
49652	:douta	=	16'h	59e6;
49653	:douta	=	16'h	59c6;
49654	:douta	=	16'h	59e6;
49655	:douta	=	16'h	59e6;
49656	:douta	=	16'h	6206;
49657	:douta	=	16'h	6206;
49658	:douta	=	16'h	5a06;
49659	:douta	=	16'h	6206;
49660	:douta	=	16'h	6206;
49661	:douta	=	16'h	6206;
49662	:douta	=	16'h	6226;
49663	:douta	=	16'h	6206;
49664	:douta	=	16'h	de16;
49665	:douta	=	16'h	bd75;
49666	:douta	=	16'h	b514;
49667	:douta	=	16'h	b555;
49668	:douta	=	16'h	b555;
49669	:douta	=	16'h	d5f6;
49670	:douta	=	16'h	bd75;
49671	:douta	=	16'h	bd55;
49672	:douta	=	16'h	ad35;
49673	:douta	=	16'h	8c32;
49674	:douta	=	16'h	9473;
49675	:douta	=	16'h	9cb4;
49676	:douta	=	16'h	94b5;
49677	:douta	=	16'h	94d5;
49678	:douta	=	16'h	94b5;
49679	:douta	=	16'h	8c74;
49680	:douta	=	16'h	8433;
49681	:douta	=	16'h	8454;
49682	:douta	=	16'h	9d58;
49683	:douta	=	16'h	0800;
49684	:douta	=	16'h	20c3;
49685	:douta	=	16'h	20a3;
49686	:douta	=	16'h	20c3;
49687	:douta	=	16'h	20a3;
49688	:douta	=	16'h	20c3;
49689	:douta	=	16'h	20e3;
49690	:douta	=	16'h	20c3;
49691	:douta	=	16'h	20c3;
49692	:douta	=	16'h	20a2;
49693	:douta	=	16'h	18a1;
49694	:douta	=	16'h	1881;
49695	:douta	=	16'h	1881;
49696	:douta	=	16'h	2082;
49697	:douta	=	16'h	20a2;
49698	:douta	=	16'h	20a2;
49699	:douta	=	16'h	20a2;
49700	:douta	=	16'h	20a2;
49701	:douta	=	16'h	20a2;
49702	:douta	=	16'h	20a2;
49703	:douta	=	16'h	20c2;
49704	:douta	=	16'h	20c2;
49705	:douta	=	16'h	28c2;
49706	:douta	=	16'h	28e2;
49707	:douta	=	16'h	30e3;
49708	:douta	=	16'h	3103;
49709	:douta	=	16'h	30e2;
49710	:douta	=	16'h	3923;
49711	:douta	=	16'h	3902;
49712	:douta	=	16'h	3a09;
49713	:douta	=	16'h	18e5;
49714	:douta	=	16'h	20a4;
49715	:douta	=	16'h	4984;
49716	:douta	=	16'h	4964;
49717	:douta	=	16'h	4983;
49718	:douta	=	16'h	51a4;
49719	:douta	=	16'h	51a4;
49720	:douta	=	16'h	59a4;
49721	:douta	=	16'h	59c4;
49722	:douta	=	16'h	61c4;
49723	:douta	=	16'h	61c3;
49724	:douta	=	16'h	6267;
49725	:douta	=	16'h	9c8f;
49726	:douta	=	16'h	6a04;
49727	:douta	=	16'h	7224;
49728	:douta	=	16'h	7224;
49729	:douta	=	16'h	7245;
49730	:douta	=	16'h	7244;
49731	:douta	=	16'h	8285;
49732	:douta	=	16'h	4984;
49733	:douta	=	16'h	7a64;
49734	:douta	=	16'h	8284;
49735	:douta	=	16'h	7a64;
49736	:douta	=	16'h	8284;
49737	:douta	=	16'h	8285;
49738	:douta	=	16'h	8285;
49739	:douta	=	16'h	8284;
49740	:douta	=	16'h	82a4;
49741	:douta	=	16'h	82a5;
49742	:douta	=	16'h	8ac5;
49743	:douta	=	16'h	8ac5;
49744	:douta	=	16'h	8ac4;
49745	:douta	=	16'h	92e5;
49746	:douta	=	16'h	9305;
49747	:douta	=	16'h	9b26;
49748	:douta	=	16'h	a346;
49749	:douta	=	16'h	a346;
49750	:douta	=	16'h	a345;
49751	:douta	=	16'h	ab85;
49752	:douta	=	16'h	ab65;
49753	:douta	=	16'h	b385;
49754	:douta	=	16'h	b3a5;
49755	:douta	=	16'h	b3a6;
49756	:douta	=	16'h	b3a5;
49757	:douta	=	16'h	bbc6;
49758	:douta	=	16'h	bbc6;
49759	:douta	=	16'h	bbe6;
49760	:douta	=	16'h	bbe6;
49761	:douta	=	16'h	bbe6;
49762	:douta	=	16'h	bc06;
49763	:douta	=	16'h	bc06;
49764	:douta	=	16'h	c406;
49765	:douta	=	16'h	c406;
49766	:douta	=	16'h	c406;
49767	:douta	=	16'h	c406;
49768	:douta	=	16'h	c426;
49769	:douta	=	16'h	c426;
49770	:douta	=	16'h	c426;
49771	:douta	=	16'h	c426;
49772	:douta	=	16'h	c426;
49773	:douta	=	16'h	c426;
49774	:douta	=	16'h	c426;
49775	:douta	=	16'h	c426;
49776	:douta	=	16'h	c446;
49777	:douta	=	16'h	c446;
49778	:douta	=	16'h	c446;
49779	:douta	=	16'h	cc47;
49780	:douta	=	16'h	cc47;
49781	:douta	=	16'h	cc47;
49782	:douta	=	16'h	cc67;
49783	:douta	=	16'h	cc47;
49784	:douta	=	16'h	cc47;
49785	:douta	=	16'h	cc47;
49786	:douta	=	16'h	cc47;
49787	:douta	=	16'h	cc47;
49788	:douta	=	16'h	cc67;
49789	:douta	=	16'h	cc47;
49790	:douta	=	16'h	cc67;
49791	:douta	=	16'h	cc67;
49792	:douta	=	16'h	cc47;
49793	:douta	=	16'h	cc47;
49794	:douta	=	16'h	cc67;
49795	:douta	=	16'h	cc67;
49796	:douta	=	16'h	cc67;
49797	:douta	=	16'h	cc47;
49798	:douta	=	16'h	cc67;
49799	:douta	=	16'h	d467;
49800	:douta	=	16'h	d467;
49801	:douta	=	16'h	d468;
49802	:douta	=	16'h	d467;
49803	:douta	=	16'h	cc67;
49804	:douta	=	16'h	d488;
49805	:douta	=	16'h	d467;
49806	:douta	=	16'h	d487;
49807	:douta	=	16'h	d487;
49808	:douta	=	16'h	d487;
49809	:douta	=	16'h	d467;
49810	:douta	=	16'h	d487;
49811	:douta	=	16'h	d487;
49812	:douta	=	16'h	d487;
49813	:douta	=	16'h	d467;
49814	:douta	=	16'h	cc67;
49815	:douta	=	16'h	d488;
49816	:douta	=	16'h	d488;
49817	:douta	=	16'h	d488;
49818	:douta	=	16'h	d487;
49819	:douta	=	16'h	cc87;
49820	:douta	=	16'h	d488;
49821	:douta	=	16'h	d487;
49822	:douta	=	16'h	d467;
49823	:douta	=	16'h	d466;
49824	:douta	=	16'h	cc66;
49825	:douta	=	16'h	d444;
49826	:douta	=	16'h	d423;
49827	:douta	=	16'h	a48c;
49828	:douta	=	16'h	ce76;
49829	:douta	=	16'h	c3e0;
49830	:douta	=	16'h	cc69;
49831	:douta	=	16'h	ccaa;
49832	:douta	=	16'h	d52d;
49833	:douta	=	16'h	d54e;
49834	:douta	=	16'h	d5f2;
49835	:douta	=	16'h	e634;
49836	:douta	=	16'h	f6f8;
49837	:douta	=	16'h	8bef;
49838	:douta	=	16'h	83af;
49839	:douta	=	16'h	5a69;
49840	:douta	=	16'h	49e7;
49841	:douta	=	16'h	41c5;
49842	:douta	=	16'h	62ca;
49843	:douta	=	16'h	6b0b;
49844	:douta	=	16'h	6aea;
49845	:douta	=	16'h	6b0a;
49846	:douta	=	16'h	6b0b;
49847	:douta	=	16'h	942f;
49848	:douta	=	16'h	9c4e;
49849	:douta	=	16'h	83ad;
49850	:douta	=	16'h	942f;
49851	:douta	=	16'h	942e;
49852	:douta	=	16'h	b510;
49853	:douta	=	16'h	acb0;
49854	:douta	=	16'h	a48f;
49855	:douta	=	16'h	cdd3;
49856	:douta	=	16'h	b511;
49857	:douta	=	16'h	bd31;
49858	:douta	=	16'h	bd31;
49859	:douta	=	16'h	c552;
49860	:douta	=	16'h	cdb3;
49861	:douta	=	16'h	d5d4;
49862	:douta	=	16'h	bd52;
49863	:douta	=	16'h	62ca;
49864	:douta	=	16'h	acd1;
49865	:douta	=	16'h	c572;
49866	:douta	=	16'h	cdb3;
49867	:douta	=	16'h	d5b3;
49868	:douta	=	16'h	cdb3;
49869	:douta	=	16'h	d5d4;
49870	:douta	=	16'h	d5b3;
49871	:douta	=	16'h	cd53;
49872	:douta	=	16'h	b4f2;
49873	:douta	=	16'h	b4d3;
49874	:douta	=	16'h	9cb3;
49875	:douta	=	16'h	a4d4;
49876	:douta	=	16'h	9cb4;
49877	:douta	=	16'h	94b4;
49878	:douta	=	16'h	94b4;
49879	:douta	=	16'h	8c93;
49880	:douta	=	16'h	8c73;
49881	:douta	=	16'h	8c73;
49882	:douta	=	16'h	8433;
49883	:douta	=	16'h	7bf1;
49884	:douta	=	16'h	7bf2;
49885	:douta	=	16'h	73b1;
49886	:douta	=	16'h	736e;
49887	:douta	=	16'h	5289;
49888	:douta	=	16'h	49e7;
49889	:douta	=	16'h	2903;
49890	:douta	=	16'h	2081;
49891	:douta	=	16'h	20c2;
49892	:douta	=	16'h	4a06;
49893	:douta	=	16'h	4a06;
49894	:douta	=	16'h	5228;
49895	:douta	=	16'h	526a;
49896	:douta	=	16'h	5aee;
49897	:douta	=	16'h	426d;
49898	:douta	=	16'h	29eb;
49899	:douta	=	16'h	62ee;
49900	:douta	=	16'h	0863;
49901	:douta	=	16'h	1883;
49902	:douta	=	16'h	10a3;
49903	:douta	=	16'h	18e4;
49904	:douta	=	16'h	0001;
49905	:douta	=	16'h	3187;
49906	:douta	=	16'h	59c5;
49907	:douta	=	16'h	59e6;
49908	:douta	=	16'h	59e7;
49909	:douta	=	16'h	6206;
49910	:douta	=	16'h	59e6;
49911	:douta	=	16'h	6206;
49912	:douta	=	16'h	6206;
49913	:douta	=	16'h	6206;
49914	:douta	=	16'h	6206;
49915	:douta	=	16'h	6226;
49916	:douta	=	16'h	6206;
49917	:douta	=	16'h	6206;
49918	:douta	=	16'h	6206;
49919	:douta	=	16'h	6a26;
49920	:douta	=	16'h	e678;
49921	:douta	=	16'h	b534;
49922	:douta	=	16'h	bd34;
49923	:douta	=	16'h	ad15;
49924	:douta	=	16'h	cdb5;
49925	:douta	=	16'h	cdd6;
49926	:douta	=	16'h	bd75;
49927	:douta	=	16'h	bd55;
49928	:douta	=	16'h	a4f5;
49929	:douta	=	16'h	9493;
49930	:douta	=	16'h	9473;
49931	:douta	=	16'h	a4f5;
49932	:douta	=	16'h	94d5;
49933	:douta	=	16'h	94b5;
49934	:douta	=	16'h	8c75;
49935	:douta	=	16'h	8453;
49936	:douta	=	16'h	8454;
49937	:douta	=	16'h	8c75;
49938	:douta	=	16'h	52cc;
49939	:douta	=	16'h	20c3;
49940	:douta	=	16'h	20c3;
49941	:douta	=	16'h	20e3;
49942	:douta	=	16'h	20e3;
49943	:douta	=	16'h	20c3;
49944	:douta	=	16'h	20c3;
49945	:douta	=	16'h	20c3;
49946	:douta	=	16'h	20a3;
49947	:douta	=	16'h	20c3;
49948	:douta	=	16'h	1881;
49949	:douta	=	16'h	1881;
49950	:douta	=	16'h	2082;
49951	:douta	=	16'h	20a2;
49952	:douta	=	16'h	1881;
49953	:douta	=	16'h	20a2;
49954	:douta	=	16'h	20a2;
49955	:douta	=	16'h	20a2;
49956	:douta	=	16'h	20a2;
49957	:douta	=	16'h	20c2;
49958	:douta	=	16'h	20c2;
49959	:douta	=	16'h	28c2;
49960	:douta	=	16'h	28e3;
49961	:douta	=	16'h	28c2;
49962	:douta	=	16'h	28e2;
49963	:douta	=	16'h	30e2;
49964	:douta	=	16'h	30e2;
49965	:douta	=	16'h	3103;
49966	:douta	=	16'h	3123;
49967	:douta	=	16'h	3903;
49968	:douta	=	16'h	3209;
49969	:douta	=	16'h	10a4;
49970	:douta	=	16'h	3104;
49971	:douta	=	16'h	4964;
49972	:douta	=	16'h	4964;
49973	:douta	=	16'h	51a4;
49974	:douta	=	16'h	59a4;
49975	:douta	=	16'h	59a4;
49976	:douta	=	16'h	59c4;
49977	:douta	=	16'h	59c4;
49978	:douta	=	16'h	61e4;
49979	:douta	=	16'h	61c3;
49980	:douta	=	16'h	6b0a;
49981	:douta	=	16'h	940c;
49982	:douta	=	16'h	69e3;
49983	:douta	=	16'h	7224;
49984	:douta	=	16'h	7244;
49985	:douta	=	16'h	7224;
49986	:douta	=	16'h	7244;
49987	:douta	=	16'h	7a44;
49988	:douta	=	16'h	4164;
49989	:douta	=	16'h	82a4;
49990	:douta	=	16'h	7a85;
49991	:douta	=	16'h	7aa5;
49992	:douta	=	16'h	7a64;
49993	:douta	=	16'h	8265;
49994	:douta	=	16'h	8285;
49995	:douta	=	16'h	8285;
49996	:douta	=	16'h	82a4;
49997	:douta	=	16'h	82a4;
49998	:douta	=	16'h	8ac5;
49999	:douta	=	16'h	8ac5;
50000	:douta	=	16'h	8ac5;
50001	:douta	=	16'h	9305;
50002	:douta	=	16'h	9305;
50003	:douta	=	16'h	9b25;
50004	:douta	=	16'h	a346;
50005	:douta	=	16'h	a346;
50006	:douta	=	16'h	a366;
50007	:douta	=	16'h	ab66;
50008	:douta	=	16'h	ab85;
50009	:douta	=	16'h	ab85;
50010	:douta	=	16'h	b3a5;
50011	:douta	=	16'h	b3c6;
50012	:douta	=	16'h	b3c6;
50013	:douta	=	16'h	b3a6;
50014	:douta	=	16'h	bbc6;
50015	:douta	=	16'h	bbe6;
50016	:douta	=	16'h	bbe6;
50017	:douta	=	16'h	bbe5;
50018	:douta	=	16'h	bbe5;
50019	:douta	=	16'h	c405;
50020	:douta	=	16'h	bbe5;
50021	:douta	=	16'h	c406;
50022	:douta	=	16'h	c406;
50023	:douta	=	16'h	c406;
50024	:douta	=	16'h	c406;
50025	:douta	=	16'h	c426;
50026	:douta	=	16'h	c426;
50027	:douta	=	16'h	c426;
50028	:douta	=	16'h	c426;
50029	:douta	=	16'h	c446;
50030	:douta	=	16'h	c426;
50031	:douta	=	16'h	cc26;
50032	:douta	=	16'h	c426;
50033	:douta	=	16'h	cc27;
50034	:douta	=	16'h	cc27;
50035	:douta	=	16'h	cc47;
50036	:douta	=	16'h	cc67;
50037	:douta	=	16'h	cc47;
50038	:douta	=	16'h	cc67;
50039	:douta	=	16'h	cc47;
50040	:douta	=	16'h	cc67;
50041	:douta	=	16'h	cc47;
50042	:douta	=	16'h	cc48;
50043	:douta	=	16'h	cc68;
50044	:douta	=	16'h	cc67;
50045	:douta	=	16'h	cc66;
50046	:douta	=	16'h	cc67;
50047	:douta	=	16'h	cc67;
50048	:douta	=	16'h	d467;
50049	:douta	=	16'h	cc67;
50050	:douta	=	16'h	cc87;
50051	:douta	=	16'h	cc87;
50052	:douta	=	16'h	d488;
50053	:douta	=	16'h	d467;
50054	:douta	=	16'h	d467;
50055	:douta	=	16'h	d468;
50056	:douta	=	16'h	d468;
50057	:douta	=	16'h	d467;
50058	:douta	=	16'h	cc67;
50059	:douta	=	16'h	cc67;
50060	:douta	=	16'h	cc68;
50061	:douta	=	16'h	d488;
50062	:douta	=	16'h	d468;
50063	:douta	=	16'h	d487;
50064	:douta	=	16'h	d467;
50065	:douta	=	16'h	d467;
50066	:douta	=	16'h	d466;
50067	:douta	=	16'h	cc45;
50068	:douta	=	16'h	cc25;
50069	:douta	=	16'h	cc25;
50070	:douta	=	16'h	cc23;
50071	:douta	=	16'h	cc25;
50072	:douta	=	16'h	cc47;
50073	:douta	=	16'h	cc89;
50074	:douta	=	16'h	cccb;
50075	:douta	=	16'h	d52e;
50076	:douta	=	16'h	d5b1;
50077	:douta	=	16'h	ddf2;
50078	:douta	=	16'h	e675;
50079	:douta	=	16'h	e6b6;
50080	:douta	=	16'h	ef19;
50081	:douta	=	16'h	f77b;
50082	:douta	=	16'h	f7bc;
50083	:douta	=	16'h	f79b;
50084	:douta	=	16'h	f77a;
50085	:douta	=	16'h	fffd;
50086	:douta	=	16'h	ff9b;
50087	:douta	=	16'h	f799;
50088	:douta	=	16'h	ef17;
50089	:douta	=	16'h	eed6;
50090	:douta	=	16'h	e652;
50091	:douta	=	16'h	e612;
50092	:douta	=	16'h	d5ae;
50093	:douta	=	16'h	cd0c;
50094	:douta	=	16'h	93ce;
50095	:douta	=	16'h	7b6c;
50096	:douta	=	16'h	83cd;
50097	:douta	=	16'h	734b;
50098	:douta	=	16'h	734b;
50099	:douta	=	16'h	7b6c;
50100	:douta	=	16'h	734c;
50101	:douta	=	16'h	7b4c;
50102	:douta	=	16'h	8bee;
50103	:douta	=	16'h	944f;
50104	:douta	=	16'h	940e;
50105	:douta	=	16'h	acd0;
50106	:douta	=	16'h	b4d0;
50107	:douta	=	16'h	acaf;
50108	:douta	=	16'h	b4f0;
50109	:douta	=	16'h	9c2e;
50110	:douta	=	16'h	de55;
50111	:douta	=	16'h	de35;
50112	:douta	=	16'h	bd12;
50113	:douta	=	16'h	d5f5;
50114	:douta	=	16'h	d614;
50115	:douta	=	16'h	d5f4;
50116	:douta	=	16'h	cdb4;
50117	:douta	=	16'h	c5b4;
50118	:douta	=	16'h	d5f4;
50119	:douta	=	16'h	c5d4;
50120	:douta	=	16'h	acd1;
50121	:douta	=	16'h	acd1;
50122	:douta	=	16'h	d5d4;
50123	:douta	=	16'h	d5b4;
50124	:douta	=	16'h	c554;
50125	:douta	=	16'h	acb3;
50126	:douta	=	16'h	9c92;
50127	:douta	=	16'h	9453;
50128	:douta	=	16'h	8452;
50129	:douta	=	16'h	8453;
50130	:douta	=	16'h	8452;
50131	:douta	=	16'h	7bf1;
50132	:douta	=	16'h	8c53;
50133	:douta	=	16'h	7bf1;
50134	:douta	=	16'h	7bd2;
50135	:douta	=	16'h	7bd1;
50136	:douta	=	16'h	7390;
50137	:douta	=	16'h	6b0d;
50138	:douta	=	16'h	4a07;
50139	:douta	=	16'h	49e7;
50140	:douta	=	16'h	2903;
50141	:douta	=	16'h	18a2;
50142	:douta	=	16'h	1881;
50143	:douta	=	16'h	3144;
50144	:douta	=	16'h	3965;
50145	:douta	=	16'h	5208;
50146	:douta	=	16'h	62ca;
50147	:douta	=	16'h	6aea;
50148	:douta	=	16'h	7b8d;
50149	:douta	=	16'h	734e;
50150	:douta	=	16'h	52cd;
50151	:douta	=	16'h	52cd;
50152	:douta	=	16'h	52cd;
50153	:douta	=	16'h	5b31;
50154	:douta	=	16'h	5310;
50155	:douta	=	16'h	6b4f;
50156	:douta	=	16'h	4aef;
50157	:douta	=	16'h	320b;
50158	:douta	=	16'h	2968;
50159	:douta	=	16'h	2127;
50160	:douta	=	16'h	08a4;
50161	:douta	=	16'h	0022;
50162	:douta	=	16'h	7267;
50163	:douta	=	16'h	6206;
50164	:douta	=	16'h	6206;
50165	:douta	=	16'h	6207;
50166	:douta	=	16'h	6a26;
50167	:douta	=	16'h	61e6;
50168	:douta	=	16'h	61c5;
50169	:douta	=	16'h	61c5;
50170	:douta	=	16'h	59a5;
50171	:douta	=	16'h	59a5;
50172	:douta	=	16'h	61e5;
50173	:douta	=	16'h	6a47;
50174	:douta	=	16'h	6a89;
50175	:douta	=	16'h	7b4b;
50176	:douta	=	16'h	e698;
50177	:douta	=	16'h	b513;
50178	:douta	=	16'h	c575;
50179	:douta	=	16'h	a4b4;
50180	:douta	=	16'h	d5f6;
50181	:douta	=	16'h	c5b5;
50182	:douta	=	16'h	bd54;
50183	:douta	=	16'h	b555;
50184	:douta	=	16'h	9cb4;
50185	:douta	=	16'h	9c94;
50186	:douta	=	16'h	9473;
50187	:douta	=	16'h	9cd5;
50188	:douta	=	16'h	94b5;
50189	:douta	=	16'h	94b5;
50190	:douta	=	16'h	8c74;
50191	:douta	=	16'h	8c54;
50192	:douta	=	16'h	8c54;
50193	:douta	=	16'h	9d17;
50194	:douta	=	16'h	18a3;
50195	:douta	=	16'h	20c3;
50196	:douta	=	16'h	20e3;
50197	:douta	=	16'h	20e3;
50198	:douta	=	16'h	20e3;
50199	:douta	=	16'h	20c3;
50200	:douta	=	16'h	20c3;
50201	:douta	=	16'h	20e3;
50202	:douta	=	16'h	20a3;
50203	:douta	=	16'h	20c3;
50204	:douta	=	16'h	1881;
50205	:douta	=	16'h	2082;
50206	:douta	=	16'h	20a2;
50207	:douta	=	16'h	20a2;
50208	:douta	=	16'h	20a2;
50209	:douta	=	16'h	20a2;
50210	:douta	=	16'h	20a2;
50211	:douta	=	16'h	20a2;
50212	:douta	=	16'h	20a2;
50213	:douta	=	16'h	20a2;
50214	:douta	=	16'h	20a2;
50215	:douta	=	16'h	28e2;
50216	:douta	=	16'h	28e2;
50217	:douta	=	16'h	28c2;
50218	:douta	=	16'h	28e2;
50219	:douta	=	16'h	30e2;
50220	:douta	=	16'h	3103;
50221	:douta	=	16'h	3103;
50222	:douta	=	16'h	3923;
50223	:douta	=	16'h	3923;
50224	:douta	=	16'h	3a09;
50225	:douta	=	16'h	10a4;
50226	:douta	=	16'h	3923;
50227	:douta	=	16'h	4984;
50228	:douta	=	16'h	4984;
50229	:douta	=	16'h	5184;
50230	:douta	=	16'h	51a4;
50231	:douta	=	16'h	51a4;
50232	:douta	=	16'h	59c4;
50233	:douta	=	16'h	59c4;
50234	:douta	=	16'h	61e4;
50235	:douta	=	16'h	61e3;
50236	:douta	=	16'h	7b6c;
50237	:douta	=	16'h	93aa;
50238	:douta	=	16'h	69c3;
50239	:douta	=	16'h	7224;
50240	:douta	=	16'h	7244;
50241	:douta	=	16'h	7244;
50242	:douta	=	16'h	7244;
50243	:douta	=	16'h	7a65;
50244	:douta	=	16'h	4984;
50245	:douta	=	16'h	8ac5;
50246	:douta	=	16'h	7aa4;
50247	:douta	=	16'h	8284;
50248	:douta	=	16'h	7a64;
50249	:douta	=	16'h	7a85;
50250	:douta	=	16'h	8285;
50251	:douta	=	16'h	8285;
50252	:douta	=	16'h	82a4;
50253	:douta	=	16'h	8ac5;
50254	:douta	=	16'h	8ac4;
50255	:douta	=	16'h	8ac5;
50256	:douta	=	16'h	8ac4;
50257	:douta	=	16'h	92e5;
50258	:douta	=	16'h	9305;
50259	:douta	=	16'h	9b26;
50260	:douta	=	16'h	a346;
50261	:douta	=	16'h	a346;
50262	:douta	=	16'h	a366;
50263	:douta	=	16'h	ab86;
50264	:douta	=	16'h	b385;
50265	:douta	=	16'h	ab85;
50266	:douta	=	16'h	b385;
50267	:douta	=	16'h	b3c6;
50268	:douta	=	16'h	b3c6;
50269	:douta	=	16'h	bbc6;
50270	:douta	=	16'h	bbc6;
50271	:douta	=	16'h	bbe6;
50272	:douta	=	16'h	bbe6;
50273	:douta	=	16'h	bbe5;
50274	:douta	=	16'h	c406;
50275	:douta	=	16'h	bc06;
50276	:douta	=	16'h	c406;
50277	:douta	=	16'h	c406;
50278	:douta	=	16'h	c406;
50279	:douta	=	16'h	c406;
50280	:douta	=	16'h	c406;
50281	:douta	=	16'h	c426;
50282	:douta	=	16'h	c426;
50283	:douta	=	16'h	c426;
50284	:douta	=	16'h	c446;
50285	:douta	=	16'h	c426;
50286	:douta	=	16'h	c426;
50287	:douta	=	16'h	c426;
50288	:douta	=	16'h	c426;
50289	:douta	=	16'h	cc47;
50290	:douta	=	16'h	cc47;
50291	:douta	=	16'h	cc47;
50292	:douta	=	16'h	cc26;
50293	:douta	=	16'h	cc47;
50294	:douta	=	16'h	cc47;
50295	:douta	=	16'h	cc67;
50296	:douta	=	16'h	cc47;
50297	:douta	=	16'h	cc67;
50298	:douta	=	16'h	cc67;
50299	:douta	=	16'h	cc67;
50300	:douta	=	16'h	cc66;
50301	:douta	=	16'h	cc68;
50302	:douta	=	16'h	cc67;
50303	:douta	=	16'h	cc67;
50304	:douta	=	16'h	cc67;
50305	:douta	=	16'h	cc67;
50306	:douta	=	16'h	d467;
50307	:douta	=	16'h	cc68;
50308	:douta	=	16'h	d468;
50309	:douta	=	16'h	d467;
50310	:douta	=	16'h	d467;
50311	:douta	=	16'h	cc87;
50312	:douta	=	16'h	cc87;
50313	:douta	=	16'h	d467;
50314	:douta	=	16'h	d467;
50315	:douta	=	16'h	d466;
50316	:douta	=	16'h	d446;
50317	:douta	=	16'h	cc23;
50318	:douta	=	16'h	cc21;
50319	:douta	=	16'h	cc23;
50320	:douta	=	16'h	cc03;
50321	:douta	=	16'h	cc25;
50322	:douta	=	16'h	cc67;
50323	:douta	=	16'h	cc89;
50324	:douta	=	16'h	d52c;
50325	:douta	=	16'h	d56d;
50326	:douta	=	16'h	ddd1;
50327	:douta	=	16'h	e655;
50328	:douta	=	16'h	e697;
50329	:douta	=	16'h	eef8;
50330	:douta	=	16'h	ef59;
50331	:douta	=	16'h	f79c;
50332	:douta	=	16'h	ffdd;
50333	:douta	=	16'h	fffd;
50334	:douta	=	16'h	fffd;
50335	:douta	=	16'h	ffdc;
50336	:douta	=	16'h	ff9b;
50337	:douta	=	16'h	f738;
50338	:douta	=	16'h	f6f7;
50339	:douta	=	16'h	e694;
50340	:douta	=	16'h	e632;
50341	:douta	=	16'h	ddd0;
50342	:douta	=	16'h	d56d;
50343	:douta	=	16'h	d52b;
50344	:douta	=	16'h	cc88;
50345	:douta	=	16'h	cc87;
50346	:douta	=	16'h	cc46;
50347	:douta	=	16'h	cc26;
50348	:douta	=	16'h	c404;
50349	:douta	=	16'h	d444;
50350	:douta	=	16'h	c48c;
50351	:douta	=	16'h	83ad;
50352	:douta	=	16'h	8c0e;
50353	:douta	=	16'h	734b;
50354	:douta	=	16'h	83cd;
50355	:douta	=	16'h	7b8c;
50356	:douta	=	16'h	83ce;
50357	:douta	=	16'h	83cd;
50358	:douta	=	16'h	944f;
50359	:douta	=	16'h	9c4e;
50360	:douta	=	16'h	a4af;
50361	:douta	=	16'h	b4f1;
50362	:douta	=	16'h	b4f0;
50363	:douta	=	16'h	b510;
50364	:douta	=	16'h	b4f0;
50365	:douta	=	16'h	9c4f;
50366	:douta	=	16'h	d616;
50367	:douta	=	16'h	cdb4;
50368	:douta	=	16'h	acd2;
50369	:douta	=	16'h	de35;
50370	:douta	=	16'h	cdb4;
50371	:douta	=	16'h	de34;
50372	:douta	=	16'h	cdd4;
50373	:douta	=	16'h	cd94;
50374	:douta	=	16'h	acd2;
50375	:douta	=	16'h	d5f6;
50376	:douta	=	16'h	bd33;
50377	:douta	=	16'h	acd3;
50378	:douta	=	16'h	d5b3;
50379	:douta	=	16'h	b514;
50380	:douta	=	16'h	a4d4;
50381	:douta	=	16'h	8c53;
50382	:douta	=	16'h	8c53;
50383	:douta	=	16'h	8432;
50384	:douta	=	16'h	83f2;
50385	:douta	=	16'h	8412;
50386	:douta	=	16'h	7bb1;
50387	:douta	=	16'h	73d1;
50388	:douta	=	16'h	7c12;
50389	:douta	=	16'h	738f;
50390	:douta	=	16'h	738e;
50391	:douta	=	16'h	62cb;
50392	:douta	=	16'h	5248;
50393	:douta	=	16'h	3144;
50394	:douta	=	16'h	1881;
50395	:douta	=	16'h	1081;
50396	:douta	=	16'h	2924;
50397	:douta	=	16'h	3165;
50398	:douta	=	16'h	3985;
50399	:douta	=	16'h	5227;
50400	:douta	=	16'h	5248;
50401	:douta	=	16'h	6aea;
50402	:douta	=	16'h	734b;
50403	:douta	=	16'h	734b;
50404	:douta	=	16'h	4a07;
50405	:douta	=	16'h	39a7;
50406	:douta	=	16'h	2925;
50407	:douta	=	16'h	2104;
50408	:douta	=	16'h	2104;
50409	:douta	=	16'h	31ea;
50410	:douta	=	16'h	4ace;
50411	:douta	=	16'h	632f;
50412	:douta	=	16'h	4acf;
50413	:douta	=	16'h	3a6c;
50414	:douta	=	16'h	2989;
50415	:douta	=	16'h	29aa;
50416	:douta	=	16'h	10a4;
50417	:douta	=	16'h	0000;
50418	:douta	=	16'h	728a;
50419	:douta	=	16'h	7247;
50420	:douta	=	16'h	59a5;
50421	:douta	=	16'h	59e5;
50422	:douta	=	16'h	59e6;
50423	:douta	=	16'h	6a47;
50424	:douta	=	16'h	72ca;
50425	:douta	=	16'h	7b4b;
50426	:douta	=	16'h	838d;
50427	:douta	=	16'h	8c0e;
50428	:douta	=	16'h	9cb0;
50429	:douta	=	16'h	ad33;
50430	:douta	=	16'h	b554;
50431	:douta	=	16'h	bdd5;
50432	:douta	=	16'h	cdf6;
50433	:douta	=	16'h	c554;
50434	:douta	=	16'h	bd55;
50435	:douta	=	16'h	ad34;
50436	:douta	=	16'h	cdb5;
50437	:douta	=	16'h	c596;
50438	:douta	=	16'h	bd75;
50439	:douta	=	16'h	ad15;
50440	:douta	=	16'h	8c53;
50441	:douta	=	16'h	9494;
50442	:douta	=	16'h	9cb4;
50443	:douta	=	16'h	94b4;
50444	:douta	=	16'h	94d5;
50445	:douta	=	16'h	94b5;
50446	:douta	=	16'h	8454;
50447	:douta	=	16'h	8c95;
50448	:douta	=	16'h	9d17;
50449	:douta	=	16'h	73f2;
50450	:douta	=	16'h	1882;
50451	:douta	=	16'h	20c3;
50452	:douta	=	16'h	20c3;
50453	:douta	=	16'h	20c3;
50454	:douta	=	16'h	20c3;
50455	:douta	=	16'h	20e3;
50456	:douta	=	16'h	20c3;
50457	:douta	=	16'h	20a3;
50458	:douta	=	16'h	20c3;
50459	:douta	=	16'h	20c3;
50460	:douta	=	16'h	1882;
50461	:douta	=	16'h	20a2;
50462	:douta	=	16'h	1881;
50463	:douta	=	16'h	1881;
50464	:douta	=	16'h	20a2;
50465	:douta	=	16'h	20a2;
50466	:douta	=	16'h	20a2;
50467	:douta	=	16'h	28e2;
50468	:douta	=	16'h	20a2;
50469	:douta	=	16'h	20c2;
50470	:douta	=	16'h	20c2;
50471	:douta	=	16'h	28c3;
50472	:douta	=	16'h	28e2;
50473	:douta	=	16'h	28e3;
50474	:douta	=	16'h	3103;
50475	:douta	=	16'h	30e2;
50476	:douta	=	16'h	3103;
50477	:douta	=	16'h	3103;
50478	:douta	=	16'h	3902;
50479	:douta	=	16'h	4185;
50480	:douta	=	16'h	422a;
50481	:douta	=	16'h	18e4;
50482	:douta	=	16'h	4963;
50483	:douta	=	16'h	4984;
50484	:douta	=	16'h	4984;
50485	:douta	=	16'h	51a4;
50486	:douta	=	16'h	59a4;
50487	:douta	=	16'h	59c4;
50488	:douta	=	16'h	59c4;
50489	:douta	=	16'h	59c4;
50490	:douta	=	16'h	61e4;
50491	:douta	=	16'h	6a25;
50492	:douta	=	16'h	8c30;
50493	:douta	=	16'h	7ae7;
50494	:douta	=	16'h	69e3;
50495	:douta	=	16'h	7245;
50496	:douta	=	16'h	7244;
50497	:douta	=	16'h	7244;
50498	:douta	=	16'h	7a64;
50499	:douta	=	16'h	7a64;
50500	:douta	=	16'h	7a64;
50501	:douta	=	16'h	7224;
50502	:douta	=	16'h	82a4;
50503	:douta	=	16'h	82a5;
50504	:douta	=	16'h	8284;
50505	:douta	=	16'h	8285;
50506	:douta	=	16'h	8285;
50507	:douta	=	16'h	8aa5;
50508	:douta	=	16'h	82a4;
50509	:douta	=	16'h	8ac5;
50510	:douta	=	16'h	8aa4;
50511	:douta	=	16'h	8ac5;
50512	:douta	=	16'h	8ac5;
50513	:douta	=	16'h	9305;
50514	:douta	=	16'h	9305;
50515	:douta	=	16'h	9b26;
50516	:douta	=	16'h	a346;
50517	:douta	=	16'h	a325;
50518	:douta	=	16'h	a366;
50519	:douta	=	16'h	ab66;
50520	:douta	=	16'h	ab65;
50521	:douta	=	16'h	ab85;
50522	:douta	=	16'h	b3a6;
50523	:douta	=	16'h	b3c6;
50524	:douta	=	16'h	b3c6;
50525	:douta	=	16'h	bbc6;
50526	:douta	=	16'h	b3c6;
50527	:douta	=	16'h	bbe6;
50528	:douta	=	16'h	bbe5;
50529	:douta	=	16'h	bbe5;
50530	:douta	=	16'h	bbe5;
50531	:douta	=	16'h	bbe5;
50532	:douta	=	16'h	c406;
50533	:douta	=	16'h	c406;
50534	:douta	=	16'h	c406;
50535	:douta	=	16'h	c406;
50536	:douta	=	16'h	c406;
50537	:douta	=	16'h	c406;
50538	:douta	=	16'h	c427;
50539	:douta	=	16'h	c427;
50540	:douta	=	16'h	c426;
50541	:douta	=	16'h	c426;
50542	:douta	=	16'h	cc47;
50543	:douta	=	16'h	c446;
50544	:douta	=	16'h	cc47;
50545	:douta	=	16'h	c446;
50546	:douta	=	16'h	c446;
50547	:douta	=	16'h	cc67;
50548	:douta	=	16'h	c446;
50549	:douta	=	16'h	cc47;
50550	:douta	=	16'h	cc67;
50551	:douta	=	16'h	cc67;
50552	:douta	=	16'h	cc48;
50553	:douta	=	16'h	cc47;
50554	:douta	=	16'h	cc67;
50555	:douta	=	16'h	cc67;
50556	:douta	=	16'h	cc66;
50557	:douta	=	16'h	cc67;
50558	:douta	=	16'h	cc47;
50559	:douta	=	16'h	cc46;
50560	:douta	=	16'h	cc25;
50561	:douta	=	16'h	cc25;
50562	:douta	=	16'h	cc04;
50563	:douta	=	16'h	cc04;
50564	:douta	=	16'h	cc04;
50565	:douta	=	16'h	cc25;
50566	:douta	=	16'h	cc45;
50567	:douta	=	16'h	ccaa;
50568	:douta	=	16'h	d50d;
50569	:douta	=	16'h	d56f;
50570	:douta	=	16'h	de13;
50571	:douta	=	16'h	e655;
50572	:douta	=	16'h	eef8;
50573	:douta	=	16'h	ef5a;
50574	:douta	=	16'h	f79b;
50575	:douta	=	16'h	f7dc;
50576	:douta	=	16'h	fffd;
50577	:douta	=	16'h	fffd;
50578	:douta	=	16'h	fffc;
50579	:douta	=	16'h	ffdb;
50580	:douta	=	16'h	f759;
50581	:douta	=	16'h	f738;
50582	:douta	=	16'h	eef7;
50583	:douta	=	16'h	e673;
50584	:douta	=	16'h	e631;
50585	:douta	=	16'h	ddaf;
50586	:douta	=	16'h	d56c;
50587	:douta	=	16'h	d4ea;
50588	:douta	=	16'h	d4a9;
50589	:douta	=	16'h	cc87;
50590	:douta	=	16'h	cc66;
50591	:douta	=	16'h	cc46;
50592	:douta	=	16'h	cc25;
50593	:douta	=	16'h	cc46;
50594	:douta	=	16'h	cc47;
50595	:douta	=	16'h	cc68;
50596	:douta	=	16'h	d488;
50597	:douta	=	16'h	d489;
50598	:douta	=	16'h	cc88;
50599	:douta	=	16'h	d489;
50600	:douta	=	16'h	cc68;
50601	:douta	=	16'h	cc68;
50602	:douta	=	16'h	cc68;
50603	:douta	=	16'h	cc68;
50604	:douta	=	16'h	cc68;
50605	:douta	=	16'h	d466;
50606	:douta	=	16'h	c44a;
50607	:douta	=	16'h	942e;
50608	:douta	=	16'h	83cd;
50609	:douta	=	16'h	9c6f;
50610	:douta	=	16'h	a4b0;
50611	:douta	=	16'h	9c6f;
50612	:douta	=	16'h	9c8f;
50613	:douta	=	16'h	9c6f;
50614	:douta	=	16'h	acd1;
50615	:douta	=	16'h	b511;
50616	:douta	=	16'h	bd52;
50617	:douta	=	16'h	c552;
50618	:douta	=	16'h	c572;
50619	:douta	=	16'h	c593;
50620	:douta	=	16'h	de36;
50621	:douta	=	16'h	ac90;
50622	:douta	=	16'h	e697;
50623	:douta	=	16'h	acd2;
50624	:douta	=	16'h	bd33;
50625	:douta	=	16'h	b514;
50626	:douta	=	16'h	b514;
50627	:douta	=	16'h	9452;
50628	:douta	=	16'h	acd3;
50629	:douta	=	16'h	b512;
50630	:douta	=	16'h	b554;
50631	:douta	=	16'h	9453;
50632	:douta	=	16'h	ddf5;
50633	:douta	=	16'h	ddf5;
50634	:douta	=	16'h	8c74;
50635	:douta	=	16'h	9494;
50636	:douta	=	16'h	8c94;
50637	:douta	=	16'h	7c11;
50638	:douta	=	16'h	73d1;
50639	:douta	=	16'h	73d1;
50640	:douta	=	16'h	630e;
50641	:douta	=	16'h	5acd;
50642	:douta	=	16'h	5229;
50643	:douta	=	16'h	49e7;
50644	:douta	=	16'h	28e3;
50645	:douta	=	16'h	1881;
50646	:douta	=	16'h	1882;
50647	:douta	=	16'h	2103;
50648	:douta	=	16'h	3164;
50649	:douta	=	16'h	41e5;
50650	:douta	=	16'h	5a89;
50651	:douta	=	16'h	5247;
50652	:douta	=	16'h	5a68;
50653	:douta	=	16'h	5a48;
50654	:douta	=	16'h	62ea;
50655	:douta	=	16'h	730c;
50656	:douta	=	16'h	7b4c;
50657	:douta	=	16'h	83cd;
50658	:douta	=	16'h	836c;
50659	:douta	=	16'h	9c2e;
50660	:douta	=	16'h	7b6c;
50661	:douta	=	16'h	5249;
50662	:douta	=	16'h	422b;
50663	:douta	=	16'h	424b;
50664	:douta	=	16'h	3a2b;
50665	:douta	=	16'h	3a2b;
50666	:douta	=	16'h	2968;
50667	:douta	=	16'h	4a4b;
50668	:douta	=	16'h	3a2b;
50669	:douta	=	16'h	3a0b;
50670	:douta	=	16'h	2189;
50671	:douta	=	16'h	2126;
50672	:douta	=	16'h	29a8;
50673	:douta	=	16'h	0883;
50674	:douta	=	16'h	18c5;
50675	:douta	=	16'h	18e4;
50676	:douta	=	16'h	9470;
50677	:douta	=	16'h	a4b2;
50678	:douta	=	16'h	9c90;
50679	:douta	=	16'h	8c0e;
50680	:douta	=	16'h	836c;
50681	:douta	=	16'h	730a;
50682	:douta	=	16'h	72a8;
50683	:douta	=	16'h	6a68;
50684	:douta	=	16'h	6247;
50685	:douta	=	16'h	6226;
50686	:douta	=	16'h	6a26;
50687	:douta	=	16'h	6a05;
50688	:douta	=	16'h	c595;
50689	:douta	=	16'h	c575;
50690	:douta	=	16'h	b535;
50691	:douta	=	16'h	bd75;
50692	:douta	=	16'h	cdb6;
50693	:douta	=	16'h	bd95;
50694	:douta	=	16'h	bd75;
50695	:douta	=	16'h	a4f5;
50696	:douta	=	16'h	8c52;
50697	:douta	=	16'h	9473;
50698	:douta	=	16'h	a4d4;
50699	:douta	=	16'h	94b4;
50700	:douta	=	16'h	94d5;
50701	:douta	=	16'h	94d5;
50702	:douta	=	16'h	8474;
50703	:douta	=	16'h	8c95;
50704	:douta	=	16'h	94f7;
50705	:douta	=	16'h	39a7;
50706	:douta	=	16'h	20e3;
50707	:douta	=	16'h	20c3;
50708	:douta	=	16'h	20c3;
50709	:douta	=	16'h	20e3;
50710	:douta	=	16'h	20c3;
50711	:douta	=	16'h	20e3;
50712	:douta	=	16'h	20c3;
50713	:douta	=	16'h	20c3;
50714	:douta	=	16'h	20c3;
50715	:douta	=	16'h	20e3;
50716	:douta	=	16'h	1882;
50717	:douta	=	16'h	20a2;
50718	:douta	=	16'h	2082;
50719	:douta	=	16'h	1881;
50720	:douta	=	16'h	20a2;
50721	:douta	=	16'h	20a2;
50722	:douta	=	16'h	20a2;
50723	:douta	=	16'h	20a2;
50724	:douta	=	16'h	20c2;
50725	:douta	=	16'h	20a2;
50726	:douta	=	16'h	28e3;
50727	:douta	=	16'h	28c2;
50728	:douta	=	16'h	28e2;
50729	:douta	=	16'h	30e3;
50730	:douta	=	16'h	30e2;
50731	:douta	=	16'h	3103;
50732	:douta	=	16'h	3103;
50733	:douta	=	16'h	3923;
50734	:douta	=	16'h	3903;
50735	:douta	=	16'h	41a6;
50736	:douta	=	16'h	31c9;
50737	:douta	=	16'h	2905;
50738	:douta	=	16'h	4963;
50739	:douta	=	16'h	4984;
50740	:douta	=	16'h	5184;
50741	:douta	=	16'h	51a4;
50742	:douta	=	16'h	51a4;
50743	:douta	=	16'h	59a4;
50744	:douta	=	16'h	59c4;
50745	:douta	=	16'h	61c4;
50746	:douta	=	16'h	61e4;
50747	:douta	=	16'h	6a67;
50748	:douta	=	16'h	94b1;
50749	:douta	=	16'h	7285;
50750	:douta	=	16'h	69e4;
50751	:douta	=	16'h	7a65;
50752	:douta	=	16'h	7244;
50753	:douta	=	16'h	7244;
50754	:douta	=	16'h	7a64;
50755	:douta	=	16'h	7a64;
50756	:douta	=	16'h	8285;
50757	:douta	=	16'h	59c4;
50758	:douta	=	16'h	8ac5;
50759	:douta	=	16'h	8285;
50760	:douta	=	16'h	8284;
50761	:douta	=	16'h	8285;
50762	:douta	=	16'h	82a4;
50763	:douta	=	16'h	8aa5;
50764	:douta	=	16'h	82a5;
50765	:douta	=	16'h	8aa5;
50766	:douta	=	16'h	8aa4;
50767	:douta	=	16'h	8ac4;
50768	:douta	=	16'h	8ac5;
50769	:douta	=	16'h	9305;
50770	:douta	=	16'h	9305;
50771	:douta	=	16'h	9b26;
50772	:douta	=	16'h	a346;
50773	:douta	=	16'h	a346;
50774	:douta	=	16'h	a366;
50775	:douta	=	16'h	ab66;
50776	:douta	=	16'h	b385;
50777	:douta	=	16'h	b385;
50778	:douta	=	16'h	b3a6;
50779	:douta	=	16'h	b3c6;
50780	:douta	=	16'h	b3c6;
50781	:douta	=	16'h	bbc6;
50782	:douta	=	16'h	bbc6;
50783	:douta	=	16'h	bbe6;
50784	:douta	=	16'h	bbe5;
50785	:douta	=	16'h	bbe5;
50786	:douta	=	16'h	c406;
50787	:douta	=	16'h	c406;
50788	:douta	=	16'h	c406;
50789	:douta	=	16'h	c406;
50790	:douta	=	16'h	c406;
50791	:douta	=	16'h	c406;
50792	:douta	=	16'h	c406;
50793	:douta	=	16'h	c426;
50794	:douta	=	16'h	c426;
50795	:douta	=	16'h	c427;
50796	:douta	=	16'h	c427;
50797	:douta	=	16'h	c427;
50798	:douta	=	16'h	c426;
50799	:douta	=	16'h	c446;
50800	:douta	=	16'h	c426;
50801	:douta	=	16'h	cc27;
50802	:douta	=	16'h	cc47;
50803	:douta	=	16'h	c447;
50804	:douta	=	16'h	cc47;
50805	:douta	=	16'h	cc47;
50806	:douta	=	16'h	cc47;
50807	:douta	=	16'h	cc47;
50808	:douta	=	16'h	cc47;
50809	:douta	=	16'h	cc46;
50810	:douta	=	16'h	cc25;
50811	:douta	=	16'h	cc25;
50812	:douta	=	16'h	cc04;
50813	:douta	=	16'h	cbe3;
50814	:douta	=	16'h	cc24;
50815	:douta	=	16'h	cc25;
50816	:douta	=	16'h	cc69;
50817	:douta	=	16'h	ccaa;
50818	:douta	=	16'h	d52d;
50819	:douta	=	16'h	d590;
50820	:douta	=	16'h	ddd1;
50821	:douta	=	16'h	e675;
50822	:douta	=	16'h	e696;
50823	:douta	=	16'h	ef39;
50824	:douta	=	16'h	f79c;
50825	:douta	=	16'h	f7bc;
50826	:douta	=	16'h	fffd;
50827	:douta	=	16'h	fffd;
50828	:douta	=	16'h	ffbc;
50829	:douta	=	16'h	f779;
50830	:douta	=	16'h	f758;
50831	:douta	=	16'h	f6f7;
50832	:douta	=	16'h	eed5;
50833	:douta	=	16'h	e673;
50834	:douta	=	16'h	e5d0;
50835	:douta	=	16'h	ddae;
50836	:douta	=	16'h	dd4c;
50837	:douta	=	16'h	d52a;
50838	:douta	=	16'h	d4c9;
50839	:douta	=	16'h	d487;
50840	:douta	=	16'h	cc87;
50841	:douta	=	16'h	cc47;
50842	:douta	=	16'h	cc46;
50843	:douta	=	16'h	cc47;
50844	:douta	=	16'h	d488;
50845	:douta	=	16'h	d488;
50846	:douta	=	16'h	d488;
50847	:douta	=	16'h	d488;
50848	:douta	=	16'h	d488;
50849	:douta	=	16'h	cc68;
50850	:douta	=	16'h	cc88;
50851	:douta	=	16'h	d488;
50852	:douta	=	16'h	d488;
50853	:douta	=	16'h	d488;
50854	:douta	=	16'h	cc68;
50855	:douta	=	16'h	cc68;
50856	:douta	=	16'h	d467;
50857	:douta	=	16'h	d488;
50858	:douta	=	16'h	d468;
50859	:douta	=	16'h	cc67;
50860	:douta	=	16'h	cc68;
50861	:douta	=	16'h	d466;
50862	:douta	=	16'h	c46a;
50863	:douta	=	16'h	9c2f;
50864	:douta	=	16'h	8bed;
50865	:douta	=	16'h	9c70;
50866	:douta	=	16'h	a4d0;
50867	:douta	=	16'h	a490;
50868	:douta	=	16'h	a4b0;
50869	:douta	=	16'h	a4b0;
50870	:douta	=	16'h	b511;
50871	:douta	=	16'h	bd32;
50872	:douta	=	16'h	c572;
50873	:douta	=	16'h	cd93;
50874	:douta	=	16'h	cdb4;
50875	:douta	=	16'h	cdd4;
50876	:douta	=	16'h	d5f4;
50877	:douta	=	16'h	a490;
50878	:douta	=	16'h	eed7;
50879	:douta	=	16'h	cd94;
50880	:douta	=	16'h	bd54;
50881	:douta	=	16'h	9494;
50882	:douta	=	16'h	acf4;
50883	:douta	=	16'h	7bf2;
50884	:douta	=	16'h	6bb2;
50885	:douta	=	16'h	acd3;
50886	:douta	=	16'h	c574;
50887	:douta	=	16'h	a4b5;
50888	:douta	=	16'h	a4d3;
50889	:douta	=	16'h	bd55;
50890	:douta	=	16'h	8c74;
50891	:douta	=	16'h	8453;
50892	:douta	=	16'h	8433;
50893	:douta	=	16'h	6bb1;
50894	:douta	=	16'h	6bd1;
50895	:douta	=	16'h	6b0d;
50896	:douta	=	16'h	4a08;
50897	:douta	=	16'h	39a5;
50898	:douta	=	16'h	2902;
50899	:douta	=	16'h	20e1;
50900	:douta	=	16'h	28e3;
50901	:douta	=	16'h	3965;
50902	:douta	=	16'h	3985;
50903	:douta	=	16'h	3985;
50904	:douta	=	16'h	39a5;
50905	:douta	=	16'h	4a06;
50906	:douta	=	16'h	5247;
50907	:douta	=	16'h	6ac9;
50908	:douta	=	16'h	6aea;
50909	:douta	=	16'h	730b;
50910	:douta	=	16'h	736c;
50911	:douta	=	16'h	7b8d;
50912	:douta	=	16'h	83cd;
50913	:douta	=	16'h	940f;
50914	:douta	=	16'h	8bed;
50915	:douta	=	16'h	9c4e;
50916	:douta	=	16'h	9c2f;
50917	:douta	=	16'h	838d;
50918	:douta	=	16'h	2967;
50919	:douta	=	16'h	2146;
50920	:douta	=	16'h	10c4;
50921	:douta	=	16'h	1905;
50922	:douta	=	16'h	10e5;
50923	:douta	=	16'h	2967;
50924	:douta	=	16'h	1906;
50925	:douta	=	16'h	2987;
50926	:douta	=	16'h	29a9;
50927	:douta	=	16'h	2147;
50928	:douta	=	16'h	2967;
50929	:douta	=	16'h	1905;
50930	:douta	=	16'h	10e6;
50931	:douta	=	16'h	08a5;
50932	:douta	=	16'h	39a6;
50933	:douta	=	16'h	6267;
50934	:douta	=	16'h	6266;
50935	:douta	=	16'h	6246;
50936	:douta	=	16'h	6226;
50937	:douta	=	16'h	6a26;
50938	:douta	=	16'h	6a26;
50939	:douta	=	16'h	6a46;
50940	:douta	=	16'h	7266;
50941	:douta	=	16'h	7267;
50942	:douta	=	16'h	7267;
50943	:douta	=	16'h	7287;
50944	:douta	=	16'h	b514;
50945	:douta	=	16'h	b555;
50946	:douta	=	16'h	a4f5;
50947	:douta	=	16'h	cdb6;
50948	:douta	=	16'h	c595;
50949	:douta	=	16'h	bd75;
50950	:douta	=	16'h	ad35;
50951	:douta	=	16'h	94b4;
50952	:douta	=	16'h	9c94;
50953	:douta	=	16'h	9cb4;
50954	:douta	=	16'h	a4f5;
50955	:douta	=	16'h	94d5;
50956	:douta	=	16'h	9cd6;
50957	:douta	=	16'h	8cb5;
50958	:douta	=	16'h	8c74;
50959	:douta	=	16'h	9d17;
50960	:douta	=	16'h	18a2;
50961	:douta	=	16'h	2061;
50962	:douta	=	16'h	28e3;
50963	:douta	=	16'h	20e3;
50964	:douta	=	16'h	20e3;
50965	:douta	=	16'h	20c3;
50966	:douta	=	16'h	20c3;
50967	:douta	=	16'h	20e3;
50968	:douta	=	16'h	20c3;
50969	:douta	=	16'h	20a3;
50970	:douta	=	16'h	20e3;
50971	:douta	=	16'h	20c3;
50972	:douta	=	16'h	2082;
50973	:douta	=	16'h	2082;
50974	:douta	=	16'h	2082;
50975	:douta	=	16'h	20a2;
50976	:douta	=	16'h	20a2;
50977	:douta	=	16'h	20a2;
50978	:douta	=	16'h	2082;
50979	:douta	=	16'h	20a2;
50980	:douta	=	16'h	20c2;
50981	:douta	=	16'h	20c2;
50982	:douta	=	16'h	20c2;
50983	:douta	=	16'h	28e2;
50984	:douta	=	16'h	28e2;
50985	:douta	=	16'h	30e2;
50986	:douta	=	16'h	3103;
50987	:douta	=	16'h	30e3;
50988	:douta	=	16'h	3103;
50989	:douta	=	16'h	3903;
50990	:douta	=	16'h	3923;
50991	:douta	=	16'h	4209;
50992	:douta	=	16'h	2988;
50993	:douta	=	16'h	3903;
50994	:douta	=	16'h	5164;
50995	:douta	=	16'h	51a4;
50996	:douta	=	16'h	51a4;
50997	:douta	=	16'h	51a3;
50998	:douta	=	16'h	59c4;
50999	:douta	=	16'h	59a4;
51000	:douta	=	16'h	61e4;
51001	:douta	=	16'h	61e4;
51002	:douta	=	16'h	61e4;
51003	:douta	=	16'h	6ac9;
51004	:douta	=	16'h	ad53;
51005	:douta	=	16'h	6a03;
51006	:douta	=	16'h	7245;
51007	:douta	=	16'h	7244;
51008	:douta	=	16'h	7244;
51009	:douta	=	16'h	7a44;
51010	:douta	=	16'h	7a44;
51011	:douta	=	16'h	7a64;
51012	:douta	=	16'h	8284;
51013	:douta	=	16'h	51c4;
51014	:douta	=	16'h	7244;
51015	:douta	=	16'h	8285;
51016	:douta	=	16'h	8285;
51017	:douta	=	16'h	82a5;
51018	:douta	=	16'h	82a4;
51019	:douta	=	16'h	8ac5;
51020	:douta	=	16'h	8ac5;
51021	:douta	=	16'h	8ac5;
51022	:douta	=	16'h	8ac5;
51023	:douta	=	16'h	8ac5;
51024	:douta	=	16'h	8ac5;
51025	:douta	=	16'h	9305;
51026	:douta	=	16'h	9b26;
51027	:douta	=	16'h	a326;
51028	:douta	=	16'h	a346;
51029	:douta	=	16'h	a346;
51030	:douta	=	16'h	ab86;
51031	:douta	=	16'h	aba6;
51032	:douta	=	16'h	b385;
51033	:douta	=	16'h	b3a5;
51034	:douta	=	16'h	b3a5;
51035	:douta	=	16'h	b3c6;
51036	:douta	=	16'h	bbc6;
51037	:douta	=	16'h	bbc6;
51038	:douta	=	16'h	bbc6;
51039	:douta	=	16'h	bbe6;
51040	:douta	=	16'h	bbe6;
51041	:douta	=	16'h	bbe6;
51042	:douta	=	16'h	c406;
51043	:douta	=	16'h	bc05;
51044	:douta	=	16'h	c406;
51045	:douta	=	16'h	c406;
51046	:douta	=	16'h	c406;
51047	:douta	=	16'h	c426;
51048	:douta	=	16'h	c426;
51049	:douta	=	16'h	c427;
51050	:douta	=	16'h	c426;
51051	:douta	=	16'h	c425;
51052	:douta	=	16'h	c405;
51053	:douta	=	16'h	c405;
51054	:douta	=	16'h	c404;
51055	:douta	=	16'h	c3e3;
51056	:douta	=	16'h	c3e3;
51057	:douta	=	16'h	c404;
51058	:douta	=	16'h	c405;
51059	:douta	=	16'h	c447;
51060	:douta	=	16'h	cc6a;
51061	:douta	=	16'h	cccb;
51062	:douta	=	16'h	d54e;
51063	:douta	=	16'h	ddb0;
51064	:douta	=	16'h	de34;
51065	:douta	=	16'h	e6d7;
51066	:douta	=	16'h	eef8;
51067	:douta	=	16'h	f77b;
51068	:douta	=	16'h	f7bb;
51069	:douta	=	16'h	ffdc;
51070	:douta	=	16'h	fffd;
51071	:douta	=	16'h	ffdc;
51072	:douta	=	16'h	ff9a;
51073	:douta	=	16'h	f759;
51074	:douta	=	16'h	ef16;
51075	:douta	=	16'h	e694;
51076	:douta	=	16'h	e653;
51077	:douta	=	16'h	ddd0;
51078	:douta	=	16'h	ddae;
51079	:douta	=	16'h	d52b;
51080	:douta	=	16'h	d4ca;
51081	:douta	=	16'h	d489;
51082	:douta	=	16'h	cc87;
51083	:douta	=	16'h	cc45;
51084	:douta	=	16'h	cc46;
51085	:douta	=	16'h	cc46;
51086	:douta	=	16'h	cc46;
51087	:douta	=	16'h	cc47;
51088	:douta	=	16'h	cc67;
51089	:douta	=	16'h	d467;
51090	:douta	=	16'h	d467;
51091	:douta	=	16'h	d467;
51092	:douta	=	16'h	d488;
51093	:douta	=	16'h	cc87;
51094	:douta	=	16'h	d487;
51095	:douta	=	16'h	d488;
51096	:douta	=	16'h	cc88;
51097	:douta	=	16'h	d488;
51098	:douta	=	16'h	d488;
51099	:douta	=	16'h	d488;
51100	:douta	=	16'h	d488;
51101	:douta	=	16'h	cc88;
51102	:douta	=	16'h	cc88;
51103	:douta	=	16'h	cc88;
51104	:douta	=	16'h	d488;
51105	:douta	=	16'h	d488;
51106	:douta	=	16'h	d488;
51107	:douta	=	16'h	cc88;
51108	:douta	=	16'h	d488;
51109	:douta	=	16'h	d488;
51110	:douta	=	16'h	cc68;
51111	:douta	=	16'h	cc88;
51112	:douta	=	16'h	cc67;
51113	:douta	=	16'h	cc67;
51114	:douta	=	16'h	cc68;
51115	:douta	=	16'h	cc68;
51116	:douta	=	16'h	cc68;
51117	:douta	=	16'h	d467;
51118	:douta	=	16'h	cc68;
51119	:douta	=	16'h	9c70;
51120	:douta	=	16'h	9c50;
51121	:douta	=	16'h	9c2f;
51122	:douta	=	16'h	9c70;
51123	:douta	=	16'h	a4b0;
51124	:douta	=	16'h	b511;
51125	:douta	=	16'h	bd31;
51126	:douta	=	16'h	bd72;
51127	:douta	=	16'h	cd94;
51128	:douta	=	16'h	cdb4;
51129	:douta	=	16'h	cdd4;
51130	:douta	=	16'h	d5f5;
51131	:douta	=	16'h	d5f5;
51132	:douta	=	16'h	cd93;
51133	:douta	=	16'h	b4d2;
51134	:douta	=	16'h	b4f3;
51135	:douta	=	16'h	acf4;
51136	:douta	=	16'h	c555;
51137	:douta	=	16'h	bd74;
51138	:douta	=	16'h	94b4;
51139	:douta	=	16'h	8c74;
51140	:douta	=	16'h	73d1;
51141	:douta	=	16'h	73f2;
51142	:douta	=	16'h	6bb2;
51143	:douta	=	16'h	8433;
51144	:douta	=	16'h	73d2;
51145	:douta	=	16'h	6370;
51146	:douta	=	16'h	6b91;
51147	:douta	=	16'h	4a6a;
51148	:douta	=	16'h	39c7;
51149	:douta	=	16'h	18a3;
51150	:douta	=	16'h	1881;
51151	:douta	=	16'h	2923;
51152	:douta	=	16'h	3965;
51153	:douta	=	16'h	3145;
51154	:douta	=	16'h	41c5;
51155	:douta	=	16'h	5227;
51156	:douta	=	16'h	5207;
51157	:douta	=	16'h	732a;
51158	:douta	=	16'h	6b0a;
51159	:douta	=	16'h	6ac9;
51160	:douta	=	16'h	6ae9;
51161	:douta	=	16'h	734b;
51162	:douta	=	16'h	734b;
51163	:douta	=	16'h	7b4b;
51164	:douta	=	16'h	7b4b;
51165	:douta	=	16'h	7b6b;
51166	:douta	=	16'h	9c4f;
51167	:douta	=	16'h	a46f;
51168	:douta	=	16'h	acaf;
51169	:douta	=	16'h	ac8f;
51170	:douta	=	16'h	b4d0;
51171	:douta	=	16'h	a46f;
51172	:douta	=	16'h	9c6f;
51173	:douta	=	16'h	8bee;
51174	:douta	=	16'h	62ed;
51175	:douta	=	16'h	3a2b;
51176	:douta	=	16'h	2967;
51177	:douta	=	16'h	18e5;
51178	:douta	=	16'h	10c3;
51179	:douta	=	16'h	0882;
51180	:douta	=	16'h	08c3;
51181	:douta	=	16'h	10a4;
51182	:douta	=	16'h	10a4;
51183	:douta	=	16'h	10e5;
51184	:douta	=	16'h	2147;
51185	:douta	=	16'h	2167;
51186	:douta	=	16'h	1906;
51187	:douta	=	16'h	1948;
51188	:douta	=	16'h	1905;
51189	:douta	=	16'h	82a7;
51190	:douta	=	16'h	7267;
51191	:douta	=	16'h	7286;
51192	:douta	=	16'h	7a67;
51193	:douta	=	16'h	7a67;
51194	:douta	=	16'h	7a87;
51195	:douta	=	16'h	7a87;
51196	:douta	=	16'h	7a87;
51197	:douta	=	16'h	7a87;
51198	:douta	=	16'h	7a86;
51199	:douta	=	16'h	7a87;
51200	:douta	=	16'h	b513;
51201	:douta	=	16'h	b515;
51202	:douta	=	16'h	a4f5;
51203	:douta	=	16'h	cdf6;
51204	:douta	=	16'h	bd75;
51205	:douta	=	16'h	bd75;
51206	:douta	=	16'h	a4f4;
51207	:douta	=	16'h	8c73;
51208	:douta	=	16'h	a4d5;
51209	:douta	=	16'h	a4d5;
51210	:douta	=	16'h	a4d5;
51211	:douta	=	16'h	94d5;
51212	:douta	=	16'h	9cd6;
51213	:douta	=	16'h	8474;
51214	:douta	=	16'h	8474;
51215	:douta	=	16'h	a559;
51216	:douta	=	16'h	1040;
51217	:douta	=	16'h	28e3;
51218	:douta	=	16'h	20c3;
51219	:douta	=	16'h	20e3;
51220	:douta	=	16'h	20c3;
51221	:douta	=	16'h	20e3;
51222	:douta	=	16'h	20e3;
51223	:douta	=	16'h	20c3;
51224	:douta	=	16'h	20a3;
51225	:douta	=	16'h	20c3;
51226	:douta	=	16'h	20e3;
51227	:douta	=	16'h	20e3;
51228	:douta	=	16'h	2082;
51229	:douta	=	16'h	20a2;
51230	:douta	=	16'h	20a2;
51231	:douta	=	16'h	2082;
51232	:douta	=	16'h	20a2;
51233	:douta	=	16'h	20a2;
51234	:douta	=	16'h	20a2;
51235	:douta	=	16'h	20a2;
51236	:douta	=	16'h	20c2;
51237	:douta	=	16'h	20c2;
51238	:douta	=	16'h	28e2;
51239	:douta	=	16'h	28e2;
51240	:douta	=	16'h	28e2;
51241	:douta	=	16'h	30e2;
51242	:douta	=	16'h	30e3;
51243	:douta	=	16'h	30e3;
51244	:douta	=	16'h	3103;
51245	:douta	=	16'h	3923;
51246	:douta	=	16'h	3924;
51247	:douta	=	16'h	422a;
51248	:douta	=	16'h	1926;
51249	:douta	=	16'h	4144;
51250	:douta	=	16'h	5184;
51251	:douta	=	16'h	5184;
51252	:douta	=	16'h	5184;
51253	:douta	=	16'h	51a4;
51254	:douta	=	16'h	59c4;
51255	:douta	=	16'h	59c4;
51256	:douta	=	16'h	61c3;
51257	:douta	=	16'h	61e4;
51258	:douta	=	16'h	6a04;
51259	:douta	=	16'h	732b;
51260	:douta	=	16'h	b595;
51261	:douta	=	16'h	69c3;
51262	:douta	=	16'h	7224;
51263	:douta	=	16'h	7244;
51264	:douta	=	16'h	7a44;
51265	:douta	=	16'h	7245;
51266	:douta	=	16'h	7a65;
51267	:douta	=	16'h	7a84;
51268	:douta	=	16'h	7a64;
51269	:douta	=	16'h	6a24;
51270	:douta	=	16'h	6a44;
51271	:douta	=	16'h	8284;
51272	:douta	=	16'h	8285;
51273	:douta	=	16'h	82a5;
51274	:douta	=	16'h	8aa4;
51275	:douta	=	16'h	8ac5;
51276	:douta	=	16'h	8aa4;
51277	:douta	=	16'h	8ac5;
51278	:douta	=	16'h	92e5;
51279	:douta	=	16'h	8ac5;
51280	:douta	=	16'h	8ac5;
51281	:douta	=	16'h	9305;
51282	:douta	=	16'h	9305;
51283	:douta	=	16'h	9b26;
51284	:douta	=	16'h	a346;
51285	:douta	=	16'h	a366;
51286	:douta	=	16'h	ab86;
51287	:douta	=	16'h	ab66;
51288	:douta	=	16'h	b3a5;
51289	:douta	=	16'h	b3a5;
51290	:douta	=	16'h	b3a6;
51291	:douta	=	16'h	b3c6;
51292	:douta	=	16'h	bbc6;
51293	:douta	=	16'h	bbc6;
51294	:douta	=	16'h	bbe6;
51295	:douta	=	16'h	bbe6;
51296	:douta	=	16'h	bbe6;
51297	:douta	=	16'h	bbe6;
51298	:douta	=	16'h	bc05;
51299	:douta	=	16'h	bbe5;
51300	:douta	=	16'h	c3e7;
51301	:douta	=	16'h	c3e6;
51302	:douta	=	16'h	c3e5;
51303	:douta	=	16'h	c3c4;
51304	:douta	=	16'h	bbc3;
51305	:douta	=	16'h	c3c3;
51306	:douta	=	16'h	c3c3;
51307	:douta	=	16'h	c3e4;
51308	:douta	=	16'h	c427;
51309	:douta	=	16'h	c448;
51310	:douta	=	16'h	ccaa;
51311	:douta	=	16'h	d52e;
51312	:douta	=	16'h	d56f;
51313	:douta	=	16'h	ddf2;
51314	:douta	=	16'h	de13;
51315	:douta	=	16'h	e696;
51316	:douta	=	16'h	ef19;
51317	:douta	=	16'h	f77a;
51318	:douta	=	16'h	f7bc;
51319	:douta	=	16'h	f7bd;
51320	:douta	=	16'h	ffdc;
51321	:douta	=	16'h	f79b;
51322	:douta	=	16'h	f77a;
51323	:douta	=	16'h	ef17;
51324	:douta	=	16'h	eef6;
51325	:douta	=	16'h	e694;
51326	:douta	=	16'h	ddf0;
51327	:douta	=	16'h	ddcf;
51328	:douta	=	16'h	d54c;
51329	:douta	=	16'h	d50b;
51330	:douta	=	16'h	cca9;
51331	:douta	=	16'h	d487;
51332	:douta	=	16'h	cc67;
51333	:douta	=	16'h	cc25;
51334	:douta	=	16'h	cc25;
51335	:douta	=	16'h	cc46;
51336	:douta	=	16'h	cc46;
51337	:douta	=	16'h	d467;
51338	:douta	=	16'h	d467;
51339	:douta	=	16'h	cc68;
51340	:douta	=	16'h	cc88;
51341	:douta	=	16'h	d488;
51342	:douta	=	16'h	cc87;
51343	:douta	=	16'h	cc87;
51344	:douta	=	16'h	d487;
51345	:douta	=	16'h	cc87;
51346	:douta	=	16'h	d487;
51347	:douta	=	16'h	d487;
51348	:douta	=	16'h	d488;
51349	:douta	=	16'h	d488;
51350	:douta	=	16'h	d488;
51351	:douta	=	16'h	cc88;
51352	:douta	=	16'h	cc88;
51353	:douta	=	16'h	d488;
51354	:douta	=	16'h	cc88;
51355	:douta	=	16'h	d488;
51356	:douta	=	16'h	d488;
51357	:douta	=	16'h	d488;
51358	:douta	=	16'h	cc88;
51359	:douta	=	16'h	d488;
51360	:douta	=	16'h	cc88;
51361	:douta	=	16'h	d488;
51362	:douta	=	16'h	d488;
51363	:douta	=	16'h	cc88;
51364	:douta	=	16'h	cc68;
51365	:douta	=	16'h	cc88;
51366	:douta	=	16'h	cc68;
51367	:douta	=	16'h	d488;
51368	:douta	=	16'h	cc67;
51369	:douta	=	16'h	d467;
51370	:douta	=	16'h	d468;
51371	:douta	=	16'h	cc69;
51372	:douta	=	16'h	cc67;
51373	:douta	=	16'h	cc68;
51374	:douta	=	16'h	d466;
51375	:douta	=	16'h	9c91;
51376	:douta	=	16'h	9c2f;
51377	:douta	=	16'h	9c6f;
51378	:douta	=	16'h	a490;
51379	:douta	=	16'h	a4b0;
51380	:douta	=	16'h	bd32;
51381	:douta	=	16'h	bd53;
51382	:douta	=	16'h	c573;
51383	:douta	=	16'h	cdd4;
51384	:douta	=	16'h	cdb4;
51385	:douta	=	16'h	d5f5;
51386	:douta	=	16'h	d5f4;
51387	:douta	=	16'h	cdb4;
51388	:douta	=	16'h	c553;
51389	:douta	=	16'h	b4d2;
51390	:douta	=	16'h	9473;
51391	:douta	=	16'h	7c13;
51392	:douta	=	16'h	a4d4;
51393	:douta	=	16'h	bd75;
51394	:douta	=	16'h	ad16;
51395	:douta	=	16'h	7bf3;
51396	:douta	=	16'h	73d2;
51397	:douta	=	16'h	6bd2;
51398	:douta	=	16'h	73d2;
51399	:douta	=	16'h	6b4f;
51400	:douta	=	16'h	6b4f;
51401	:douta	=	16'h	5acd;
51402	:douta	=	16'h	3186;
51403	:douta	=	16'h	2903;
51404	:douta	=	16'h	28e3;
51405	:douta	=	16'h	3185;
51406	:douta	=	16'h	39a5;
51407	:douta	=	16'h	62a9;
51408	:douta	=	16'h	5a68;
51409	:douta	=	16'h	5a68;
51410	:douta	=	16'h	5227;
51411	:douta	=	16'h	5a47;
51412	:douta	=	16'h	4a06;
51413	:douta	=	16'h	732b;
51414	:douta	=	16'h	83ac;
51415	:douta	=	16'h	836c;
51416	:douta	=	16'h	7b2b;
51417	:douta	=	16'h	838c;
51418	:douta	=	16'h	8bcb;
51419	:douta	=	16'h	93ec;
51420	:douta	=	16'h	a44e;
51421	:douta	=	16'h	942d;
51422	:douta	=	16'h	a46f;
51423	:douta	=	16'h	accf;
51424	:douta	=	16'h	b510;
51425	:douta	=	16'h	c551;
51426	:douta	=	16'h	bd30;
51427	:douta	=	16'h	ac8f;
51428	:douta	=	16'h	9c2f;
51429	:douta	=	16'h	8bce;
51430	:douta	=	16'h	6b4d;
51431	:douta	=	16'h	52ac;
51432	:douta	=	16'h	3209;
51433	:douta	=	16'h	2967;
51434	:douta	=	16'h	2126;
51435	:douta	=	16'h	10a3;
51436	:douta	=	16'h	1083;
51437	:douta	=	16'h	0882;
51438	:douta	=	16'h	10c3;
51439	:douta	=	16'h	10e4;
51440	:douta	=	16'h	1927;
51441	:douta	=	16'h	2168;
51442	:douta	=	16'h	08a4;
51443	:douta	=	16'h	2188;
51444	:douta	=	16'h	08e6;
51445	:douta	=	16'h	8ac7;
51446	:douta	=	16'h	7267;
51447	:douta	=	16'h	7a87;
51448	:douta	=	16'h	8287;
51449	:douta	=	16'h	7aa7;
51450	:douta	=	16'h	7a87;
51451	:douta	=	16'h	7a87;
51452	:douta	=	16'h	82a7;
51453	:douta	=	16'h	7a87;
51454	:douta	=	16'h	7a87;
51455	:douta	=	16'h	7aa7;
51456	:douta	=	16'h	c575;
51457	:douta	=	16'h	acf5;
51458	:douta	=	16'h	ad35;
51459	:douta	=	16'h	cdf6;
51460	:douta	=	16'h	c575;
51461	:douta	=	16'h	bd75;
51462	:douta	=	16'h	9474;
51463	:douta	=	16'h	8412;
51464	:douta	=	16'h	a516;
51465	:douta	=	16'h	a4f5;
51466	:douta	=	16'h	9cd5;
51467	:douta	=	16'h	94d5;
51468	:douta	=	16'h	9cf6;
51469	:douta	=	16'h	8454;
51470	:douta	=	16'h	9cf7;
51471	:douta	=	16'h	8453;
51472	:douta	=	16'h	20a2;
51473	:douta	=	16'h	20e3;
51474	:douta	=	16'h	20e3;
51475	:douta	=	16'h	20c3;
51476	:douta	=	16'h	28e3;
51477	:douta	=	16'h	20c3;
51478	:douta	=	16'h	20e3;
51479	:douta	=	16'h	20e3;
51480	:douta	=	16'h	20c3;
51481	:douta	=	16'h	20c3;
51482	:douta	=	16'h	20e3;
51483	:douta	=	16'h	1882;
51484	:douta	=	16'h	2082;
51485	:douta	=	16'h	20a2;
51486	:douta	=	16'h	20a2;
51487	:douta	=	16'h	20a2;
51488	:douta	=	16'h	20a2;
51489	:douta	=	16'h	20a2;
51490	:douta	=	16'h	20a2;
51491	:douta	=	16'h	20c2;
51492	:douta	=	16'h	20c2;
51493	:douta	=	16'h	28e3;
51494	:douta	=	16'h	28c2;
51495	:douta	=	16'h	28e2;
51496	:douta	=	16'h	28e2;
51497	:douta	=	16'h	3103;
51498	:douta	=	16'h	3103;
51499	:douta	=	16'h	3103;
51500	:douta	=	16'h	3923;
51501	:douta	=	16'h	3923;
51502	:douta	=	16'h	41a5;
51503	:douta	=	16'h	424b;
51504	:douta	=	16'h	10e5;
51505	:douta	=	16'h	5184;
51506	:douta	=	16'h	4984;
51507	:douta	=	16'h	5184;
51508	:douta	=	16'h	5184;
51509	:douta	=	16'h	51a4;
51510	:douta	=	16'h	59c4;
51511	:douta	=	16'h	61c4;
51512	:douta	=	16'h	61e4;
51513	:douta	=	16'h	61e4;
51514	:douta	=	16'h	61c3;
51515	:douta	=	16'h	8c2f;
51516	:douta	=	16'h	b573;
51517	:douta	=	16'h	71e3;
51518	:douta	=	16'h	7245;
51519	:douta	=	16'h	7244;
51520	:douta	=	16'h	7a64;
51521	:douta	=	16'h	7a64;
51522	:douta	=	16'h	7a64;
51523	:douta	=	16'h	7a64;
51524	:douta	=	16'h	7a85;
51525	:douta	=	16'h	7a85;
51526	:douta	=	16'h	51c4;
51527	:douta	=	16'h	8aa5;
51528	:douta	=	16'h	8285;
51529	:douta	=	16'h	8284;
51530	:douta	=	16'h	8aa5;
51531	:douta	=	16'h	8aa5;
51532	:douta	=	16'h	8ac5;
51533	:douta	=	16'h	8ac5;
51534	:douta	=	16'h	8ac5;
51535	:douta	=	16'h	8ac5;
51536	:douta	=	16'h	92e6;
51537	:douta	=	16'h	9306;
51538	:douta	=	16'h	9b26;
51539	:douta	=	16'h	9b26;
51540	:douta	=	16'h	a346;
51541	:douta	=	16'h	a345;
51542	:douta	=	16'h	ab85;
51543	:douta	=	16'h	ab85;
51544	:douta	=	16'h	b385;
51545	:douta	=	16'h	ab65;
51546	:douta	=	16'h	ab64;
51547	:douta	=	16'h	b384;
51548	:douta	=	16'h	b364;
51549	:douta	=	16'h	b364;
51550	:douta	=	16'h	b364;
51551	:douta	=	16'h	bbc6;
51552	:douta	=	16'h	c428;
51553	:douta	=	16'h	c44a;
51554	:douta	=	16'h	c4ec;
51555	:douta	=	16'h	cd2d;
51556	:douta	=	16'h	d5b0;
51557	:douta	=	16'h	de54;
51558	:douta	=	16'h	e6b5;
51559	:douta	=	16'h	ef18;
51560	:douta	=	16'h	f75a;
51561	:douta	=	16'h	f79b;
51562	:douta	=	16'h	f7bc;
51563	:douta	=	16'h	f7bb;
51564	:douta	=	16'h	f779;
51565	:douta	=	16'h	ef58;
51566	:douta	=	16'h	eef6;
51567	:douta	=	16'h	e694;
51568	:douta	=	16'h	e652;
51569	:douta	=	16'h	ddcf;
51570	:douta	=	16'h	d58e;
51571	:douta	=	16'h	d50b;
51572	:douta	=	16'h	cca8;
51573	:douta	=	16'h	cc87;
51574	:douta	=	16'h	cc46;
51575	:douta	=	16'h	cc27;
51576	:douta	=	16'h	cc25;
51577	:douta	=	16'h	cc25;
51578	:douta	=	16'h	cc25;
51579	:douta	=	16'h	cc46;
51580	:douta	=	16'h	cc46;
51581	:douta	=	16'h	cc47;
51582	:douta	=	16'h	d467;
51583	:douta	=	16'h	d468;
51584	:douta	=	16'h	cc68;
51585	:douta	=	16'h	cc68;
51586	:douta	=	16'h	cc67;
51587	:douta	=	16'h	cc68;
51588	:douta	=	16'h	cc67;
51589	:douta	=	16'h	d488;
51590	:douta	=	16'h	cc67;
51591	:douta	=	16'h	d488;
51592	:douta	=	16'h	d488;
51593	:douta	=	16'h	d488;
51594	:douta	=	16'h	cc68;
51595	:douta	=	16'h	d488;
51596	:douta	=	16'h	d488;
51597	:douta	=	16'h	d488;
51598	:douta	=	16'h	d488;
51599	:douta	=	16'h	d488;
51600	:douta	=	16'h	d488;
51601	:douta	=	16'h	d487;
51602	:douta	=	16'h	cc68;
51603	:douta	=	16'h	d488;
51604	:douta	=	16'h	cc87;
51605	:douta	=	16'h	cc67;
51606	:douta	=	16'h	cc88;
51607	:douta	=	16'h	cc88;
51608	:douta	=	16'h	d488;
51609	:douta	=	16'h	d488;
51610	:douta	=	16'h	d488;
51611	:douta	=	16'h	d488;
51612	:douta	=	16'h	cc88;
51613	:douta	=	16'h	d488;
51614	:douta	=	16'h	d468;
51615	:douta	=	16'h	cc68;
51616	:douta	=	16'h	d4a9;
51617	:douta	=	16'h	cc88;
51618	:douta	=	16'h	cc68;
51619	:douta	=	16'h	d488;
51620	:douta	=	16'h	d488;
51621	:douta	=	16'h	d488;
51622	:douta	=	16'h	cc68;
51623	:douta	=	16'h	d488;
51624	:douta	=	16'h	cc68;
51625	:douta	=	16'h	d488;
51626	:douta	=	16'h	cc68;
51627	:douta	=	16'h	cc68;
51628	:douta	=	16'h	d488;
51629	:douta	=	16'h	d467;
51630	:douta	=	16'h	cc47;
51631	:douta	=	16'h	9c4e;
51632	:douta	=	16'h	9c4f;
51633	:douta	=	16'h	acd2;
51634	:douta	=	16'h	acd1;
51635	:douta	=	16'h	b4f2;
51636	:douta	=	16'h	bd32;
51637	:douta	=	16'h	bd52;
51638	:douta	=	16'h	c573;
51639	:douta	=	16'h	c594;
51640	:douta	=	16'h	c553;
51641	:douta	=	16'h	acf4;
51642	:douta	=	16'h	a4b3;
51643	:douta	=	16'h	9473;
51644	:douta	=	16'h	7bf2;
51645	:douta	=	16'h	8432;
51646	:douta	=	16'h	8c53;
51647	:douta	=	16'h	6bb1;
51648	:douta	=	16'h	7c13;
51649	:douta	=	16'h	6bb1;
51650	:douta	=	16'h	7391;
51651	:douta	=	16'h	736f;
51652	:douta	=	16'h	62cd;
51653	:douta	=	16'h	39a6;
51654	:douta	=	16'h	3144;
51655	:douta	=	16'h	3124;
51656	:douta	=	16'h	2902;
51657	:douta	=	16'h	0860;
51658	:douta	=	16'h	8bcd;
51659	:douta	=	16'h	62ca;
51660	:douta	=	16'h	6b0a;
51661	:douta	=	16'h	7b6b;
51662	:douta	=	16'h	940e;
51663	:douta	=	16'h	8bad;
51664	:douta	=	16'h	940e;
51665	:douta	=	16'h	83ad;
51666	:douta	=	16'h	8bed;
51667	:douta	=	16'h	838c;
51668	:douta	=	16'h	8bcc;
51669	:douta	=	16'h	7b6b;
51670	:douta	=	16'h	7309;
51671	:douta	=	16'h	9c2e;
51672	:douta	=	16'h	9c6f;
51673	:douta	=	16'h	ac8f;
51674	:douta	=	16'h	b4d0;
51675	:douta	=	16'h	b510;
51676	:douta	=	16'h	c551;
51677	:douta	=	16'h	cd71;
51678	:douta	=	16'h	cd92;
51679	:douta	=	16'h	cd72;
51680	:douta	=	16'h	bd12;
51681	:douta	=	16'h	c551;
51682	:douta	=	16'h	cd92;
51683	:douta	=	16'h	ac8f;
51684	:douta	=	16'h	a470;
51685	:douta	=	16'h	9410;
51686	:douta	=	16'h	736e;
51687	:douta	=	16'h	632d;
51688	:douta	=	16'h	424b;
51689	:douta	=	16'h	31a8;
51690	:douta	=	16'h	31c8;
51691	:douta	=	16'h	2126;
51692	:douta	=	16'h	1905;
51693	:douta	=	16'h	2987;
51694	:douta	=	16'h	0883;
51695	:douta	=	16'h	10c4;
51696	:douta	=	16'h	1083;
51697	:douta	=	16'h	10c4;
51698	:douta	=	16'h	10e5;
51699	:douta	=	16'h	2169;
51700	:douta	=	16'h	2188;
51701	:douta	=	16'h	59e6;
51702	:douta	=	16'h	8ae8;
51703	:douta	=	16'h	7aa6;
51704	:douta	=	16'h	82a7;
51705	:douta	=	16'h	82a7;
51706	:douta	=	16'h	82a7;
51707	:douta	=	16'h	82a7;
51708	:douta	=	16'h	82a7;
51709	:douta	=	16'h	82a7;
51710	:douta	=	16'h	82a7;
51711	:douta	=	16'h	82a7;
51712	:douta	=	16'h	bd75;
51713	:douta	=	16'h	ad15;
51714	:douta	=	16'h	bd75;
51715	:douta	=	16'h	cdd6;
51716	:douta	=	16'h	c575;
51717	:douta	=	16'h	bd75;
51718	:douta	=	16'h	8c32;
51719	:douta	=	16'h	8c73;
51720	:douta	=	16'h	94b5;
51721	:douta	=	16'h	a4f5;
51722	:douta	=	16'h	9cd5;
51723	:douta	=	16'h	9cf6;
51724	:douta	=	16'h	94d5;
51725	:douta	=	16'h	8454;
51726	:douta	=	16'h	a579;
51727	:douta	=	16'h	5b0c;
51728	:douta	=	16'h	28e3;
51729	:douta	=	16'h	28e4;
51730	:douta	=	16'h	20c3;
51731	:douta	=	16'h	28e3;
51732	:douta	=	16'h	20a3;
51733	:douta	=	16'h	20e3;
51734	:douta	=	16'h	20c3;
51735	:douta	=	16'h	20e3;
51736	:douta	=	16'h	20c3;
51737	:douta	=	16'h	20a3;
51738	:douta	=	16'h	20e3;
51739	:douta	=	16'h	1882;
51740	:douta	=	16'h	20a2;
51741	:douta	=	16'h	1881;
51742	:douta	=	16'h	1881;
51743	:douta	=	16'h	20a2;
51744	:douta	=	16'h	20a2;
51745	:douta	=	16'h	20a2;
51746	:douta	=	16'h	20a2;
51747	:douta	=	16'h	20c2;
51748	:douta	=	16'h	20c2;
51749	:douta	=	16'h	28e2;
51750	:douta	=	16'h	28c2;
51751	:douta	=	16'h	28c2;
51752	:douta	=	16'h	28e2;
51753	:douta	=	16'h	28e2;
51754	:douta	=	16'h	3103;
51755	:douta	=	16'h	3103;
51756	:douta	=	16'h	3103;
51757	:douta	=	16'h	3923;
51758	:douta	=	16'h	41c7;
51759	:douta	=	16'h	424b;
51760	:douta	=	16'h	18e6;
51761	:douta	=	16'h	5163;
51762	:douta	=	16'h	5184;
51763	:douta	=	16'h	5184;
51764	:douta	=	16'h	51a4;
51765	:douta	=	16'h	59c4;
51766	:douta	=	16'h	59c4;
51767	:douta	=	16'h	59c4;
51768	:douta	=	16'h	61e4;
51769	:douta	=	16'h	6204;
51770	:douta	=	16'h	61c3;
51771	:douta	=	16'h	9491;
51772	:douta	=	16'h	b572;
51773	:douta	=	16'h	6a04;
51774	:douta	=	16'h	7245;
51775	:douta	=	16'h	7244;
51776	:douta	=	16'h	7a64;
51777	:douta	=	16'h	7a85;
51778	:douta	=	16'h	7a64;
51779	:douta	=	16'h	7a84;
51780	:douta	=	16'h	8285;
51781	:douta	=	16'h	8aa5;
51782	:douta	=	16'h	51c4;
51783	:douta	=	16'h	82a4;
51784	:douta	=	16'h	7aa5;
51785	:douta	=	16'h	82a4;
51786	:douta	=	16'h	8aa5;
51787	:douta	=	16'h	8ac5;
51788	:douta	=	16'h	8ac5;
51789	:douta	=	16'h	8ae5;
51790	:douta	=	16'h	8ae5;
51791	:douta	=	16'h	92e5;
51792	:douta	=	16'h	8ac5;
51793	:douta	=	16'h	92e5;
51794	:douta	=	16'h	92c4;
51795	:douta	=	16'h	9ae4;
51796	:douta	=	16'h	9ae4;
51797	:douta	=	16'h	9ae4;
51798	:douta	=	16'h	a304;
51799	:douta	=	16'h	a344;
51800	:douta	=	16'h	ab85;
51801	:douta	=	16'h	abc6;
51802	:douta	=	16'h	b408;
51803	:douta	=	16'h	c4ac;
51804	:douta	=	16'h	c4ee;
51805	:douta	=	16'h	cd90;
51806	:douta	=	16'h	d5b1;
51807	:douta	=	16'h	de54;
51808	:douta	=	16'h	e6d7;
51809	:douta	=	16'h	ef18;
51810	:douta	=	16'h	f77a;
51811	:douta	=	16'h	f79a;
51812	:douta	=	16'h	f79a;
51813	:douta	=	16'h	f77a;
51814	:douta	=	16'h	ef58;
51815	:douta	=	16'h	eef6;
51816	:douta	=	16'h	e6b5;
51817	:douta	=	16'h	e633;
51818	:douta	=	16'h	ddcf;
51819	:douta	=	16'h	d56e;
51820	:douta	=	16'h	d50b;
51821	:douta	=	16'h	ccea;
51822	:douta	=	16'h	c467;
51823	:douta	=	16'h	cc46;
51824	:douta	=	16'h	c425;
51825	:douta	=	16'h	c404;
51826	:douta	=	16'h	c404;
51827	:douta	=	16'h	c405;
51828	:douta	=	16'h	cc25;
51829	:douta	=	16'h	cc26;
51830	:douta	=	16'h	cc47;
51831	:douta	=	16'h	cc47;
51832	:douta	=	16'h	cc68;
51833	:douta	=	16'h	cc68;
51834	:douta	=	16'h	cc68;
51835	:douta	=	16'h	cc68;
51836	:douta	=	16'h	cc67;
51837	:douta	=	16'h	cc68;
51838	:douta	=	16'h	cc68;
51839	:douta	=	16'h	cc68;
51840	:douta	=	16'h	cc68;
51841	:douta	=	16'h	cc68;
51842	:douta	=	16'h	cc68;
51843	:douta	=	16'h	d488;
51844	:douta	=	16'h	cc68;
51845	:douta	=	16'h	d488;
51846	:douta	=	16'h	d468;
51847	:douta	=	16'h	cc68;
51848	:douta	=	16'h	d488;
51849	:douta	=	16'h	d488;
51850	:douta	=	16'h	d488;
51851	:douta	=	16'h	d488;
51852	:douta	=	16'h	d488;
51853	:douta	=	16'h	d488;
51854	:douta	=	16'h	d488;
51855	:douta	=	16'h	d488;
51856	:douta	=	16'h	d488;
51857	:douta	=	16'h	cc68;
51858	:douta	=	16'h	cc88;
51859	:douta	=	16'h	cc88;
51860	:douta	=	16'h	d488;
51861	:douta	=	16'h	d488;
51862	:douta	=	16'h	d488;
51863	:douta	=	16'h	cc88;
51864	:douta	=	16'h	d488;
51865	:douta	=	16'h	d488;
51866	:douta	=	16'h	d488;
51867	:douta	=	16'h	d489;
51868	:douta	=	16'h	d4a9;
51869	:douta	=	16'h	d4a9;
51870	:douta	=	16'h	cc88;
51871	:douta	=	16'h	d488;
51872	:douta	=	16'h	d4a9;
51873	:douta	=	16'h	d488;
51874	:douta	=	16'h	cc68;
51875	:douta	=	16'h	cc88;
51876	:douta	=	16'h	d488;
51877	:douta	=	16'h	cc88;
51878	:douta	=	16'h	d4a9;
51879	:douta	=	16'h	d488;
51880	:douta	=	16'h	cc67;
51881	:douta	=	16'h	cc68;
51882	:douta	=	16'h	d4c8;
51883	:douta	=	16'h	d4c9;
51884	:douta	=	16'h	d4c9;
51885	:douta	=	16'h	cc67;
51886	:douta	=	16'h	d468;
51887	:douta	=	16'h	ac6f;
51888	:douta	=	16'h	9c91;
51889	:douta	=	16'h	b513;
51890	:douta	=	16'h	acd2;
51891	:douta	=	16'h	b512;
51892	:douta	=	16'h	bd12;
51893	:douta	=	16'h	b532;
51894	:douta	=	16'h	b513;
51895	:douta	=	16'h	b534;
51896	:douta	=	16'h	acf3;
51897	:douta	=	16'h	9c93;
51898	:douta	=	16'h	8c53;
51899	:douta	=	16'h	8433;
51900	:douta	=	16'h	7bf2;
51901	:douta	=	16'h	73d1;
51902	:douta	=	16'h	7bd1;
51903	:douta	=	16'h	6bb1;
51904	:douta	=	16'h	73b0;
51905	:douta	=	16'h	7bd1;
51906	:douta	=	16'h	62cc;
51907	:douta	=	16'h	2903;
51908	:douta	=	16'h	3965;
51909	:douta	=	16'h	4a27;
51910	:douta	=	16'h	5226;
51911	:douta	=	16'h	41a5;
51912	:douta	=	16'h	5a68;
51913	:douta	=	16'h	3985;
51914	:douta	=	16'h	a490;
51915	:douta	=	16'h	836c;
51916	:douta	=	16'h	836c;
51917	:douta	=	16'h	9c2e;
51918	:douta	=	16'h	7b4b;
51919	:douta	=	16'h	acd1;
51920	:douta	=	16'h	9c4f;
51921	:douta	=	16'h	ac8f;
51922	:douta	=	16'h	a46e;
51923	:douta	=	16'h	a46e;
51924	:douta	=	16'h	a46e;
51925	:douta	=	16'h	acd0;
51926	:douta	=	16'h	942d;
51927	:douta	=	16'h	a490;
51928	:douta	=	16'h	bd11;
51929	:douta	=	16'h	c551;
51930	:douta	=	16'h	cdb3;
51931	:douta	=	16'h	cd93;
51932	:douta	=	16'h	cdb2;
51933	:douta	=	16'h	cdb2;
51934	:douta	=	16'h	d5b3;
51935	:douta	=	16'h	d5d4;
51936	:douta	=	16'h	d5b3;
51937	:douta	=	16'h	c511;
51938	:douta	=	16'h	c571;
51939	:douta	=	16'h	b4d0;
51940	:douta	=	16'h	a450;
51941	:douta	=	16'h	9c30;
51942	:douta	=	16'h	7bae;
51943	:douta	=	16'h	736e;
51944	:douta	=	16'h	4a6b;
51945	:douta	=	16'h	39c9;
51946	:douta	=	16'h	39e9;
51947	:douta	=	16'h	2146;
51948	:douta	=	16'h	2125;
51949	:douta	=	16'h	1906;
51950	:douta	=	16'h	10c4;
51951	:douta	=	16'h	10a4;
51952	:douta	=	16'h	18e4;
51953	:douta	=	16'h	18e4;
51954	:douta	=	16'h	10a3;
51955	:douta	=	16'h	2168;
51956	:douta	=	16'h	1968;
51957	:douta	=	16'h	3945;
51958	:douta	=	16'h	8ae7;
51959	:douta	=	16'h	82a7;
51960	:douta	=	16'h	82a7;
51961	:douta	=	16'h	82c7;
51962	:douta	=	16'h	82a7;
51963	:douta	=	16'h	82c7;
51964	:douta	=	16'h	82a7;
51965	:douta	=	16'h	82a7;
51966	:douta	=	16'h	8ac7;
51967	:douta	=	16'h	82a7;
51968	:douta	=	16'h	ad14;
51969	:douta	=	16'h	ad35;
51970	:douta	=	16'h	cdf6;
51971	:douta	=	16'h	c5b5;
51972	:douta	=	16'h	bd55;
51973	:douta	=	16'h	b555;
51974	:douta	=	16'h	8c53;
51975	:douta	=	16'h	a557;
51976	:douta	=	16'h	94b4;
51977	:douta	=	16'h	9cf5;
51978	:douta	=	16'h	9cd5;
51979	:douta	=	16'h	94d5;
51980	:douta	=	16'h	94b5;
51981	:douta	=	16'h	8c95;
51982	:douta	=	16'h	6b90;
51983	:douta	=	16'h	1060;
51984	:douta	=	16'h	20e3;
51985	:douta	=	16'h	20e3;
51986	:douta	=	16'h	28e3;
51987	:douta	=	16'h	20e3;
51988	:douta	=	16'h	20e3;
51989	:douta	=	16'h	20c3;
51990	:douta	=	16'h	20c3;
51991	:douta	=	16'h	20c3;
51992	:douta	=	16'h	20e3;
51993	:douta	=	16'h	20c3;
51994	:douta	=	16'h	20a2;
51995	:douta	=	16'h	1882;
51996	:douta	=	16'h	20a2;
51997	:douta	=	16'h	20a2;
51998	:douta	=	16'h	20a2;
51999	:douta	=	16'h	20a2;
52000	:douta	=	16'h	20a2;
52001	:douta	=	16'h	20a2;
52002	:douta	=	16'h	20a2;
52003	:douta	=	16'h	20c2;
52004	:douta	=	16'h	28e3;
52005	:douta	=	16'h	28e2;
52006	:douta	=	16'h	28e2;
52007	:douta	=	16'h	28e2;
52008	:douta	=	16'h	28e2;
52009	:douta	=	16'h	3123;
52010	:douta	=	16'h	3123;
52011	:douta	=	16'h	3103;
52012	:douta	=	16'h	3923;
52013	:douta	=	16'h	3923;
52014	:douta	=	16'h	422a;
52015	:douta	=	16'h	424a;
52016	:douta	=	16'h	18c5;
52017	:douta	=	16'h	51a4;
52018	:douta	=	16'h	5184;
52019	:douta	=	16'h	51a4;
52020	:douta	=	16'h	51a4;
52021	:douta	=	16'h	59a4;
52022	:douta	=	16'h	59c4;
52023	:douta	=	16'h	59c4;
52024	:douta	=	16'h	61e3;
52025	:douta	=	16'h	61e4;
52026	:douta	=	16'h	61a3;
52027	:douta	=	16'h	b594;
52028	:douta	=	16'h	acaf;
52029	:douta	=	16'h	7224;
52030	:douta	=	16'h	7264;
52031	:douta	=	16'h	7244;
52032	:douta	=	16'h	7a85;
52033	:douta	=	16'h	7a64;
52034	:douta	=	16'h	7a85;
52035	:douta	=	16'h	7a85;
52036	:douta	=	16'h	7a64;
52037	:douta	=	16'h	8aa4;
52038	:douta	=	16'h	6204;
52039	:douta	=	16'h	8244;
52040	:douta	=	16'h	7a24;
52041	:douta	=	16'h	7a24;
52042	:douta	=	16'h	82a5;
52043	:douta	=	16'h	82c6;
52044	:douta	=	16'h	9327;
52045	:douta	=	16'h	9369;
52046	:douta	=	16'h	a40c;
52047	:douta	=	16'h	b4af;
52048	:douta	=	16'h	bd10;
52049	:douta	=	16'h	c592;
52050	:douta	=	16'h	cdf3;
52051	:douta	=	16'h	de96;
52052	:douta	=	16'h	e6f8;
52053	:douta	=	16'h	e718;
52054	:douta	=	16'h	ef59;
52055	:douta	=	16'h	f779;
52056	:douta	=	16'h	ef37;
52057	:douta	=	16'h	ef17;
52058	:douta	=	16'h	e6b5;
52059	:douta	=	16'h	de32;
52060	:douta	=	16'h	d5f0;
52061	:douta	=	16'h	d54d;
52062	:douta	=	16'h	cd2d;
52063	:douta	=	16'h	c4ca;
52064	:douta	=	16'h	c448;
52065	:douta	=	16'h	bc27;
52066	:douta	=	16'h	bc05;
52067	:douta	=	16'h	bbe5;
52068	:douta	=	16'h	bbc4;
52069	:douta	=	16'h	c3c5;
52070	:douta	=	16'h	bbe5;
52071	:douta	=	16'h	c3e5;
52072	:douta	=	16'h	c405;
52073	:douta	=	16'h	c426;
52074	:douta	=	16'h	c406;
52075	:douta	=	16'h	c427;
52076	:douta	=	16'h	cc47;
52077	:douta	=	16'h	c446;
52078	:douta	=	16'h	cc48;
52079	:douta	=	16'h	cc47;
52080	:douta	=	16'h	cc47;
52081	:douta	=	16'h	cc67;
52082	:douta	=	16'h	cc46;
52083	:douta	=	16'h	cc47;
52084	:douta	=	16'h	cc48;
52085	:douta	=	16'h	cc68;
52086	:douta	=	16'h	cc67;
52087	:douta	=	16'h	cc47;
52088	:douta	=	16'h	cc67;
52089	:douta	=	16'h	cc67;
52090	:douta	=	16'h	cc68;
52091	:douta	=	16'h	cc48;
52092	:douta	=	16'h	cc68;
52093	:douta	=	16'h	cc67;
52094	:douta	=	16'h	cc68;
52095	:douta	=	16'h	cc68;
52096	:douta	=	16'h	cc68;
52097	:douta	=	16'h	cc68;
52098	:douta	=	16'h	cc67;
52099	:douta	=	16'h	cc68;
52100	:douta	=	16'h	cc68;
52101	:douta	=	16'h	cc88;
52102	:douta	=	16'h	cc88;
52103	:douta	=	16'h	cc68;
52104	:douta	=	16'h	cc68;
52105	:douta	=	16'h	cc68;
52106	:douta	=	16'h	d488;
52107	:douta	=	16'h	d488;
52108	:douta	=	16'h	d488;
52109	:douta	=	16'h	d488;
52110	:douta	=	16'h	d488;
52111	:douta	=	16'h	d488;
52112	:douta	=	16'h	d488;
52113	:douta	=	16'h	d487;
52114	:douta	=	16'h	d487;
52115	:douta	=	16'h	d488;
52116	:douta	=	16'h	d488;
52117	:douta	=	16'h	cc88;
52118	:douta	=	16'h	d488;
52119	:douta	=	16'h	cc88;
52120	:douta	=	16'h	d488;
52121	:douta	=	16'h	cc88;
52122	:douta	=	16'h	cc88;
52123	:douta	=	16'h	d488;
52124	:douta	=	16'h	d488;
52125	:douta	=	16'h	d488;
52126	:douta	=	16'h	cc88;
52127	:douta	=	16'h	d488;
52128	:douta	=	16'h	d488;
52129	:douta	=	16'h	d488;
52130	:douta	=	16'h	d4a9;
52131	:douta	=	16'h	cc68;
52132	:douta	=	16'h	d488;
52133	:douta	=	16'h	d489;
52134	:douta	=	16'h	d488;
52135	:douta	=	16'h	d488;
52136	:douta	=	16'h	d487;
52137	:douta	=	16'h	cc46;
52138	:douta	=	16'h	cc25;
52139	:douta	=	16'h	cc25;
52140	:douta	=	16'h	cc45;
52141	:douta	=	16'h	cc67;
52142	:douta	=	16'h	cc87;
52143	:douta	=	16'h	ccec;
52144	:douta	=	16'h	a490;
52145	:douta	=	16'h	acd2;
52146	:douta	=	16'h	a4b2;
52147	:douta	=	16'h	acd2;
52148	:douta	=	16'h	acd3;
52149	:douta	=	16'h	acd3;
52150	:douta	=	16'h	a4b3;
52151	:douta	=	16'h	9cb4;
52152	:douta	=	16'h	9494;
52153	:douta	=	16'h	8412;
52154	:douta	=	16'h	8412;
52155	:douta	=	16'h	7bf2;
52156	:douta	=	16'h	8411;
52157	:douta	=	16'h	738f;
52158	:douta	=	16'h	39a6;
52159	:douta	=	16'h	3944;
52160	:douta	=	16'h	28e3;
52161	:douta	=	16'h	41c4;
52162	:douta	=	16'h	4a05;
52163	:douta	=	16'h	72e9;
52164	:douta	=	16'h	6ae8;
52165	:douta	=	16'h	838b;
52166	:douta	=	16'h	8bcc;
52167	:douta	=	16'h	8bcd;
52168	:douta	=	16'h	734a;
52169	:douta	=	16'h	942e;
52170	:douta	=	16'h	41e6;
52171	:douta	=	16'h	9c6f;
52172	:douta	=	16'h	940d;
52173	:douta	=	16'h	bd51;
52174	:douta	=	16'h	b4f0;
52175	:douta	=	16'h	730b;
52176	:douta	=	16'h	c572;
52177	:douta	=	16'h	acd1;
52178	:douta	=	16'h	bd53;
52179	:douta	=	16'h	bd52;
52180	:douta	=	16'h	cd93;
52181	:douta	=	16'h	bd31;
52182	:douta	=	16'h	bd32;
52183	:douta	=	16'h	d5b3;
52184	:douta	=	16'h	d5b2;
52185	:douta	=	16'h	d5b3;
52186	:douta	=	16'h	d5b3;
52187	:douta	=	16'h	d5b3;
52188	:douta	=	16'h	cd72;
52189	:douta	=	16'h	cd52;
52190	:douta	=	16'h	cd72;
52191	:douta	=	16'h	c532;
52192	:douta	=	16'h	c532;
52193	:douta	=	16'h	b4d1;
52194	:douta	=	16'h	acb1;
52195	:douta	=	16'h	ac91;
52196	:douta	=	16'h	8c10;
52197	:douta	=	16'h	8bf0;
52198	:douta	=	16'h	9c71;
52199	:douta	=	16'h	8c10;
52200	:douta	=	16'h	6b4f;
52201	:douta	=	16'h	5b0d;
52202	:douta	=	16'h	5b0d;
52203	:douta	=	16'h	3a2a;
52204	:douta	=	16'h	39e9;
52205	:douta	=	16'h	2126;
52206	:douta	=	16'h	3a09;
52207	:douta	=	16'h	1906;
52208	:douta	=	16'h	10c4;
52209	:douta	=	16'h	18c4;
52210	:douta	=	16'h	1926;
52211	:douta	=	16'h	1128;
52212	:douta	=	16'h	3a6d;
52213	:douta	=	16'h	936a;
52214	:douta	=	16'h	8aa6;
52215	:douta	=	16'h	8ac7;
52216	:douta	=	16'h	8ac7;
52217	:douta	=	16'h	8ac7;
52218	:douta	=	16'h	8ac7;
52219	:douta	=	16'h	8ac7;
52220	:douta	=	16'h	8ac7;
52221	:douta	=	16'h	8ac7;
52222	:douta	=	16'h	8ac7;
52223	:douta	=	16'h	8ae7;
52224	:douta	=	16'h	ad15;
52225	:douta	=	16'h	b555;
52226	:douta	=	16'h	d616;
52227	:douta	=	16'h	c5b5;
52228	:douta	=	16'h	bd55;
52229	:douta	=	16'h	ad35;
52230	:douta	=	16'h	9494;
52231	:douta	=	16'h	ad57;
52232	:douta	=	16'h	9cd5;
52233	:douta	=	16'h	94d5;
52234	:douta	=	16'h	9cd5;
52235	:douta	=	16'h	94d5;
52236	:douta	=	16'h	8c74;
52237	:douta	=	16'h	8cb5;
52238	:douta	=	16'h	4208;
52239	:douta	=	16'h	1040;
52240	:douta	=	16'h	28e3;
52241	:douta	=	16'h	2103;
52242	:douta	=	16'h	20c3;
52243	:douta	=	16'h	20e3;
52244	:douta	=	16'h	20c3;
52245	:douta	=	16'h	20e3;
52246	:douta	=	16'h	20c3;
52247	:douta	=	16'h	20e3;
52248	:douta	=	16'h	20e3;
52249	:douta	=	16'h	20e3;
52250	:douta	=	16'h	20a3;
52251	:douta	=	16'h	1882;
52252	:douta	=	16'h	20a2;
52253	:douta	=	16'h	20a2;
52254	:douta	=	16'h	20a2;
52255	:douta	=	16'h	1881;
52256	:douta	=	16'h	20a2;
52257	:douta	=	16'h	20a2;
52258	:douta	=	16'h	20a2;
52259	:douta	=	16'h	28e2;
52260	:douta	=	16'h	28e3;
52261	:douta	=	16'h	28c2;
52262	:douta	=	16'h	28e2;
52263	:douta	=	16'h	28e2;
52264	:douta	=	16'h	30e2;
52265	:douta	=	16'h	3103;
52266	:douta	=	16'h	3103;
52267	:douta	=	16'h	3903;
52268	:douta	=	16'h	3923;
52269	:douta	=	16'h	3923;
52270	:douta	=	16'h	4a4b;
52271	:douta	=	16'h	3a09;
52272	:douta	=	16'h	18e5;
52273	:douta	=	16'h	5184;
52274	:douta	=	16'h	5184;
52275	:douta	=	16'h	51a4;
52276	:douta	=	16'h	51a4;
52277	:douta	=	16'h	59c4;
52278	:douta	=	16'h	59c4;
52279	:douta	=	16'h	61e4;
52280	:douta	=	16'h	61e4;
52281	:douta	=	16'h	6a04;
52282	:douta	=	16'h	61c3;
52283	:douta	=	16'h	b594;
52284	:douta	=	16'h	9c2c;
52285	:douta	=	16'h	7224;
52286	:douta	=	16'h	7a44;
52287	:douta	=	16'h	7224;
52288	:douta	=	16'h	7224;
52289	:douta	=	16'h	7203;
52290	:douta	=	16'h	7203;
52291	:douta	=	16'h	7224;
52292	:douta	=	16'h	7224;
52293	:douta	=	16'h	82c6;
52294	:douta	=	16'h	7aa6;
52295	:douta	=	16'h	8b49;
52296	:douta	=	16'h	9beb;
52297	:douta	=	16'h	ac8d;
52298	:douta	=	16'h	bd51;
52299	:douta	=	16'h	bd71;
52300	:douta	=	16'h	cdf3;
52301	:douta	=	16'h	d634;
52302	:douta	=	16'h	deb6;
52303	:douta	=	16'h	ded6;
52304	:douta	=	16'h	ded6;
52305	:douta	=	16'h	e6b5;
52306	:douta	=	16'h	de95;
52307	:douta	=	16'h	de94;
52308	:douta	=	16'h	d631;
52309	:douta	=	16'h	d5f0;
52310	:douta	=	16'h	c54d;
52311	:douta	=	16'h	c50c;
52312	:douta	=	16'h	c4aa;
52313	:douta	=	16'h	bc69;
52314	:douta	=	16'h	b3e7;
52315	:douta	=	16'h	b3c5;
52316	:douta	=	16'h	b3a4;
52317	:douta	=	16'h	b384;
52318	:douta	=	16'h	b3a4;
52319	:douta	=	16'h	bba4;
52320	:douta	=	16'h	bbc4;
52321	:douta	=	16'h	bbc6;
52322	:douta	=	16'h	c3e7;
52323	:douta	=	16'h	c3e7;
52324	:douta	=	16'h	c407;
52325	:douta	=	16'h	c407;
52326	:douta	=	16'h	c406;
52327	:douta	=	16'h	c426;
52328	:douta	=	16'h	c426;
52329	:douta	=	16'h	c427;
52330	:douta	=	16'h	c446;
52331	:douta	=	16'h	c446;
52332	:douta	=	16'h	c447;
52333	:douta	=	16'h	c447;
52334	:douta	=	16'h	c446;
52335	:douta	=	16'h	cc48;
52336	:douta	=	16'h	cc47;
52337	:douta	=	16'h	cc47;
52338	:douta	=	16'h	cc47;
52339	:douta	=	16'h	cc67;
52340	:douta	=	16'h	cc47;
52341	:douta	=	16'h	cc48;
52342	:douta	=	16'h	cc67;
52343	:douta	=	16'h	cc68;
52344	:douta	=	16'h	cc67;
52345	:douta	=	16'h	cc67;
52346	:douta	=	16'h	cc48;
52347	:douta	=	16'h	cc68;
52348	:douta	=	16'h	cc68;
52349	:douta	=	16'h	cc68;
52350	:douta	=	16'h	cc88;
52351	:douta	=	16'h	cc68;
52352	:douta	=	16'h	cc88;
52353	:douta	=	16'h	cc68;
52354	:douta	=	16'h	cc67;
52355	:douta	=	16'h	d488;
52356	:douta	=	16'h	cc68;
52357	:douta	=	16'h	cc68;
52358	:douta	=	16'h	cc68;
52359	:douta	=	16'h	cc68;
52360	:douta	=	16'h	cc67;
52361	:douta	=	16'h	d488;
52362	:douta	=	16'h	d488;
52363	:douta	=	16'h	d488;
52364	:douta	=	16'h	d488;
52365	:douta	=	16'h	d488;
52366	:douta	=	16'h	cc67;
52367	:douta	=	16'h	d488;
52368	:douta	=	16'h	d488;
52369	:douta	=	16'h	cc87;
52370	:douta	=	16'h	d488;
52371	:douta	=	16'h	d488;
52372	:douta	=	16'h	d488;
52373	:douta	=	16'h	d488;
52374	:douta	=	16'h	d488;
52375	:douta	=	16'h	d488;
52376	:douta	=	16'h	d488;
52377	:douta	=	16'h	d488;
52378	:douta	=	16'h	d488;
52379	:douta	=	16'h	d488;
52380	:douta	=	16'h	d488;
52381	:douta	=	16'h	d488;
52382	:douta	=	16'h	d488;
52383	:douta	=	16'h	cc88;
52384	:douta	=	16'h	d487;
52385	:douta	=	16'h	d467;
52386	:douta	=	16'h	d467;
52387	:douta	=	16'h	cc25;
52388	:douta	=	16'h	cc46;
52389	:douta	=	16'h	cc46;
52390	:douta	=	16'h	cca9;
52391	:douta	=	16'h	ccc9;
52392	:douta	=	16'h	cd0b;
52393	:douta	=	16'h	d52c;
52394	:douta	=	16'h	d58f;
52395	:douta	=	16'h	d5d0;
52396	:douta	=	16'h	de53;
52397	:douta	=	16'h	e696;
52398	:douta	=	16'h	eed7;
52399	:douta	=	16'h	ffba;
52400	:douta	=	16'h	e6d7;
52401	:douta	=	16'h	a492;
52402	:douta	=	16'h	a492;
52403	:douta	=	16'h	9cb2;
52404	:douta	=	16'h	a4b3;
52405	:douta	=	16'h	9cb2;
52406	:douta	=	16'h	9472;
52407	:douta	=	16'h	8c53;
52408	:douta	=	16'h	8c93;
52409	:douta	=	16'h	8412;
52410	:douta	=	16'h	7bf2;
52411	:douta	=	16'h	738f;
52412	:douta	=	16'h	4a06;
52413	:douta	=	16'h	3964;
52414	:douta	=	16'h	3124;
52415	:douta	=	16'h	41a5;
52416	:douta	=	16'h	5a68;
52417	:douta	=	16'h	72e9;
52418	:douta	=	16'h	7309;
52419	:douta	=	16'h	7b4a;
52420	:douta	=	16'h	7b2a;
52421	:douta	=	16'h	7b4b;
52422	:douta	=	16'h	940d;
52423	:douta	=	16'h	940d;
52424	:douta	=	16'h	a46e;
52425	:douta	=	16'h	acaf;
52426	:douta	=	16'h	940e;
52427	:douta	=	16'h	6b0a;
52428	:douta	=	16'h	9c2e;
52429	:douta	=	16'h	e654;
52430	:douta	=	16'h	de14;
52431	:douta	=	16'h	5a69;
52432	:douta	=	16'h	c573;
52433	:douta	=	16'h	bd32;
52434	:douta	=	16'h	c594;
52435	:douta	=	16'h	c573;
52436	:douta	=	16'h	bd12;
52437	:douta	=	16'h	bd12;
52438	:douta	=	16'h	bcf2;
52439	:douta	=	16'h	a471;
52440	:douta	=	16'h	b4f2;
52441	:douta	=	16'h	b4f1;
52442	:douta	=	16'h	b4d2;
52443	:douta	=	16'h	b4d2;
52444	:douta	=	16'h	b4d2;
52445	:douta	=	16'h	b4f2;
52446	:douta	=	16'h	acd2;
52447	:douta	=	16'h	acd2;
52448	:douta	=	16'h	acd3;
52449	:douta	=	16'h	9c72;
52450	:douta	=	16'h	9c71;
52451	:douta	=	16'h	a472;
52452	:douta	=	16'h	8c10;
52453	:douta	=	16'h	8c11;
52454	:douta	=	16'h	9451;
52455	:douta	=	16'h	8c11;
52456	:douta	=	16'h	73b0;
52457	:douta	=	16'h	6b6f;
52458	:douta	=	16'h	6b6f;
52459	:douta	=	16'h	4a6c;
52460	:douta	=	16'h	3a4a;
52461	:douta	=	16'h	29a8;
52462	:douta	=	16'h	39e9;
52463	:douta	=	16'h	2188;
52464	:douta	=	16'h	2167;
52465	:douta	=	16'h	18e4;
52466	:douta	=	16'h	1905;
52467	:douta	=	16'h	1106;
52468	:douta	=	16'h	08e6;
52469	:douta	=	16'h	8309;
52470	:douta	=	16'h	82a8;
52471	:douta	=	16'h	8ac7;
52472	:douta	=	16'h	8ae7;
52473	:douta	=	16'h	8ac7;
52474	:douta	=	16'h	8b08;
52475	:douta	=	16'h	8ae7;
52476	:douta	=	16'h	8ac7;
52477	:douta	=	16'h	8ae7;
52478	:douta	=	16'h	8ae7;
52479	:douta	=	16'h	8ae7;
52480	:douta	=	16'h	ad56;
52481	:douta	=	16'h	cdb5;
52482	:douta	=	16'h	cdf6;
52483	:douta	=	16'h	c596;
52484	:douta	=	16'h	b555;
52485	:douta	=	16'h	9494;
52486	:douta	=	16'h	a516;
52487	:douta	=	16'h	ad57;
52488	:douta	=	16'h	a4f5;
52489	:douta	=	16'h	9cf6;
52490	:douta	=	16'h	9cd5;
52491	:douta	=	16'h	8c75;
52492	:douta	=	16'h	8454;
52493	:douta	=	16'h	a558;
52494	:douta	=	16'h	2965;
52495	:douta	=	16'h	3165;
52496	:douta	=	16'h	2082;
52497	:douta	=	16'h	1882;
52498	:douta	=	16'h	20c3;
52499	:douta	=	16'h	20e3;
52500	:douta	=	16'h	20c3;
52501	:douta	=	16'h	20e3;
52502	:douta	=	16'h	20c3;
52503	:douta	=	16'h	20e3;
52504	:douta	=	16'h	20c3;
52505	:douta	=	16'h	20c3;
52506	:douta	=	16'h	1882;
52507	:douta	=	16'h	18a2;
52508	:douta	=	16'h	20a2;
52509	:douta	=	16'h	20a2;
52510	:douta	=	16'h	20a2;
52511	:douta	=	16'h	20c2;
52512	:douta	=	16'h	20a2;
52513	:douta	=	16'h	20a2;
52514	:douta	=	16'h	20a2;
52515	:douta	=	16'h	20a2;
52516	:douta	=	16'h	28e2;
52517	:douta	=	16'h	28e2;
52518	:douta	=	16'h	28e2;
52519	:douta	=	16'h	28e2;
52520	:douta	=	16'h	30e2;
52521	:douta	=	16'h	3103;
52522	:douta	=	16'h	3123;
52523	:douta	=	16'h	3923;
52524	:douta	=	16'h	3923;
52525	:douta	=	16'h	3923;
52526	:douta	=	16'h	4a4b;
52527	:douta	=	16'h	31a8;
52528	:douta	=	16'h	2904;
52529	:douta	=	16'h	5184;
52530	:douta	=	16'h	5184;
52531	:douta	=	16'h	5163;
52532	:douta	=	16'h	5163;
52533	:douta	=	16'h	5163;
52534	:douta	=	16'h	5983;
52535	:douta	=	16'h	5984;
52536	:douta	=	16'h	61a4;
52537	:douta	=	16'h	61e4;
52538	:douta	=	16'h	7266;
52539	:douta	=	16'h	ad51;
52540	:douta	=	16'h	9c0d;
52541	:douta	=	16'h	9c4c;
52542	:douta	=	16'h	a48d;
52543	:douta	=	16'h	b4f1;
52544	:douta	=	16'h	c5b2;
52545	:douta	=	16'h	ce13;
52546	:douta	=	16'h	d654;
52547	:douta	=	16'h	d674;
52548	:douta	=	16'h	d674;
52549	:douta	=	16'h	d654;
52550	:douta	=	16'h	deb5;
52551	:douta	=	16'h	8ba9;
52552	:douta	=	16'h	cdf2;
52553	:douta	=	16'h	b4cd;
52554	:douta	=	16'h	a44b;
52555	:douta	=	16'h	a42b;
52556	:douta	=	16'h	9ba9;
52557	:douta	=	16'h	9b88;
52558	:douta	=	16'h	9326;
52559	:douta	=	16'h	8ae5;
52560	:douta	=	16'h	8ac5;
52561	:douta	=	16'h	92c5;
52562	:douta	=	16'h	9b05;
52563	:douta	=	16'h	9b05;
52564	:douta	=	16'h	a346;
52565	:douta	=	16'h	ab46;
52566	:douta	=	16'h	ab86;
52567	:douta	=	16'h	ab87;
52568	:douta	=	16'h	b3a7;
52569	:douta	=	16'h	b3c7;
52570	:douta	=	16'h	b3c7;
52571	:douta	=	16'h	bbc7;
52572	:douta	=	16'h	bbc7;
52573	:douta	=	16'h	bbc6;
52574	:douta	=	16'h	bbe6;
52575	:douta	=	16'h	bbe7;
52576	:douta	=	16'h	c406;
52577	:douta	=	16'h	c406;
52578	:douta	=	16'h	c406;
52579	:douta	=	16'h	c406;
52580	:douta	=	16'h	c406;
52581	:douta	=	16'h	c427;
52582	:douta	=	16'h	c426;
52583	:douta	=	16'h	c447;
52584	:douta	=	16'h	c426;
52585	:douta	=	16'h	c427;
52586	:douta	=	16'h	c427;
52587	:douta	=	16'h	c427;
52588	:douta	=	16'h	c428;
52589	:douta	=	16'h	cc47;
52590	:douta	=	16'h	cc27;
52591	:douta	=	16'h	cc47;
52592	:douta	=	16'h	cc47;
52593	:douta	=	16'h	cc67;
52594	:douta	=	16'h	cc67;
52595	:douta	=	16'h	cc67;
52596	:douta	=	16'h	cc67;
52597	:douta	=	16'h	cc67;
52598	:douta	=	16'h	cc67;
52599	:douta	=	16'h	cc68;
52600	:douta	=	16'h	cc68;
52601	:douta	=	16'h	cc67;
52602	:douta	=	16'h	cc67;
52603	:douta	=	16'h	cc67;
52604	:douta	=	16'h	cc67;
52605	:douta	=	16'h	cc68;
52606	:douta	=	16'h	cc68;
52607	:douta	=	16'h	cc68;
52608	:douta	=	16'h	cc68;
52609	:douta	=	16'h	cc88;
52610	:douta	=	16'h	cc67;
52611	:douta	=	16'h	cc68;
52612	:douta	=	16'h	cc68;
52613	:douta	=	16'h	d488;
52614	:douta	=	16'h	cc67;
52615	:douta	=	16'h	cc68;
52616	:douta	=	16'h	d488;
52617	:douta	=	16'h	d488;
52618	:douta	=	16'h	cc68;
52619	:douta	=	16'h	cc88;
52620	:douta	=	16'h	cc88;
52621	:douta	=	16'h	d488;
52622	:douta	=	16'h	cc68;
52623	:douta	=	16'h	d488;
52624	:douta	=	16'h	cc67;
52625	:douta	=	16'h	d487;
52626	:douta	=	16'h	cc66;
52627	:douta	=	16'h	cc46;
52628	:douta	=	16'h	cc45;
52629	:douta	=	16'h	cc25;
52630	:douta	=	16'h	cc25;
52631	:douta	=	16'h	cc26;
52632	:douta	=	16'h	cc47;
52633	:douta	=	16'h	cc89;
52634	:douta	=	16'h	d4aa;
52635	:douta	=	16'h	d50d;
52636	:douta	=	16'h	d56f;
52637	:douta	=	16'h	ddb1;
52638	:douta	=	16'h	de14;
52639	:douta	=	16'h	e655;
52640	:douta	=	16'h	eed7;
52641	:douta	=	16'h	ef19;
52642	:douta	=	16'h	f75b;
52643	:douta	=	16'h	f79c;
52644	:douta	=	16'h	f79c;
52645	:douta	=	16'h	fffe;
52646	:douta	=	16'h	f77a;
52647	:douta	=	16'h	f758;
52648	:douta	=	16'h	eed6;
52649	:douta	=	16'h	ee94;
52650	:douta	=	16'h	de11;
52651	:douta	=	16'h	e5d0;
52652	:douta	=	16'h	dd6d;
52653	:douta	=	16'h	d50a;
52654	:douta	=	16'h	d4e9;
52655	:douta	=	16'h	d486;
52656	:douta	=	16'h	c469;
52657	:douta	=	16'h	a4b2;
52658	:douta	=	16'h	a4b3;
52659	:douta	=	16'h	a492;
52660	:douta	=	16'h	9452;
52661	:douta	=	16'h	9432;
52662	:douta	=	16'h	83f1;
52663	:douta	=	16'h	83f0;
52664	:douta	=	16'h	6b2c;
52665	:douta	=	16'h	49c6;
52666	:douta	=	16'h	51e6;
52667	:douta	=	16'h	49e6;
52668	:douta	=	16'h	6aca;
52669	:douta	=	16'h	62a9;
52670	:douta	=	16'h	836b;
52671	:douta	=	16'h	7b2b;
52672	:douta	=	16'h	8bcd;
52673	:douta	=	16'h	838b;
52674	:douta	=	16'h	8bac;
52675	:douta	=	16'h	a42e;
52676	:douta	=	16'h	9c2e;
52677	:douta	=	16'h	ac8f;
52678	:douta	=	16'h	a46e;
52679	:douta	=	16'h	8bed;
52680	:douta	=	16'h	cd92;
52681	:douta	=	16'h	d593;
52682	:douta	=	16'h	d5d3;
52683	:douta	=	16'h	acd1;
52684	:douta	=	16'h	a490;
52685	:douta	=	16'h	736d;
52686	:douta	=	16'h	9451;
52687	:douta	=	16'h	e615;
52688	:douta	=	16'h	9430;
52689	:douta	=	16'h	c573;
52690	:douta	=	16'h	acd2;
52691	:douta	=	16'h	b513;
52692	:douta	=	16'h	a493;
52693	:douta	=	16'h	9472;
52694	:douta	=	16'h	8412;
52695	:douta	=	16'h	7bf1;
52696	:douta	=	16'h	6b4f;
52697	:douta	=	16'h	7bd1;
52698	:douta	=	16'h	8453;
52699	:douta	=	16'h	8c74;
52700	:douta	=	16'h	8c54;
52701	:douta	=	16'h	8c74;
52702	:douta	=	16'h	9494;
52703	:douta	=	16'h	8c74;
52704	:douta	=	16'h	8c74;
52705	:douta	=	16'h	9473;
52706	:douta	=	16'h	8c53;
52707	:douta	=	16'h	9473;
52708	:douta	=	16'h	8c32;
52709	:douta	=	16'h	8412;
52710	:douta	=	16'h	8c32;
52711	:douta	=	16'h	9453;
52712	:douta	=	16'h	8452;
52713	:douta	=	16'h	73d2;
52714	:douta	=	16'h	7c53;
52715	:douta	=	16'h	73f2;
52716	:douta	=	16'h	6370;
52717	:douta	=	16'h	428e;
52718	:douta	=	16'h	3a2b;
52719	:douta	=	16'h	320a;
52720	:douta	=	16'h	2147;
52721	:douta	=	16'h	2946;
52722	:douta	=	16'h	2126;
52723	:douta	=	16'h	1907;
52724	:douta	=	16'h	2169;
52725	:douta	=	16'h	5acb;
52726	:douta	=	16'h	7245;
52727	:douta	=	16'h	92e8;
52728	:douta	=	16'h	92e8;
52729	:douta	=	16'h	92e8;
52730	:douta	=	16'h	8ae7;
52731	:douta	=	16'h	8ae7;
52732	:douta	=	16'h	8ae7;
52733	:douta	=	16'h	8ae8;
52734	:douta	=	16'h	8ae7;
52735	:douta	=	16'h	9307;
52736	:douta	=	16'h	ad36;
52737	:douta	=	16'h	d5f6;
52738	:douta	=	16'h	cdf6;
52739	:douta	=	16'h	c5b5;
52740	:douta	=	16'h	ad15;
52741	:douta	=	16'h	9453;
52742	:douta	=	16'h	ad77;
52743	:douta	=	16'h	a516;
52744	:douta	=	16'h	9cf5;
52745	:douta	=	16'h	9cd6;
52746	:douta	=	16'h	9cd5;
52747	:douta	=	16'h	8c74;
52748	:douta	=	16'h	8454;
52749	:douta	=	16'h	8474;
52750	:douta	=	16'h	3a2a;
52751	:douta	=	16'h	4aac;
52752	:douta	=	16'h	39c8;
52753	:douta	=	16'h	3146;
52754	:douta	=	16'h	20a2;
52755	:douta	=	16'h	20c2;
52756	:douta	=	16'h	20c3;
52757	:douta	=	16'h	20e3;
52758	:douta	=	16'h	20c3;
52759	:douta	=	16'h	28e3;
52760	:douta	=	16'h	20e3;
52761	:douta	=	16'h	20e3;
52762	:douta	=	16'h	1882;
52763	:douta	=	16'h	18a2;
52764	:douta	=	16'h	20a2;
52765	:douta	=	16'h	18a2;
52766	:douta	=	16'h	18a2;
52767	:douta	=	16'h	20c2;
52768	:douta	=	16'h	20a2;
52769	:douta	=	16'h	20a2;
52770	:douta	=	16'h	20c2;
52771	:douta	=	16'h	20c2;
52772	:douta	=	16'h	28e3;
52773	:douta	=	16'h	28e3;
52774	:douta	=	16'h	28e2;
52775	:douta	=	16'h	30e2;
52776	:douta	=	16'h	30e2;
52777	:douta	=	16'h	3903;
52778	:douta	=	16'h	3103;
52779	:douta	=	16'h	3103;
52780	:douta	=	16'h	30e2;
52781	:douta	=	16'h	38e2;
52782	:douta	=	16'h	422a;
52783	:douta	=	16'h	2947;
52784	:douta	=	16'h	28e4;
52785	:douta	=	16'h	4943;
52786	:douta	=	16'h	5184;
52787	:douta	=	16'h	51c4;
52788	:douta	=	16'h	5a05;
52789	:douta	=	16'h	6a87;
52790	:douta	=	16'h	7308;
52791	:douta	=	16'h	836a;
52792	:douta	=	16'h	93ec;
52793	:douta	=	16'h	9c6e;
52794	:douta	=	16'h	b530;
52795	:douta	=	16'h	bd91;
52796	:douta	=	16'h	c5f3;
52797	:douta	=	16'h	ce34;
52798	:douta	=	16'h	ce33;
52799	:douta	=	16'h	cdf2;
52800	:douta	=	16'h	c591;
52801	:douta	=	16'h	bd70;
52802	:douta	=	16'h	acee;
52803	:douta	=	16'h	ac8d;
52804	:douta	=	16'h	a40b;
52805	:douta	=	16'h	93ca;
52806	:douta	=	16'h	9bea;
52807	:douta	=	16'h	49c4;
52808	:douta	=	16'h	9327;
52809	:douta	=	16'h	8285;
52810	:douta	=	16'h	8284;
52811	:douta	=	16'h	8283;
52812	:douta	=	16'h	8284;
52813	:douta	=	16'h	8aa4;
52814	:douta	=	16'h	8aa4;
52815	:douta	=	16'h	92c6;
52816	:douta	=	16'h	9306;
52817	:douta	=	16'h	9306;
52818	:douta	=	16'h	9b26;
52819	:douta	=	16'h	a366;
52820	:douta	=	16'h	a386;
52821	:douta	=	16'h	ab67;
52822	:douta	=	16'h	ab86;
52823	:douta	=	16'h	b3a6;
52824	:douta	=	16'h	b3a6;
52825	:douta	=	16'h	b3c7;
52826	:douta	=	16'h	b3c6;
52827	:douta	=	16'h	bbc6;
52828	:douta	=	16'h	bbe6;
52829	:douta	=	16'h	bbe6;
52830	:douta	=	16'h	bbe6;
52831	:douta	=	16'h	bbe6;
52832	:douta	=	16'h	bc06;
52833	:douta	=	16'h	bbe6;
52834	:douta	=	16'h	c427;
52835	:douta	=	16'h	c427;
52836	:douta	=	16'h	c407;
52837	:douta	=	16'h	c407;
52838	:douta	=	16'h	c427;
52839	:douta	=	16'h	cc47;
52840	:douta	=	16'h	c427;
52841	:douta	=	16'h	c446;
52842	:douta	=	16'h	c426;
52843	:douta	=	16'h	c427;
52844	:douta	=	16'h	cc47;
52845	:douta	=	16'h	c446;
52846	:douta	=	16'h	cc47;
52847	:douta	=	16'h	cc47;
52848	:douta	=	16'h	cc47;
52849	:douta	=	16'h	cc47;
52850	:douta	=	16'h	c447;
52851	:douta	=	16'h	cc47;
52852	:douta	=	16'h	cc48;
52853	:douta	=	16'h	cc47;
52854	:douta	=	16'h	cc67;
52855	:douta	=	16'h	cc68;
52856	:douta	=	16'h	cc47;
52857	:douta	=	16'h	cc68;
52858	:douta	=	16'h	cc68;
52859	:douta	=	16'h	cc68;
52860	:douta	=	16'h	cc69;
52861	:douta	=	16'h	cc68;
52862	:douta	=	16'h	cc88;
52863	:douta	=	16'h	cc88;
52864	:douta	=	16'h	cc67;
52865	:douta	=	16'h	cc68;
52866	:douta	=	16'h	cc68;
52867	:douta	=	16'h	d488;
52868	:douta	=	16'h	d488;
52869	:douta	=	16'h	cc67;
52870	:douta	=	16'h	cc67;
52871	:douta	=	16'h	cc68;
52872	:douta	=	16'h	cc87;
52873	:douta	=	16'h	cc87;
52874	:douta	=	16'h	d467;
52875	:douta	=	16'h	cc66;
52876	:douta	=	16'h	d446;
52877	:douta	=	16'h	d446;
52878	:douta	=	16'h	cc45;
52879	:douta	=	16'h	cc25;
52880	:douta	=	16'h	cc45;
52881	:douta	=	16'h	cc66;
52882	:douta	=	16'h	cca9;
52883	:douta	=	16'h	cccb;
52884	:douta	=	16'h	d52d;
52885	:douta	=	16'h	d54e;
52886	:douta	=	16'h	ddb1;
52887	:douta	=	16'h	de33;
52888	:douta	=	16'h	e675;
52889	:douta	=	16'h	e6d7;
52890	:douta	=	16'h	ef18;
52891	:douta	=	16'h	f77b;
52892	:douta	=	16'h	f7bc;
52893	:douta	=	16'h	ffdd;
52894	:douta	=	16'h	fffc;
52895	:douta	=	16'h	ffdc;
52896	:douta	=	16'h	ff9a;
52897	:douta	=	16'h	f759;
52898	:douta	=	16'h	ef17;
52899	:douta	=	16'h	f6d6;
52900	:douta	=	16'h	f75a;
52901	:douta	=	16'h	ee10;
52902	:douta	=	16'h	d50b;
52903	:douta	=	16'h	d50a;
52904	:douta	=	16'h	d4c9;
52905	:douta	=	16'h	cca8;
52906	:douta	=	16'h	cc67;
52907	:douta	=	16'h	cc46;
52908	:douta	=	16'h	cc47;
52909	:douta	=	16'h	cc67;
52910	:douta	=	16'h	d468;
52911	:douta	=	16'h	d447;
52912	:douta	=	16'h	cc68;
52913	:douta	=	16'h	9c93;
52914	:douta	=	16'h	a492;
52915	:douta	=	16'h	9472;
52916	:douta	=	16'h	8411;
52917	:douta	=	16'h	8411;
52918	:douta	=	16'h	734e;
52919	:douta	=	16'h	5226;
52920	:douta	=	16'h	3163;
52921	:douta	=	16'h	5227;
52922	:douta	=	16'h	5a68;
52923	:douta	=	16'h	732b;
52924	:douta	=	16'h	7b4b;
52925	:douta	=	16'h	734b;
52926	:douta	=	16'h	7b4b;
52927	:douta	=	16'h	836b;
52928	:douta	=	16'h	9c4e;
52929	:douta	=	16'h	9c0d;
52930	:douta	=	16'h	a44e;
52931	:douta	=	16'h	a46e;
52932	:douta	=	16'h	ac8f;
52933	:douta	=	16'h	b4f0;
52934	:douta	=	16'h	c531;
52935	:douta	=	16'h	940e;
52936	:douta	=	16'h	d5b3;
52937	:douta	=	16'h	d615;
52938	:douta	=	16'h	c552;
52939	:douta	=	16'h	de16;
52940	:douta	=	16'h	d5b3;
52941	:douta	=	16'h	838e;
52942	:douta	=	16'h	6b6f;
52943	:douta	=	16'h	a491;
52944	:douta	=	16'h	8390;
52945	:douta	=	16'h	acd2;
52946	:douta	=	16'h	a4b3;
52947	:douta	=	16'h	a473;
52948	:douta	=	16'h	9c72;
52949	:douta	=	16'h	8c32;
52950	:douta	=	16'h	8412;
52951	:douta	=	16'h	73b0;
52952	:douta	=	16'h	6b4f;
52953	:douta	=	16'h	7390;
52954	:douta	=	16'h	7bd1;
52955	:douta	=	16'h	7bf1;
52956	:douta	=	16'h	8453;
52957	:douta	=	16'h	8432;
52958	:douta	=	16'h	8453;
52959	:douta	=	16'h	8c94;
52960	:douta	=	16'h	8c75;
52961	:douta	=	16'h	8453;
52962	:douta	=	16'h	9474;
52963	:douta	=	16'h	8c53;
52964	:douta	=	16'h	8c73;
52965	:douta	=	16'h	8c32;
52966	:douta	=	16'h	83f1;
52967	:douta	=	16'h	8c52;
52968	:douta	=	16'h	8c74;
52969	:douta	=	16'h	6bd2;
52970	:douta	=	16'h	7c13;
52971	:douta	=	16'h	7c54;
52972	:douta	=	16'h	73f3;
52973	:douta	=	16'h	530f;
52974	:douta	=	16'h	320a;
52975	:douta	=	16'h	3a2b;
52976	:douta	=	16'h	2947;
52977	:douta	=	16'h	2146;
52978	:douta	=	16'h	2125;
52979	:douta	=	16'h	428b;
52980	:douta	=	16'h	b5b6;
52981	:douta	=	16'h	8c10;
52982	:douta	=	16'h	61c4;
52983	:douta	=	16'h	9309;
52984	:douta	=	16'h	92e8;
52985	:douta	=	16'h	8b07;
52986	:douta	=	16'h	9307;
52987	:douta	=	16'h	9307;
52988	:douta	=	16'h	9307;
52989	:douta	=	16'h	9308;
52990	:douta	=	16'h	9308;
52991	:douta	=	16'h	9308;
52992	:douta	=	16'h	ad36;
52993	:douta	=	16'h	cdd6;
52994	:douta	=	16'h	c5b5;
52995	:douta	=	16'h	bd95;
52996	:douta	=	16'h	9c94;
52997	:douta	=	16'h	9453;
52998	:douta	=	16'h	ad57;
52999	:douta	=	16'h	9cf5;
53000	:douta	=	16'h	9cd5;
53001	:douta	=	16'h	94d5;
53002	:douta	=	16'h	9cd5;
53003	:douta	=	16'h	8433;
53004	:douta	=	16'h	94d7;
53005	:douta	=	16'h	2103;
53006	:douta	=	16'h	20c3;
53007	:douta	=	16'h	20c3;
53008	:douta	=	16'h	2904;
53009	:douta	=	16'h	3987;
53010	:douta	=	16'h	426b;
53011	:douta	=	16'h	426b;
53012	:douta	=	16'h	3a29;
53013	:douta	=	16'h	2104;
53014	:douta	=	16'h	20c2;
53015	:douta	=	16'h	20a2;
53016	:douta	=	16'h	20e3;
53017	:douta	=	16'h	20e3;
53018	:douta	=	16'h	2082;
53019	:douta	=	16'h	20a2;
53020	:douta	=	16'h	1881;
53021	:douta	=	16'h	2082;
53022	:douta	=	16'h	1881;
53023	:douta	=	16'h	1861;
53024	:douta	=	16'h	1881;
53025	:douta	=	16'h	2081;
53026	:douta	=	16'h	2082;
53027	:douta	=	16'h	2082;
53028	:douta	=	16'h	28e3;
53029	:douta	=	16'h	28e3;
53030	:douta	=	16'h	3144;
53031	:douta	=	16'h	3965;
53032	:douta	=	16'h	41a5;
53033	:douta	=	16'h	5227;
53034	:douta	=	16'h	5248;
53035	:douta	=	16'h	62c9;
53036	:douta	=	16'h	736c;
53037	:douta	=	16'h	7b6c;
53038	:douta	=	16'h	39c8;
53039	:douta	=	16'h	1906;
53040	:douta	=	16'h	7b6c;
53041	:douta	=	16'h	9c90;
53042	:douta	=	16'h	948f;
53043	:douta	=	16'h	944e;
53044	:douta	=	16'h	942e;
53045	:douta	=	16'h	8bcb;
53046	:douta	=	16'h	834a;
53047	:douta	=	16'h	7b29;
53048	:douta	=	16'h	72c7;
53049	:douta	=	16'h	72a6;
53050	:douta	=	16'h	6a45;
53051	:douta	=	16'h	7224;
53052	:douta	=	16'h	7224;
53053	:douta	=	16'h	7224;
53054	:douta	=	16'h	7204;
53055	:douta	=	16'h	7203;
53056	:douta	=	16'h	7244;
53057	:douta	=	16'h	7a44;
53058	:douta	=	16'h	7a65;
53059	:douta	=	16'h	8285;
53060	:douta	=	16'h	82a5;
53061	:douta	=	16'h	82a6;
53062	:douta	=	16'h	82c5;
53063	:douta	=	16'h	51a4;
53064	:douta	=	16'h	7a65;
53065	:douta	=	16'h	8ac6;
53066	:douta	=	16'h	8ae5;
53067	:douta	=	16'h	92e5;
53068	:douta	=	16'h	92c6;
53069	:douta	=	16'h	92e5;
53070	:douta	=	16'h	9306;
53071	:douta	=	16'h	9306;
53072	:douta	=	16'h	9306;
53073	:douta	=	16'h	9306;
53074	:douta	=	16'h	9b46;
53075	:douta	=	16'h	a366;
53076	:douta	=	16'h	ab87;
53077	:douta	=	16'h	ab86;
53078	:douta	=	16'h	ab86;
53079	:douta	=	16'h	b3a6;
53080	:douta	=	16'h	b3a7;
53081	:douta	=	16'h	b3c7;
53082	:douta	=	16'h	b3c7;
53083	:douta	=	16'h	bbe7;
53084	:douta	=	16'h	bbe7;
53085	:douta	=	16'h	bbc6;
53086	:douta	=	16'h	bbe7;
53087	:douta	=	16'h	bbe6;
53088	:douta	=	16'h	c407;
53089	:douta	=	16'h	c407;
53090	:douta	=	16'h	bc07;
53091	:douta	=	16'h	c407;
53092	:douta	=	16'h	c407;
53093	:douta	=	16'h	c406;
53094	:douta	=	16'h	c426;
53095	:douta	=	16'h	c426;
53096	:douta	=	16'h	c427;
53097	:douta	=	16'h	c447;
53098	:douta	=	16'h	c427;
53099	:douta	=	16'h	cc47;
53100	:douta	=	16'h	cc27;
53101	:douta	=	16'h	c446;
53102	:douta	=	16'h	cc47;
53103	:douta	=	16'h	cc47;
53104	:douta	=	16'h	cc47;
53105	:douta	=	16'h	cc47;
53106	:douta	=	16'h	cc48;
53107	:douta	=	16'h	cc67;
53108	:douta	=	16'h	cc67;
53109	:douta	=	16'h	cc68;
53110	:douta	=	16'h	cc47;
53111	:douta	=	16'h	cc48;
53112	:douta	=	16'h	cc68;
53113	:douta	=	16'h	cc67;
53114	:douta	=	16'h	cc67;
53115	:douta	=	16'h	cc67;
53116	:douta	=	16'h	cc67;
53117	:douta	=	16'h	cc25;
53118	:douta	=	16'h	cc25;
53119	:douta	=	16'h	cc25;
53120	:douta	=	16'h	cc25;
53121	:douta	=	16'h	c404;
53122	:douta	=	16'h	cc46;
53123	:douta	=	16'h	cc68;
53124	:douta	=	16'h	cca9;
53125	:douta	=	16'h	d50b;
53126	:douta	=	16'h	d52c;
53127	:douta	=	16'h	dd8f;
53128	:douta	=	16'h	de13;
53129	:douta	=	16'h	de34;
53130	:douta	=	16'h	e6b7;
53131	:douta	=	16'h	eef8;
53132	:douta	=	16'h	f75a;
53133	:douta	=	16'h	f79c;
53134	:douta	=	16'h	f7bd;
53135	:douta	=	16'h	ffdc;
53136	:douta	=	16'h	ffdc;
53137	:douta	=	16'h	ffdb;
53138	:douta	=	16'h	f77a;
53139	:douta	=	16'h	f738;
53140	:douta	=	16'h	eed6;
53141	:douta	=	16'h	eeb5;
53142	:douta	=	16'h	e653;
53143	:douta	=	16'h	ddcf;
53144	:douta	=	16'h	dd8f;
53145	:douta	=	16'h	d54d;
53146	:douta	=	16'h	d50b;
53147	:douta	=	16'h	cca9;
53148	:douta	=	16'h	cc67;
53149	:douta	=	16'h	cc66;
53150	:douta	=	16'h	cc46;
53151	:douta	=	16'h	cc26;
53152	:douta	=	16'h	cc66;
53153	:douta	=	16'h	cc46;
53154	:douta	=	16'h	d425;
53155	:douta	=	16'h	ad11;
53156	:douta	=	16'h	de97;
53157	:douta	=	16'h	cc26;
53158	:douta	=	16'h	d489;
53159	:douta	=	16'h	d4a9;
53160	:douta	=	16'h	d488;
53161	:douta	=	16'h	d488;
53162	:douta	=	16'h	cc88;
53163	:douta	=	16'h	cc88;
53164	:douta	=	16'h	d489;
53165	:douta	=	16'h	cc89;
53166	:douta	=	16'h	cc69;
53167	:douta	=	16'h	cc68;
53168	:douta	=	16'h	dc87;
53169	:douta	=	16'h	9493;
53170	:douta	=	16'h	83ae;
53171	:douta	=	16'h	62aa;
53172	:douta	=	16'h	4185;
53173	:douta	=	16'h	3985;
53174	:douta	=	16'h	62a8;
53175	:douta	=	16'h	730a;
53176	:douta	=	16'h	7b4b;
53177	:douta	=	16'h	7b4b;
53178	:douta	=	16'h	7b6b;
53179	:douta	=	16'h	8c0e;
53180	:douta	=	16'h	8c0d;
53181	:douta	=	16'h	940d;
53182	:douta	=	16'h	a48f;
53183	:douta	=	16'h	acaf;
53184	:douta	=	16'h	b4f0;
53185	:douta	=	16'h	bd11;
53186	:douta	=	16'h	bd10;
53187	:douta	=	16'h	cd73;
53188	:douta	=	16'h	cdb4;
53189	:douta	=	16'h	c572;
53190	:douta	=	16'h	acb0;
53191	:douta	=	16'h	8bad;
53192	:douta	=	16'h	ddd4;
53193	:douta	=	16'h	d5b3;
53194	:douta	=	16'h	cd93;
53195	:douta	=	16'h	acb3;
53196	:douta	=	16'h	9c52;
53197	:douta	=	16'h	9473;
53198	:douta	=	16'h	8412;
53199	:douta	=	16'h	7390;
53200	:douta	=	16'h	a4b2;
53201	:douta	=	16'h	acb3;
53202	:douta	=	16'h	9452;
53203	:douta	=	16'h	8c32;
53204	:douta	=	16'h	83f1;
53205	:douta	=	16'h	83f1;
53206	:douta	=	16'h	7bb1;
53207	:douta	=	16'h	7390;
53208	:douta	=	16'h	6b4f;
53209	:douta	=	16'h	630e;
53210	:douta	=	16'h	736f;
53211	:douta	=	16'h	738f;
53212	:douta	=	16'h	7390;
53213	:douta	=	16'h	73b0;
53214	:douta	=	16'h	7390;
53215	:douta	=	16'h	6b4f;
53216	:douta	=	16'h	736f;
53217	:douta	=	16'h	7390;
53218	:douta	=	16'h	6b6f;
53219	:douta	=	16'h	73b1;
53220	:douta	=	16'h	73b0;
53221	:douta	=	16'h	73d1;
53222	:douta	=	16'h	73b1;
53223	:douta	=	16'h	6b70;
53224	:douta	=	16'h	7c12;
53225	:douta	=	16'h	7bf3;
53226	:douta	=	16'h	7433;
53227	:douta	=	16'h	6370;
53228	:douta	=	16'h	6391;
53229	:douta	=	16'h	7c75;
53230	:douta	=	16'h	6350;
53231	:douta	=	16'h	3a2a;
53232	:douta	=	16'h	2147;
53233	:douta	=	16'h	29c9;
53234	:douta	=	16'h	2a4c;
53235	:douta	=	16'h	ffff;
53236	:douta	=	16'h	ffff;
53237	:douta	=	16'h	ffff;
53238	:douta	=	16'h	938e;
53239	:douta	=	16'h	9b49;
53240	:douta	=	16'h	9328;
53241	:douta	=	16'h	9308;
53242	:douta	=	16'h	9307;
53243	:douta	=	16'h	9328;
53244	:douta	=	16'h	9307;
53245	:douta	=	16'h	9307;
53246	:douta	=	16'h	9b28;
53247	:douta	=	16'h	9328;
53248	:douta	=	16'h	b556;
53249	:douta	=	16'h	cdd6;
53250	:douta	=	16'h	cdb5;
53251	:douta	=	16'h	bd75;
53252	:douta	=	16'h	8c53;
53253	:douta	=	16'h	9cb5;
53254	:douta	=	16'h	a516;
53255	:douta	=	16'h	a4f5;
53256	:douta	=	16'h	9cd5;
53257	:douta	=	16'h	9cf6;
53258	:douta	=	16'h	9cb5;
53259	:douta	=	16'h	8c74;
53260	:douta	=	16'h	9d79;
53261	:douta	=	16'h	1020;
53262	:douta	=	16'h	28e3;
53263	:douta	=	16'h	28e3;
53264	:douta	=	16'h	20a2;
53265	:douta	=	16'h	20c2;
53266	:douta	=	16'h	2924;
53267	:douta	=	16'h	320a;
53268	:douta	=	16'h	428c;
53269	:douta	=	16'h	42ad;
53270	:douta	=	16'h	3a4a;
53271	:douta	=	16'h	2925;
53272	:douta	=	16'h	2082;
53273	:douta	=	16'h	1881;
53274	:douta	=	16'h	1881;
53275	:douta	=	16'h	1881;
53276	:douta	=	16'h	1881;
53277	:douta	=	16'h	20a3;
53278	:douta	=	16'h	20a3;
53279	:douta	=	16'h	2904;
53280	:douta	=	16'h	2924;
53281	:douta	=	16'h	3145;
53282	:douta	=	16'h	39a6;
53283	:douta	=	16'h	39a7;
53284	:douta	=	16'h	4a29;
53285	:douta	=	16'h	4a49;
53286	:douta	=	16'h	52aa;
53287	:douta	=	16'h	630b;
53288	:douta	=	16'h	630b;
53289	:douta	=	16'h	734b;
53290	:douta	=	16'h	734b;
53291	:douta	=	16'h	734b;
53292	:douta	=	16'h	734b;
53293	:douta	=	16'h	6aea;
53294	:douta	=	16'h	39c9;
53295	:douta	=	16'h	10e6;
53296	:douta	=	16'h	6247;
53297	:douta	=	16'h	6246;
53298	:douta	=	16'h	5a25;
53299	:douta	=	16'h	5a05;
53300	:douta	=	16'h	59c4;
53301	:douta	=	16'h	59a4;
53302	:douta	=	16'h	59a3;
53303	:douta	=	16'h	59a3;
53304	:douta	=	16'h	61c4;
53305	:douta	=	16'h	69c3;
53306	:douta	=	16'h	69e3;
53307	:douta	=	16'h	7224;
53308	:douta	=	16'h	7244;
53309	:douta	=	16'h	7244;
53310	:douta	=	16'h	7a64;
53311	:douta	=	16'h	7a64;
53312	:douta	=	16'h	8285;
53313	:douta	=	16'h	7a85;
53314	:douta	=	16'h	82a5;
53315	:douta	=	16'h	8285;
53316	:douta	=	16'h	82a5;
53317	:douta	=	16'h	82a6;
53318	:douta	=	16'h	8ac5;
53319	:douta	=	16'h	51c4;
53320	:douta	=	16'h	6a25;
53321	:douta	=	16'h	8ac6;
53322	:douta	=	16'h	8ae5;
53323	:douta	=	16'h	9306;
53324	:douta	=	16'h	8ac5;
53325	:douta	=	16'h	92e6;
53326	:douta	=	16'h	92e6;
53327	:douta	=	16'h	9306;
53328	:douta	=	16'h	9326;
53329	:douta	=	16'h	9306;
53330	:douta	=	16'h	9b46;
53331	:douta	=	16'h	a366;
53332	:douta	=	16'h	ab87;
53333	:douta	=	16'h	ab86;
53334	:douta	=	16'h	aba6;
53335	:douta	=	16'h	aba6;
53336	:douta	=	16'h	b3c7;
53337	:douta	=	16'h	b3c7;
53338	:douta	=	16'h	b3e6;
53339	:douta	=	16'h	bbe7;
53340	:douta	=	16'h	bbe6;
53341	:douta	=	16'h	bbe6;
53342	:douta	=	16'h	bbe6;
53343	:douta	=	16'h	c3e7;
53344	:douta	=	16'h	c406;
53345	:douta	=	16'h	c407;
53346	:douta	=	16'h	c427;
53347	:douta	=	16'h	c407;
53348	:douta	=	16'h	c427;
53349	:douta	=	16'h	c426;
53350	:douta	=	16'h	cc27;
53351	:douta	=	16'h	c427;
53352	:douta	=	16'h	c427;
53353	:douta	=	16'h	c447;
53354	:douta	=	16'h	cc47;
53355	:douta	=	16'h	cc47;
53356	:douta	=	16'h	cc47;
53357	:douta	=	16'h	cc27;
53358	:douta	=	16'h	cc47;
53359	:douta	=	16'h	cc48;
53360	:douta	=	16'h	cc47;
53361	:douta	=	16'h	cc47;
53362	:douta	=	16'h	cc47;
53363	:douta	=	16'h	cc47;
53364	:douta	=	16'h	cc47;
53365	:douta	=	16'h	cc26;
53366	:douta	=	16'h	c404;
53367	:douta	=	16'h	cc05;
53368	:douta	=	16'h	c403;
53369	:douta	=	16'h	c404;
53370	:douta	=	16'h	cc25;
53371	:douta	=	16'h	c445;
53372	:douta	=	16'h	cc47;
53373	:douta	=	16'h	ccaa;
53374	:douta	=	16'h	d52d;
53375	:douta	=	16'h	d56e;
53376	:douta	=	16'h	ddd1;
53377	:douta	=	16'h	de11;
53378	:douta	=	16'h	de74;
53379	:douta	=	16'h	eed8;
53380	:douta	=	16'h	ef19;
53381	:douta	=	16'h	f77b;
53382	:douta	=	16'h	f77c;
53383	:douta	=	16'h	ffbc;
53384	:douta	=	16'h	ffdc;
53385	:douta	=	16'h	ffdc;
53386	:douta	=	16'h	f79a;
53387	:douta	=	16'h	f77a;
53388	:douta	=	16'h	ef17;
53389	:douta	=	16'h	eeb5;
53390	:douta	=	16'h	e674;
53391	:douta	=	16'h	e611;
53392	:douta	=	16'h	ddef;
53393	:douta	=	16'h	dd8d;
53394	:douta	=	16'h	d52c;
53395	:douta	=	16'h	d50b;
53396	:douta	=	16'h	cca9;
53397	:douta	=	16'h	d489;
53398	:douta	=	16'h	cc67;
53399	:douta	=	16'h	cc46;
53400	:douta	=	16'h	cc47;
53401	:douta	=	16'h	cc47;
53402	:douta	=	16'h	cc47;
53403	:douta	=	16'h	d468;
53404	:douta	=	16'h	d468;
53405	:douta	=	16'h	d488;
53406	:douta	=	16'h	d488;
53407	:douta	=	16'h	cc88;
53408	:douta	=	16'h	d488;
53409	:douta	=	16'h	d488;
53410	:douta	=	16'h	d466;
53411	:douta	=	16'h	ad31;
53412	:douta	=	16'h	deb8;
53413	:douta	=	16'h	cc45;
53414	:douta	=	16'h	cc68;
53415	:douta	=	16'h	d4a9;
53416	:douta	=	16'h	cc89;
53417	:douta	=	16'h	cc88;
53418	:douta	=	16'h	cc68;
53419	:douta	=	16'h	cc88;
53420	:douta	=	16'h	cc68;
53421	:douta	=	16'h	d489;
53422	:douta	=	16'h	cc69;
53423	:douta	=	16'h	cc49;
53424	:douta	=	16'h	d468;
53425	:douta	=	16'h	9430;
53426	:douta	=	16'h	49c5;
53427	:douta	=	16'h	4184;
53428	:douta	=	16'h	5227;
53429	:douta	=	16'h	6b2b;
53430	:douta	=	16'h	838c;
53431	:douta	=	16'h	838c;
53432	:douta	=	16'h	8bcc;
53433	:douta	=	16'h	93ed;
53434	:douta	=	16'h	940d;
53435	:douta	=	16'h	9c8f;
53436	:douta	=	16'h	944e;
53437	:douta	=	16'h	9c6f;
53438	:douta	=	16'h	bd30;
53439	:douta	=	16'h	bd10;
53440	:douta	=	16'h	bd11;
53441	:douta	=	16'h	c572;
53442	:douta	=	16'h	c572;
53443	:douta	=	16'h	cd93;
53444	:douta	=	16'h	d5f4;
53445	:douta	=	16'h	cd73;
53446	:douta	=	16'h	cd93;
53447	:douta	=	16'h	940f;
53448	:douta	=	16'h	bd12;
53449	:douta	=	16'h	cd72;
53450	:douta	=	16'h	cd72;
53451	:douta	=	16'h	a492;
53452	:douta	=	16'h	9c92;
53453	:douta	=	16'h	9433;
53454	:douta	=	16'h	8433;
53455	:douta	=	16'h	73b0;
53456	:douta	=	16'h	6b6f;
53457	:douta	=	16'h	7bb0;
53458	:douta	=	16'h	83f1;
53459	:douta	=	16'h	8411;
53460	:douta	=	16'h	83d1;
53461	:douta	=	16'h	7bd0;
53462	:douta	=	16'h	7bb1;
53463	:douta	=	16'h	6b4f;
53464	:douta	=	16'h	6b4f;
53465	:douta	=	16'h	6b2f;
53466	:douta	=	16'h	6b4e;
53467	:douta	=	16'h	6b2e;
53468	:douta	=	16'h	6b4f;
53469	:douta	=	16'h	7370;
53470	:douta	=	16'h	6b4e;
53471	:douta	=	16'h	6b0d;
53472	:douta	=	16'h	5a8b;
53473	:douta	=	16'h	6b2e;
53474	:douta	=	16'h	6b2e;
53475	:douta	=	16'h	6b4f;
53476	:douta	=	16'h	6b4f;
53477	:douta	=	16'h	6b4f;
53478	:douta	=	16'h	6b6f;
53479	:douta	=	16'h	6b4f;
53480	:douta	=	16'h	6370;
53481	:douta	=	16'h	73f2;
53482	:douta	=	16'h	7413;
53483	:douta	=	16'h	73f3;
53484	:douta	=	16'h	6391;
53485	:douta	=	16'h	4aef;
53486	:douta	=	16'h	7bf1;
53487	:douta	=	16'h	424c;
53488	:douta	=	16'h	2967;
53489	:douta	=	16'h	2168;
53490	:douta	=	16'h	5b6e;
53491	:douta	=	16'h	ffff;
53492	:douta	=	16'h	ffff;
53493	:douta	=	16'h	ffff;
53494	:douta	=	16'h	d5b6;
53495	:douta	=	16'h	9309;
53496	:douta	=	16'h	9b28;
53497	:douta	=	16'h	9b28;
53498	:douta	=	16'h	9328;
53499	:douta	=	16'h	9b28;
53500	:douta	=	16'h	9b28;
53501	:douta	=	16'h	9b28;
53502	:douta	=	16'h	9b28;
53503	:douta	=	16'h	9b28;
53504	:douta	=	16'h	cdd6;
53505	:douta	=	16'h	cdd6;
53506	:douta	=	16'h	cdb6;
53507	:douta	=	16'h	b555;
53508	:douta	=	16'h	9453;
53509	:douta	=	16'h	ad57;
53510	:douta	=	16'h	a515;
53511	:douta	=	16'h	a516;
53512	:douta	=	16'h	9cd5;
53513	:douta	=	16'h	9cf6;
53514	:douta	=	16'h	8c74;
53515	:douta	=	16'h	a558;
53516	:douta	=	16'h	5b2e;
53517	:douta	=	16'h	28e3;
53518	:douta	=	16'h	28e3;
53519	:douta	=	16'h	28e3;
53520	:douta	=	16'h	20e3;
53521	:douta	=	16'h	20c3;
53522	:douta	=	16'h	28e3;
53523	:douta	=	16'h	28c3;
53524	:douta	=	16'h	20a2;
53525	:douta	=	16'h	20e3;
53526	:douta	=	16'h	20e3;
53527	:douta	=	16'h	31c8;
53528	:douta	=	16'h	3a2a;
53529	:douta	=	16'h	39e9;
53530	:douta	=	16'h	31c7;
53531	:douta	=	16'h	31c7;
53532	:douta	=	16'h	31c7;
53533	:douta	=	16'h	31c7;
53534	:douta	=	16'h	31a6;
53535	:douta	=	16'h	3165;
53536	:douta	=	16'h	3165;
53537	:douta	=	16'h	3144;
53538	:douta	=	16'h	3144;
53539	:douta	=	16'h	3124;
53540	:douta	=	16'h	2903;
53541	:douta	=	16'h	3103;
53542	:douta	=	16'h	30e2;
53543	:douta	=	16'h	30e2;
53544	:douta	=	16'h	30e2;
53545	:douta	=	16'h	30e2;
53546	:douta	=	16'h	30e2;
53547	:douta	=	16'h	3902;
53548	:douta	=	16'h	3902;
53549	:douta	=	16'h	41a6;
53550	:douta	=	16'h	2987;
53551	:douta	=	16'h	10a5;
53552	:douta	=	16'h	51a4;
53553	:douta	=	16'h	51a4;
53554	:douta	=	16'h	59c4;
53555	:douta	=	16'h	59c4;
53556	:douta	=	16'h	59c4;
53557	:douta	=	16'h	61e4;
53558	:douta	=	16'h	61e4;
53559	:douta	=	16'h	69e4;
53560	:douta	=	16'h	6a04;
53561	:douta	=	16'h	7224;
53562	:douta	=	16'h	7224;
53563	:douta	=	16'h	7244;
53564	:douta	=	16'h	7a44;
53565	:douta	=	16'h	7a65;
53566	:douta	=	16'h	7a85;
53567	:douta	=	16'h	7a64;
53568	:douta	=	16'h	8285;
53569	:douta	=	16'h	8285;
53570	:douta	=	16'h	8285;
53571	:douta	=	16'h	82a5;
53572	:douta	=	16'h	82c6;
53573	:douta	=	16'h	82c6;
53574	:douta	=	16'h	8ac6;
53575	:douta	=	16'h	6a24;
53576	:douta	=	16'h	51a4;
53577	:douta	=	16'h	8ac6;
53578	:douta	=	16'h	9306;
53579	:douta	=	16'h	9306;
53580	:douta	=	16'h	9306;
53581	:douta	=	16'h	9306;
53582	:douta	=	16'h	9306;
53583	:douta	=	16'h	9306;
53584	:douta	=	16'h	9306;
53585	:douta	=	16'h	9b47;
53586	:douta	=	16'h	9b46;
53587	:douta	=	16'h	ab87;
53588	:douta	=	16'h	ab87;
53589	:douta	=	16'h	aba7;
53590	:douta	=	16'h	b3a7;
53591	:douta	=	16'h	b3a7;
53592	:douta	=	16'h	b3a7;
53593	:douta	=	16'h	b3c7;
53594	:douta	=	16'h	b3e6;
53595	:douta	=	16'h	bbe7;
53596	:douta	=	16'h	bbe7;
53597	:douta	=	16'h	bbe6;
53598	:douta	=	16'h	c3e7;
53599	:douta	=	16'h	c3e7;
53600	:douta	=	16'h	c407;
53601	:douta	=	16'h	c407;
53602	:douta	=	16'h	c407;
53603	:douta	=	16'h	c427;
53604	:douta	=	16'h	c406;
53605	:douta	=	16'h	c406;
53606	:douta	=	16'h	c406;
53607	:douta	=	16'h	c406;
53608	:douta	=	16'h	c404;
53609	:douta	=	16'h	c3e3;
53610	:douta	=	16'h	c3e3;
53611	:douta	=	16'h	c404;
53612	:douta	=	16'h	cc26;
53613	:douta	=	16'h	cc28;
53614	:douta	=	16'h	cc89;
53615	:douta	=	16'h	cccb;
53616	:douta	=	16'h	ccec;
53617	:douta	=	16'h	d56f;
53618	:douta	=	16'h	ddb1;
53619	:douta	=	16'h	de33;
53620	:douta	=	16'h	e6b6;
53621	:douta	=	16'h	eed8;
53622	:douta	=	16'h	ef39;
53623	:douta	=	16'h	f77a;
53624	:douta	=	16'h	f79c;
53625	:douta	=	16'h	f7dc;
53626	:douta	=	16'h	f7bc;
53627	:douta	=	16'h	f79b;
53628	:douta	=	16'h	f77a;
53629	:douta	=	16'h	ef37;
53630	:douta	=	16'h	eed5;
53631	:douta	=	16'h	eeb4;
53632	:douta	=	16'h	e612;
53633	:douta	=	16'h	ddd1;
53634	:douta	=	16'h	d5ae;
53635	:douta	=	16'h	d52c;
53636	:douta	=	16'h	d50b;
53637	:douta	=	16'h	cca8;
53638	:douta	=	16'h	cc88;
53639	:douta	=	16'h	cc66;
53640	:douta	=	16'h	cc46;
53641	:douta	=	16'h	cc26;
53642	:douta	=	16'h	cc46;
53643	:douta	=	16'h	cc45;
53644	:douta	=	16'h	d467;
53645	:douta	=	16'h	d467;
53646	:douta	=	16'h	d468;
53647	:douta	=	16'h	d488;
53648	:douta	=	16'h	d488;
53649	:douta	=	16'h	cc88;
53650	:douta	=	16'h	d488;
53651	:douta	=	16'h	d488;
53652	:douta	=	16'h	cc88;
53653	:douta	=	16'h	d488;
53654	:douta	=	16'h	d488;
53655	:douta	=	16'h	d488;
53656	:douta	=	16'h	d489;
53657	:douta	=	16'h	d488;
53658	:douta	=	16'h	d488;
53659	:douta	=	16'h	cc88;
53660	:douta	=	16'h	d4a9;
53661	:douta	=	16'h	d488;
53662	:douta	=	16'h	d4a9;
53663	:douta	=	16'h	d4a9;
53664	:douta	=	16'h	d488;
53665	:douta	=	16'h	cc69;
53666	:douta	=	16'h	d488;
53667	:douta	=	16'h	ad31;
53668	:douta	=	16'h	deb7;
53669	:douta	=	16'h	cc25;
53670	:douta	=	16'h	d488;
53671	:douta	=	16'h	cc68;
53672	:douta	=	16'h	cc68;
53673	:douta	=	16'h	cc88;
53674	:douta	=	16'h	cc88;
53675	:douta	=	16'h	cc68;
53676	:douta	=	16'h	cc68;
53677	:douta	=	16'h	cc68;
53678	:douta	=	16'h	cc89;
53679	:douta	=	16'h	cc69;
53680	:douta	=	16'h	cc68;
53681	:douta	=	16'h	9beb;
53682	:douta	=	16'h	72c9;
53683	:douta	=	16'h	7b4a;
53684	:douta	=	16'h	836c;
53685	:douta	=	16'h	83ad;
53686	:douta	=	16'h	940e;
53687	:douta	=	16'h	ac90;
53688	:douta	=	16'h	9c4e;
53689	:douta	=	16'h	ac8f;
53690	:douta	=	16'h	b4d0;
53691	:douta	=	16'h	b4f0;
53692	:douta	=	16'h	b4f0;
53693	:douta	=	16'h	c552;
53694	:douta	=	16'h	cd93;
53695	:douta	=	16'h	d5b3;
53696	:douta	=	16'h	cd93;
53697	:douta	=	16'h	cd93;
53698	:douta	=	16'h	cdb4;
53699	:douta	=	16'h	cd53;
53700	:douta	=	16'h	c553;
53701	:douta	=	16'h	b511;
53702	:douta	=	16'h	9c71;
53703	:douta	=	16'h	acb2;
53704	:douta	=	16'h	7bb0;
53705	:douta	=	16'h	83d1;
53706	:douta	=	16'h	8c11;
53707	:douta	=	16'h	9474;
53708	:douta	=	16'h	9473;
53709	:douta	=	16'h	8c74;
53710	:douta	=	16'h	8c53;
53711	:douta	=	16'h	6b70;
53712	:douta	=	16'h	6b6f;
53713	:douta	=	16'h	7b90;
53714	:douta	=	16'h	7b90;
53715	:douta	=	16'h	736f;
53716	:douta	=	16'h	6b4e;
53717	:douta	=	16'h	6b4f;
53718	:douta	=	16'h	6b2e;
53719	:douta	=	16'h	6b6f;
53720	:douta	=	16'h	630e;
53721	:douta	=	16'h	634e;
53722	:douta	=	16'h	6b4f;
53723	:douta	=	16'h	632f;
53724	:douta	=	16'h	630d;
53725	:douta	=	16'h	62cd;
53726	:douta	=	16'h	6b2e;
53727	:douta	=	16'h	62cd;
53728	:douta	=	16'h	630e;
53729	:douta	=	16'h	62cc;
53730	:douta	=	16'h	5a8b;
53731	:douta	=	16'h	62cc;
53732	:douta	=	16'h	62cc;
53733	:douta	=	16'h	6b0d;
53734	:douta	=	16'h	62ed;
53735	:douta	=	16'h	6b4f;
53736	:douta	=	16'h	6370;
53737	:douta	=	16'h	4aad;
53738	:douta	=	16'h	530f;
53739	:douta	=	16'h	6bb1;
53740	:douta	=	16'h	6370;
53741	:douta	=	16'h	8c73;
53742	:douta	=	16'h	4acf;
53743	:douta	=	16'h	4acf;
53744	:douta	=	16'h	5b51;
53745	:douta	=	16'h	39cc;
53746	:douta	=	16'h	d71c;
53747	:douta	=	16'h	ffff;
53748	:douta	=	16'h	ffff;
53749	:douta	=	16'h	ffff;
53750	:douta	=	16'h	ff1a;
53751	:douta	=	16'h	7aa6;
53752	:douta	=	16'h	9b28;
53753	:douta	=	16'h	9b28;
53754	:douta	=	16'h	9b48;
53755	:douta	=	16'h	9b48;
53756	:douta	=	16'h	9b48;
53757	:douta	=	16'h	9b28;
53758	:douta	=	16'h	9b48;
53759	:douta	=	16'h	9b48;
53760	:douta	=	16'h	d5f6;
53761	:douta	=	16'h	cdd6;
53762	:douta	=	16'h	c596;
53763	:douta	=	16'h	ad15;
53764	:douta	=	16'h	9cb4;
53765	:douta	=	16'h	b577;
53766	:douta	=	16'h	a4f5;
53767	:douta	=	16'h	a4f5;
53768	:douta	=	16'h	9cd5;
53769	:douta	=	16'h	94d5;
53770	:douta	=	16'h	8434;
53771	:douta	=	16'h	94d6;
53772	:douta	=	16'h	3166;
53773	:douta	=	16'h	20e3;
53774	:douta	=	16'h	20e3;
53775	:douta	=	16'h	20e3;
53776	:douta	=	16'h	20c3;
53777	:douta	=	16'h	20c3;
53778	:douta	=	16'h	28e3;
53779	:douta	=	16'h	20e3;
53780	:douta	=	16'h	20c3;
53781	:douta	=	16'h	20c3;
53782	:douta	=	16'h	20a3;
53783	:douta	=	16'h	20c3;
53784	:douta	=	16'h	20e3;
53785	:douta	=	16'h	20e3;
53786	:douta	=	16'h	2103;
53787	:douta	=	16'h	2103;
53788	:douta	=	16'h	20a3;
53789	:douta	=	16'h	20c3;
53790	:douta	=	16'h	20c3;
53791	:douta	=	16'h	20a2;
53792	:douta	=	16'h	20a2;
53793	:douta	=	16'h	20a1;
53794	:douta	=	16'h	20a2;
53795	:douta	=	16'h	28a2;
53796	:douta	=	16'h	28c2;
53797	:douta	=	16'h	28c2;
53798	:douta	=	16'h	28c2;
53799	:douta	=	16'h	30e2;
53800	:douta	=	16'h	3102;
53801	:douta	=	16'h	3923;
53802	:douta	=	16'h	3903;
53803	:douta	=	16'h	4123;
53804	:douta	=	16'h	4123;
53805	:douta	=	16'h	49e7;
53806	:douta	=	16'h	2947;
53807	:douta	=	16'h	0884;
53808	:douta	=	16'h	5184;
53809	:douta	=	16'h	59a4;
53810	:douta	=	16'h	59c4;
53811	:douta	=	16'h	59c4;
53812	:douta	=	16'h	59c4;
53813	:douta	=	16'h	61e4;
53814	:douta	=	16'h	61e4;
53815	:douta	=	16'h	6204;
53816	:douta	=	16'h	6a24;
53817	:douta	=	16'h	6a24;
53818	:douta	=	16'h	7224;
53819	:douta	=	16'h	7244;
53820	:douta	=	16'h	7a65;
53821	:douta	=	16'h	7a64;
53822	:douta	=	16'h	7a64;
53823	:douta	=	16'h	7a85;
53824	:douta	=	16'h	7a85;
53825	:douta	=	16'h	8285;
53826	:douta	=	16'h	8285;
53827	:douta	=	16'h	82a6;
53828	:douta	=	16'h	8aa6;
53829	:douta	=	16'h	82c6;
53830	:douta	=	16'h	82c6;
53831	:douta	=	16'h	7a85;
53832	:douta	=	16'h	5184;
53833	:douta	=	16'h	92e6;
53834	:douta	=	16'h	8ac5;
53835	:douta	=	16'h	9306;
53836	:douta	=	16'h	9306;
53837	:douta	=	16'h	9306;
53838	:douta	=	16'h	9306;
53839	:douta	=	16'h	9306;
53840	:douta	=	16'h	9326;
53841	:douta	=	16'h	9326;
53842	:douta	=	16'h	9b26;
53843	:douta	=	16'h	a366;
53844	:douta	=	16'h	ab87;
53845	:douta	=	16'h	ab86;
53846	:douta	=	16'h	b3c6;
53847	:douta	=	16'h	b3a6;
53848	:douta	=	16'h	b3c6;
53849	:douta	=	16'h	b3c6;
53850	:douta	=	16'h	b3c7;
53851	:douta	=	16'h	bbe6;
53852	:douta	=	16'h	b3c6;
53853	:douta	=	16'h	bbe7;
53854	:douta	=	16'h	bbe6;
53855	:douta	=	16'h	bbe6;
53856	:douta	=	16'h	bbc5;
53857	:douta	=	16'h	bbe5;
53858	:douta	=	16'h	bba4;
53859	:douta	=	16'h	c3c4;
53860	:douta	=	16'h	bbc4;
53861	:douta	=	16'h	bc05;
53862	:douta	=	16'h	c426;
53863	:douta	=	16'h	c468;
53864	:douta	=	16'h	c4a9;
53865	:douta	=	16'h	cced;
53866	:douta	=	16'h	d58f;
53867	:douta	=	16'h	d5d1;
53868	:douta	=	16'h	de54;
53869	:douta	=	16'h	e675;
53870	:douta	=	16'h	eef8;
53871	:douta	=	16'h	ef59;
53872	:douta	=	16'h	f77a;
53873	:douta	=	16'h	f79b;
53874	:douta	=	16'h	f7bc;
53875	:douta	=	16'h	f7bb;
53876	:douta	=	16'h	f77a;
53877	:douta	=	16'h	f759;
53878	:douta	=	16'h	eef6;
53879	:douta	=	16'h	e6b6;
53880	:douta	=	16'h	e673;
53881	:douta	=	16'h	ddd0;
53882	:douta	=	16'h	ddaf;
53883	:douta	=	16'h	d54d;
53884	:douta	=	16'h	d52b;
53885	:douta	=	16'h	ccea;
53886	:douta	=	16'h	cca8;
53887	:douta	=	16'h	cc88;
53888	:douta	=	16'h	cc46;
53889	:douta	=	16'h	cc46;
53890	:douta	=	16'h	cc25;
53891	:douta	=	16'h	cc46;
53892	:douta	=	16'h	cc46;
53893	:douta	=	16'h	cc47;
53894	:douta	=	16'h	cc47;
53895	:douta	=	16'h	cc68;
53896	:douta	=	16'h	d488;
53897	:douta	=	16'h	cc88;
53898	:douta	=	16'h	cc88;
53899	:douta	=	16'h	cc88;
53900	:douta	=	16'h	cc88;
53901	:douta	=	16'h	d488;
53902	:douta	=	16'h	d488;
53903	:douta	=	16'h	cc88;
53904	:douta	=	16'h	cc88;
53905	:douta	=	16'h	d488;
53906	:douta	=	16'h	cc88;
53907	:douta	=	16'h	d488;
53908	:douta	=	16'h	cc88;
53909	:douta	=	16'h	d488;
53910	:douta	=	16'h	d4a9;
53911	:douta	=	16'h	cc68;
53912	:douta	=	16'h	d469;
53913	:douta	=	16'h	d488;
53914	:douta	=	16'h	d488;
53915	:douta	=	16'h	cc69;
53916	:douta	=	16'h	d488;
53917	:douta	=	16'h	d488;
53918	:douta	=	16'h	d488;
53919	:douta	=	16'h	d488;
53920	:douta	=	16'h	d4a9;
53921	:douta	=	16'h	cc88;
53922	:douta	=	16'h	d487;
53923	:douta	=	16'h	ad11;
53924	:douta	=	16'h	deb8;
53925	:douta	=	16'h	cc05;
53926	:douta	=	16'h	cc88;
53927	:douta	=	16'h	cc88;
53928	:douta	=	16'h	cc88;
53929	:douta	=	16'h	cc88;
53930	:douta	=	16'h	cc68;
53931	:douta	=	16'h	cc68;
53932	:douta	=	16'h	cc68;
53933	:douta	=	16'h	cc68;
53934	:douta	=	16'h	cc68;
53935	:douta	=	16'h	cc69;
53936	:douta	=	16'h	cc68;
53937	:douta	=	16'h	a3ea;
53938	:douta	=	16'h	730a;
53939	:douta	=	16'h	8bac;
53940	:douta	=	16'h	8bee;
53941	:douta	=	16'h	8bcd;
53942	:douta	=	16'h	acb0;
53943	:douta	=	16'h	ac90;
53944	:douta	=	16'h	a490;
53945	:douta	=	16'h	bd11;
53946	:douta	=	16'h	c552;
53947	:douta	=	16'h	bd11;
53948	:douta	=	16'h	c553;
53949	:douta	=	16'h	c593;
53950	:douta	=	16'h	cdb4;
53951	:douta	=	16'h	d5d4;
53952	:douta	=	16'h	d5b4;
53953	:douta	=	16'h	c553;
53954	:douta	=	16'h	c573;
53955	:douta	=	16'h	bd12;
53956	:douta	=	16'h	acd3;
53957	:douta	=	16'h	a4d2;
53958	:douta	=	16'h	8c12;
53959	:douta	=	16'h	8bf1;
53960	:douta	=	16'h	9452;
53961	:douta	=	16'h	9452;
53962	:douta	=	16'h	83b0;
53963	:douta	=	16'h	8c53;
53964	:douta	=	16'h	9474;
53965	:douta	=	16'h	7bf1;
53966	:douta	=	16'h	7bf2;
53967	:douta	=	16'h	7390;
53968	:douta	=	16'h	632f;
53969	:douta	=	16'h	738f;
53970	:douta	=	16'h	6b2e;
53971	:douta	=	16'h	734f;
53972	:douta	=	16'h	630d;
53973	:douta	=	16'h	62ed;
53974	:douta	=	16'h	630e;
53975	:douta	=	16'h	6b2e;
53976	:douta	=	16'h	630e;
53977	:douta	=	16'h	5aed;
53978	:douta	=	16'h	5acd;
53979	:douta	=	16'h	528c;
53980	:douta	=	16'h	734f;
53981	:douta	=	16'h	62ed;
53982	:douta	=	16'h	62cd;
53983	:douta	=	16'h	62ed;
53984	:douta	=	16'h	5a6b;
53985	:douta	=	16'h	5a8b;
53986	:douta	=	16'h	528a;
53987	:douta	=	16'h	49e9;
53988	:douta	=	16'h	7b6f;
53989	:douta	=	16'h	6b0e;
53990	:douta	=	16'h	62ac;
53991	:douta	=	16'h	62ed;
53992	:douta	=	16'h	5b0e;
53993	:douta	=	16'h	4ace;
53994	:douta	=	16'h	320b;
53995	:douta	=	16'h	8433;
53996	:douta	=	16'h	7390;
53997	:douta	=	16'h	5b2f;
53998	:douta	=	16'h	6bb3;
53999	:douta	=	16'h	5b72;
54000	:douta	=	16'h	53d3;
54001	:douta	=	16'h	5c13;
54002	:douta	=	16'h	ffff;
54003	:douta	=	16'h	feba;
54004	:douta	=	16'h	ee58;
54005	:douta	=	16'h	c4b0;
54006	:douta	=	16'h	ab49;
54007	:douta	=	16'h	a349;
54008	:douta	=	16'h	9b29;
54009	:douta	=	16'h	9b28;
54010	:douta	=	16'h	9b48;
54011	:douta	=	16'h	9b48;
54012	:douta	=	16'h	9b48;
54013	:douta	=	16'h	9b48;
54014	:douta	=	16'h	9b48;
54015	:douta	=	16'h	9b48;
54016	:douta	=	16'h	de16;
54017	:douta	=	16'h	c595;
54018	:douta	=	16'h	bd55;
54019	:douta	=	16'h	9494;
54020	:douta	=	16'h	ad36;
54021	:douta	=	16'h	ad36;
54022	:douta	=	16'h	a515;
54023	:douta	=	16'h	a4f5;
54024	:douta	=	16'h	9cd5;
54025	:douta	=	16'h	8c94;
54026	:douta	=	16'h	8cb6;
54027	:douta	=	16'h	31c7;
54028	:douta	=	16'h	1040;
54029	:douta	=	16'h	28e4;
54030	:douta	=	16'h	28e3;
54031	:douta	=	16'h	28e3;
54032	:douta	=	16'h	28e3;
54033	:douta	=	16'h	28e3;
54034	:douta	=	16'h	28e3;
54035	:douta	=	16'h	20e3;
54036	:douta	=	16'h	20e3;
54037	:douta	=	16'h	20e3;
54038	:douta	=	16'h	20e3;
54039	:douta	=	16'h	20e3;
54040	:douta	=	16'h	20e3;
54041	:douta	=	16'h	18a2;
54042	:douta	=	16'h	20a2;
54043	:douta	=	16'h	20a2;
54044	:douta	=	16'h	20a2;
54045	:douta	=	16'h	20c2;
54046	:douta	=	16'h	20a2;
54047	:douta	=	16'h	20a2;
54048	:douta	=	16'h	20a2;
54049	:douta	=	16'h	20c2;
54050	:douta	=	16'h	28e2;
54051	:douta	=	16'h	28e3;
54052	:douta	=	16'h	30e3;
54053	:douta	=	16'h	28e3;
54054	:douta	=	16'h	3103;
54055	:douta	=	16'h	3123;
54056	:douta	=	16'h	3903;
54057	:douta	=	16'h	3943;
54058	:douta	=	16'h	4123;
54059	:douta	=	16'h	4144;
54060	:douta	=	16'h	4165;
54061	:douta	=	16'h	4a49;
54062	:douta	=	16'h	2126;
54063	:douta	=	16'h	18a5;
54064	:douta	=	16'h	59a4;
54065	:douta	=	16'h	51a4;
54066	:douta	=	16'h	51a4;
54067	:douta	=	16'h	61e4;
54068	:douta	=	16'h	61c4;
54069	:douta	=	16'h	61e4;
54070	:douta	=	16'h	6204;
54071	:douta	=	16'h	6a04;
54072	:douta	=	16'h	6a04;
54073	:douta	=	16'h	7224;
54074	:douta	=	16'h	7244;
54075	:douta	=	16'h	7a64;
54076	:douta	=	16'h	7a64;
54077	:douta	=	16'h	7a65;
54078	:douta	=	16'h	7a85;
54079	:douta	=	16'h	8286;
54080	:douta	=	16'h	82a5;
54081	:douta	=	16'h	7a85;
54082	:douta	=	16'h	82a6;
54083	:douta	=	16'h	82a5;
54084	:douta	=	16'h	82c6;
54085	:douta	=	16'h	82c5;
54086	:douta	=	16'h	8ac6;
54087	:douta	=	16'h	9326;
54088	:douta	=	16'h	61e5;
54089	:douta	=	16'h	9b26;
54090	:douta	=	16'h	9306;
54091	:douta	=	16'h	9306;
54092	:douta	=	16'h	9305;
54093	:douta	=	16'h	9305;
54094	:douta	=	16'h	92e6;
54095	:douta	=	16'h	9326;
54096	:douta	=	16'h	9306;
54097	:douta	=	16'h	9306;
54098	:douta	=	16'h	9b05;
54099	:douta	=	16'h	a326;
54100	:douta	=	16'h	a325;
54101	:douta	=	16'h	a325;
54102	:douta	=	16'h	ab45;
54103	:douta	=	16'h	ab64;
54104	:douta	=	16'h	ab85;
54105	:douta	=	16'h	b3c6;
54106	:douta	=	16'h	bc08;
54107	:douta	=	16'h	c4ac;
54108	:douta	=	16'h	c50d;
54109	:douta	=	16'h	cd70;
54110	:douta	=	16'h	d5b1;
54111	:douta	=	16'h	de53;
54112	:douta	=	16'h	e6d6;
54113	:douta	=	16'h	e718;
54114	:douta	=	16'h	ef7a;
54115	:douta	=	16'h	f77a;
54116	:douta	=	16'h	f7bb;
54117	:douta	=	16'h	f79a;
54118	:douta	=	16'h	f77a;
54119	:douta	=	16'h	ef38;
54120	:douta	=	16'h	eef6;
54121	:douta	=	16'h	e6b4;
54122	:douta	=	16'h	de32;
54123	:douta	=	16'h	ddf1;
54124	:douta	=	16'h	d58e;
54125	:douta	=	16'h	cd4d;
54126	:douta	=	16'h	ccea;
54127	:douta	=	16'h	cca8;
54128	:douta	=	16'h	c468;
54129	:douta	=	16'h	cc46;
54130	:douta	=	16'h	c425;
54131	:douta	=	16'h	cc25;
54132	:douta	=	16'h	cc25;
54133	:douta	=	16'h	cc25;
54134	:douta	=	16'h	cc46;
54135	:douta	=	16'h	cc46;
54136	:douta	=	16'h	cc67;
54137	:douta	=	16'h	cc67;
54138	:douta	=	16'h	cc68;
54139	:douta	=	16'h	cc67;
54140	:douta	=	16'h	cc68;
54141	:douta	=	16'h	cc68;
54142	:douta	=	16'h	d488;
54143	:douta	=	16'h	cc67;
54144	:douta	=	16'h	cc68;
54145	:douta	=	16'h	cc68;
54146	:douta	=	16'h	cc68;
54147	:douta	=	16'h	d488;
54148	:douta	=	16'h	cc68;
54149	:douta	=	16'h	cc68;
54150	:douta	=	16'h	cc68;
54151	:douta	=	16'h	cc88;
54152	:douta	=	16'h	cc88;
54153	:douta	=	16'h	cc88;
54154	:douta	=	16'h	cc88;
54155	:douta	=	16'h	cc88;
54156	:douta	=	16'h	d488;
54157	:douta	=	16'h	d488;
54158	:douta	=	16'h	cc88;
54159	:douta	=	16'h	cc88;
54160	:douta	=	16'h	cc88;
54161	:douta	=	16'h	cc88;
54162	:douta	=	16'h	d4a9;
54163	:douta	=	16'h	cc88;
54164	:douta	=	16'h	d4a9;
54165	:douta	=	16'h	d488;
54166	:douta	=	16'h	cc88;
54167	:douta	=	16'h	d4a9;
54168	:douta	=	16'h	d489;
54169	:douta	=	16'h	d489;
54170	:douta	=	16'h	d489;
54171	:douta	=	16'h	d4a9;
54172	:douta	=	16'h	d4a9;
54173	:douta	=	16'h	d488;
54174	:douta	=	16'h	d4a9;
54175	:douta	=	16'h	d488;
54176	:douta	=	16'h	d488;
54177	:douta	=	16'h	d488;
54178	:douta	=	16'h	d487;
54179	:douta	=	16'h	ad31;
54180	:douta	=	16'h	ded7;
54181	:douta	=	16'h	cc26;
54182	:douta	=	16'h	cc68;
54183	:douta	=	16'h	cc68;
54184	:douta	=	16'h	cc88;
54185	:douta	=	16'h	cc68;
54186	:douta	=	16'h	cc88;
54187	:douta	=	16'h	cc88;
54188	:douta	=	16'h	cc88;
54189	:douta	=	16'h	cc68;
54190	:douta	=	16'h	d488;
54191	:douta	=	16'h	cc68;
54192	:douta	=	16'h	cc88;
54193	:douta	=	16'h	a40a;
54194	:douta	=	16'h	8bad;
54195	:douta	=	16'h	8bcd;
54196	:douta	=	16'h	93ee;
54197	:douta	=	16'h	9c2f;
54198	:douta	=	16'h	bd32;
54199	:douta	=	16'h	bd12;
54200	:douta	=	16'h	bd33;
54201	:douta	=	16'h	c553;
54202	:douta	=	16'h	c573;
54203	:douta	=	16'h	bd73;
54204	:douta	=	16'h	cdb5;
54205	:douta	=	16'h	cdb4;
54206	:douta	=	16'h	d5d4;
54207	:douta	=	16'h	cd92;
54208	:douta	=	16'h	cd73;
54209	:douta	=	16'h	acd2;
54210	:douta	=	16'h	b4d3;
54211	:douta	=	16'h	8c32;
54212	:douta	=	16'h	9453;
54213	:douta	=	16'h	9432;
54214	:douta	=	16'h	9473;
54215	:douta	=	16'h	8c32;
54216	:douta	=	16'h	7bb0;
54217	:douta	=	16'h	83f2;
54218	:douta	=	16'h	6b4f;
54219	:douta	=	16'h	7bb0;
54220	:douta	=	16'h	732f;
54221	:douta	=	16'h	630d;
54222	:douta	=	16'h	6b2e;
54223	:douta	=	16'h	630e;
54224	:douta	=	16'h	632e;
54225	:douta	=	16'h	62ed;
54226	:douta	=	16'h	8432;
54227	:douta	=	16'h	736f;
54228	:douta	=	16'h	62ed;
54229	:douta	=	16'h	5acc;
54230	:douta	=	16'h	4a2a;
54231	:douta	=	16'h	5acc;
54232	:douta	=	16'h	62cc;
54233	:douta	=	16'h	5aab;
54234	:douta	=	16'h	5a8b;
54235	:douta	=	16'h	526a;
54236	:douta	=	16'h	41e8;
54237	:douta	=	16'h	62ac;
54238	:douta	=	16'h	736f;
54239	:douta	=	16'h	8c32;
54240	:douta	=	16'h	9453;
54241	:douta	=	16'h	8413;
54242	:douta	=	16'h	8c74;
54243	:douta	=	16'h	8432;
54244	:douta	=	16'h	6b4f;
54245	:douta	=	16'h	632f;
54246	:douta	=	16'h	6b2e;
54247	:douta	=	16'h	634e;
54248	:douta	=	16'h	9c92;
54249	:douta	=	16'h	b5d7;
54250	:douta	=	16'h	a575;
54251	:douta	=	16'h	6c94;
54252	:douta	=	16'h	8557;
54253	:douta	=	16'h	ce7b;
54254	:douta	=	16'h	cdb3;
54255	:douta	=	16'h	ddb2;
54256	:douta	=	16'h	c388;
54257	:douta	=	16'h	b2c5;
54258	:douta	=	16'h	9ac4;
54259	:douta	=	16'h	a368;
54260	:douta	=	16'h	a368;
54261	:douta	=	16'h	a368;
54262	:douta	=	16'h	9b47;
54263	:douta	=	16'h	a369;
54264	:douta	=	16'h	a369;
54265	:douta	=	16'h	a369;
54266	:douta	=	16'h	9b48;
54267	:douta	=	16'h	9b48;
54268	:douta	=	16'h	9b48;
54269	:douta	=	16'h	a349;
54270	:douta	=	16'h	9b48;
54271	:douta	=	16'h	9b48;
54272	:douta	=	16'h	d616;
54273	:douta	=	16'h	bd95;
54274	:douta	=	16'h	bd96;
54275	:douta	=	16'h	8433;
54276	:douta	=	16'h	b577;
54277	:douta	=	16'h	a536;
54278	:douta	=	16'h	a4f5;
54279	:douta	=	16'h	9cf5;
54280	:douta	=	16'h	a4d5;
54281	:douta	=	16'h	8474;
54282	:douta	=	16'h	a539;
54283	:douta	=	16'h	1881;
54284	:douta	=	16'h	28e3;
54285	:douta	=	16'h	28e3;
54286	:douta	=	16'h	28e3;
54287	:douta	=	16'h	28e3;
54288	:douta	=	16'h	20e3;
54289	:douta	=	16'h	28e3;
54290	:douta	=	16'h	20c3;
54291	:douta	=	16'h	20c3;
54292	:douta	=	16'h	28e3;
54293	:douta	=	16'h	20e3;
54294	:douta	=	16'h	20e3;
54295	:douta	=	16'h	20c3;
54296	:douta	=	16'h	20e3;
54297	:douta	=	16'h	1881;
54298	:douta	=	16'h	20c2;
54299	:douta	=	16'h	2082;
54300	:douta	=	16'h	20a2;
54301	:douta	=	16'h	20c2;
54302	:douta	=	16'h	20a2;
54303	:douta	=	16'h	20a2;
54304	:douta	=	16'h	20a2;
54305	:douta	=	16'h	20c2;
54306	:douta	=	16'h	28e3;
54307	:douta	=	16'h	28e3;
54308	:douta	=	16'h	30e3;
54309	:douta	=	16'h	28e3;
54310	:douta	=	16'h	3123;
54311	:douta	=	16'h	3103;
54312	:douta	=	16'h	3923;
54313	:douta	=	16'h	3923;
54314	:douta	=	16'h	4143;
54315	:douta	=	16'h	4143;
54316	:douta	=	16'h	4185;
54317	:douta	=	16'h	4a4a;
54318	:douta	=	16'h	1905;
54319	:douta	=	16'h	20c5;
54320	:douta	=	16'h	51a4;
54321	:douta	=	16'h	51a4;
54322	:douta	=	16'h	59e4;
54323	:douta	=	16'h	59c4;
54324	:douta	=	16'h	61c4;
54325	:douta	=	16'h	61e4;
54326	:douta	=	16'h	61e4;
54327	:douta	=	16'h	69e4;
54328	:douta	=	16'h	6a04;
54329	:douta	=	16'h	7224;
54330	:douta	=	16'h	7244;
54331	:douta	=	16'h	7a65;
54332	:douta	=	16'h	7a65;
54333	:douta	=	16'h	7a64;
54334	:douta	=	16'h	7a85;
54335	:douta	=	16'h	82a5;
54336	:douta	=	16'h	8285;
54337	:douta	=	16'h	82a5;
54338	:douta	=	16'h	8aa6;
54339	:douta	=	16'h	8aa6;
54340	:douta	=	16'h	82c6;
54341	:douta	=	16'h	82c6;
54342	:douta	=	16'h	8ac6;
54343	:douta	=	16'h	9306;
54344	:douta	=	16'h	6a25;
54345	:douta	=	16'h	9305;
54346	:douta	=	16'h	8ac4;
54347	:douta	=	16'h	8ac4;
54348	:douta	=	16'h	8aa4;
54349	:douta	=	16'h	8aa4;
54350	:douta	=	16'h	8a84;
54351	:douta	=	16'h	8aa5;
54352	:douta	=	16'h	8ac6;
54353	:douta	=	16'h	9305;
54354	:douta	=	16'h	9b67;
54355	:douta	=	16'h	a3e8;
54356	:douta	=	16'h	b46b;
54357	:douta	=	16'h	bcac;
54358	:douta	=	16'h	cd4f;
54359	:douta	=	16'h	cd90;
54360	:douta	=	16'h	de13;
54361	:douta	=	16'h	de53;
54362	:douta	=	16'h	e6b6;
54363	:douta	=	16'h	ef38;
54364	:douta	=	16'h	ef59;
54365	:douta	=	16'h	f779;
54366	:douta	=	16'h	f77a;
54367	:douta	=	16'h	ef59;
54368	:douta	=	16'h	eef7;
54369	:douta	=	16'h	e6b5;
54370	:douta	=	16'h	e653;
54371	:douta	=	16'h	de32;
54372	:douta	=	16'h	d5d0;
54373	:douta	=	16'h	d56e;
54374	:douta	=	16'h	cd2d;
54375	:douta	=	16'h	ccca;
54376	:douta	=	16'h	cca9;
54377	:douta	=	16'h	c467;
54378	:douta	=	16'h	c425;
54379	:douta	=	16'h	c425;
54380	:douta	=	16'h	c404;
54381	:douta	=	16'h	c404;
54382	:douta	=	16'h	cc07;
54383	:douta	=	16'h	cc27;
54384	:douta	=	16'h	cc26;
54385	:douta	=	16'h	cc67;
54386	:douta	=	16'h	cc67;
54387	:douta	=	16'h	cc67;
54388	:douta	=	16'h	cc67;
54389	:douta	=	16'h	cc67;
54390	:douta	=	16'h	cc67;
54391	:douta	=	16'h	cc67;
54392	:douta	=	16'h	cc67;
54393	:douta	=	16'h	cc67;
54394	:douta	=	16'h	cc67;
54395	:douta	=	16'h	cc67;
54396	:douta	=	16'h	cc68;
54397	:douta	=	16'h	cc68;
54398	:douta	=	16'h	cc68;
54399	:douta	=	16'h	cc68;
54400	:douta	=	16'h	d488;
54401	:douta	=	16'h	cc88;
54402	:douta	=	16'h	cc68;
54403	:douta	=	16'h	cc68;
54404	:douta	=	16'h	cc68;
54405	:douta	=	16'h	cc88;
54406	:douta	=	16'h	cc68;
54407	:douta	=	16'h	cc88;
54408	:douta	=	16'h	cc88;
54409	:douta	=	16'h	cc88;
54410	:douta	=	16'h	d488;
54411	:douta	=	16'h	cc88;
54412	:douta	=	16'h	cc88;
54413	:douta	=	16'h	d488;
54414	:douta	=	16'h	d488;
54415	:douta	=	16'h	cc88;
54416	:douta	=	16'h	cc88;
54417	:douta	=	16'h	d488;
54418	:douta	=	16'h	d488;
54419	:douta	=	16'h	cc88;
54420	:douta	=	16'h	cc88;
54421	:douta	=	16'h	d488;
54422	:douta	=	16'h	cc88;
54423	:douta	=	16'h	d488;
54424	:douta	=	16'h	d4a9;
54425	:douta	=	16'h	cc89;
54426	:douta	=	16'h	d488;
54427	:douta	=	16'h	cc88;
54428	:douta	=	16'h	d488;
54429	:douta	=	16'h	cc88;
54430	:douta	=	16'h	cc88;
54431	:douta	=	16'h	d488;
54432	:douta	=	16'h	d488;
54433	:douta	=	16'h	d488;
54434	:douta	=	16'h	d487;
54435	:douta	=	16'h	ad31;
54436	:douta	=	16'h	e6d8;
54437	:douta	=	16'h	cc25;
54438	:douta	=	16'h	cc88;
54439	:douta	=	16'h	cc88;
54440	:douta	=	16'h	cc68;
54441	:douta	=	16'h	cc68;
54442	:douta	=	16'h	cc88;
54443	:douta	=	16'h	cc88;
54444	:douta	=	16'h	cc88;
54445	:douta	=	16'h	cc88;
54446	:douta	=	16'h	cc88;
54447	:douta	=	16'h	cc88;
54448	:douta	=	16'h	cc68;
54449	:douta	=	16'h	ac0a;
54450	:douta	=	16'h	93ee;
54451	:douta	=	16'h	940e;
54452	:douta	=	16'h	940e;
54453	:douta	=	16'h	a450;
54454	:douta	=	16'h	bd32;
54455	:douta	=	16'h	bd32;
54456	:douta	=	16'h	c573;
54457	:douta	=	16'h	c574;
54458	:douta	=	16'h	bd33;
54459	:douta	=	16'h	c594;
54460	:douta	=	16'h	cdd5;
54461	:douta	=	16'h	cd94;
54462	:douta	=	16'h	c553;
54463	:douta	=	16'h	bd13;
54464	:douta	=	16'h	b4d3;
54465	:douta	=	16'h	acb3;
54466	:douta	=	16'h	a492;
54467	:douta	=	16'h	8412;
54468	:douta	=	16'h	8432;
54469	:douta	=	16'h	7bd1;
54470	:douta	=	16'h	83f1;
54471	:douta	=	16'h	8412;
54472	:douta	=	16'h	7390;
54473	:douta	=	16'h	7b90;
54474	:douta	=	16'h	632e;
54475	:douta	=	16'h	7bb0;
54476	:douta	=	16'h	736f;
54477	:douta	=	16'h	6b2e;
54478	:douta	=	16'h	6b2e;
54479	:douta	=	16'h	62ed;
54480	:douta	=	16'h	6b4e;
54481	:douta	=	16'h	632e;
54482	:douta	=	16'h	7c12;
54483	:douta	=	16'h	6b6f;
54484	:douta	=	16'h	6b0d;
54485	:douta	=	16'h	5aad;
54486	:douta	=	16'h	526c;
54487	:douta	=	16'h	526b;
54488	:douta	=	16'h	52ab;
54489	:douta	=	16'h	62ac;
54490	:douta	=	16'h	6b2e;
54491	:douta	=	16'h	736f;
54492	:douta	=	16'h	8bf0;
54493	:douta	=	16'h	8c31;
54494	:douta	=	16'h	8c73;
54495	:douta	=	16'h	632f;
54496	:douta	=	16'h	528d;
54497	:douta	=	16'h	7391;
54498	:douta	=	16'h	7bb1;
54499	:douta	=	16'h	630e;
54500	:douta	=	16'h	52ce;
54501	:douta	=	16'h	636f;
54502	:douta	=	16'h	9d55;
54503	:douta	=	16'h	c67a;
54504	:douta	=	16'h	f7ff;
54505	:douta	=	16'h	ffff;
54506	:douta	=	16'h	ffff;
54507	:douta	=	16'h	fefa;
54508	:douta	=	16'h	f636;
54509	:douta	=	16'h	dcad;
54510	:douta	=	16'h	bb47;
54511	:douta	=	16'h	9aa3;
54512	:douta	=	16'h	9b47;
54513	:douta	=	16'h	9b67;
54514	:douta	=	16'h	a388;
54515	:douta	=	16'h	a368;
54516	:douta	=	16'h	a368;
54517	:douta	=	16'h	9b47;
54518	:douta	=	16'h	a368;
54519	:douta	=	16'h	a368;
54520	:douta	=	16'h	a349;
54521	:douta	=	16'h	a348;
54522	:douta	=	16'h	a348;
54523	:douta	=	16'h	a348;
54524	:douta	=	16'h	9b48;
54525	:douta	=	16'h	a348;
54526	:douta	=	16'h	a348;
54527	:douta	=	16'h	9b48;
54528	:douta	=	16'h	cdd6;
54529	:douta	=	16'h	bd95;
54530	:douta	=	16'h	b556;
54531	:douta	=	16'h	8c53;
54532	:douta	=	16'h	ad57;
54533	:douta	=	16'h	a515;
54534	:douta	=	16'h	a4f5;
54535	:douta	=	16'h	a4d5;
54536	:douta	=	16'h	9cd5;
54537	:douta	=	16'h	9d38;
54538	:douta	=	16'h	7c74;
54539	:douta	=	16'h	2041;
54540	:douta	=	16'h	2082;
54541	:douta	=	16'h	28e3;
54542	:douta	=	16'h	20e3;
54543	:douta	=	16'h	28e3;
54544	:douta	=	16'h	28e3;
54545	:douta	=	16'h	28e3;
54546	:douta	=	16'h	2904;
54547	:douta	=	16'h	28e3;
54548	:douta	=	16'h	28e3;
54549	:douta	=	16'h	20e3;
54550	:douta	=	16'h	20e3;
54551	:douta	=	16'h	20e3;
54552	:douta	=	16'h	20a2;
54553	:douta	=	16'h	1882;
54554	:douta	=	16'h	20a2;
54555	:douta	=	16'h	20a2;
54556	:douta	=	16'h	20a2;
54557	:douta	=	16'h	20a2;
54558	:douta	=	16'h	20a2;
54559	:douta	=	16'h	20a2;
54560	:douta	=	16'h	20a2;
54561	:douta	=	16'h	28e3;
54562	:douta	=	16'h	28c2;
54563	:douta	=	16'h	28e3;
54564	:douta	=	16'h	28e2;
54565	:douta	=	16'h	3103;
54566	:douta	=	16'h	3103;
54567	:douta	=	16'h	3123;
54568	:douta	=	16'h	3923;
54569	:douta	=	16'h	3944;
54570	:douta	=	16'h	3923;
54571	:douta	=	16'h	4143;
54572	:douta	=	16'h	41c7;
54573	:douta	=	16'h	424a;
54574	:douta	=	16'h	18a5;
54575	:douta	=	16'h	3104;
54576	:douta	=	16'h	51a4;
54577	:douta	=	16'h	59a4;
54578	:douta	=	16'h	59c4;
54579	:douta	=	16'h	61c4;
54580	:douta	=	16'h	61e4;
54581	:douta	=	16'h	6204;
54582	:douta	=	16'h	61e4;
54583	:douta	=	16'h	6a24;
54584	:douta	=	16'h	6a04;
54585	:douta	=	16'h	7224;
54586	:douta	=	16'h	7224;
54587	:douta	=	16'h	7a64;
54588	:douta	=	16'h	7244;
54589	:douta	=	16'h	7a44;
54590	:douta	=	16'h	7224;
54591	:douta	=	16'h	7a24;
54592	:douta	=	16'h	7a24;
54593	:douta	=	16'h	7a44;
54594	:douta	=	16'h	7a64;
54595	:douta	=	16'h	8285;
54596	:douta	=	16'h	82c7;
54597	:douta	=	16'h	8b28;
54598	:douta	=	16'h	9369;
54599	:douta	=	16'h	a42b;
54600	:douta	=	16'h	b4ae;
54601	:douta	=	16'h	9bcb;
54602	:douta	=	16'h	c591;
54603	:douta	=	16'h	cdf2;
54604	:douta	=	16'h	d653;
54605	:douta	=	16'h	d674;
54606	:douta	=	16'h	de94;
54607	:douta	=	16'h	de73;
54608	:douta	=	16'h	d674;
54609	:douta	=	16'h	d653;
54610	:douta	=	16'h	cdf1;
54611	:douta	=	16'h	d5d1;
54612	:douta	=	16'h	cd6e;
54613	:douta	=	16'h	c52e;
54614	:douta	=	16'h	c4ec;
54615	:douta	=	16'h	bcab;
54616	:douta	=	16'h	bc49;
54617	:douta	=	16'h	bc28;
54618	:douta	=	16'h	b3e7;
54619	:douta	=	16'h	bbe6;
54620	:douta	=	16'h	bbc5;
54621	:douta	=	16'h	bba5;
54622	:douta	=	16'h	b3a5;
54623	:douta	=	16'h	bba4;
54624	:douta	=	16'h	bbc5;
54625	:douta	=	16'h	bbe5;
54626	:douta	=	16'h	c406;
54627	:douta	=	16'h	c406;
54628	:douta	=	16'h	c426;
54629	:douta	=	16'h	c426;
54630	:douta	=	16'h	c446;
54631	:douta	=	16'h	c447;
54632	:douta	=	16'h	cc48;
54633	:douta	=	16'h	c447;
54634	:douta	=	16'h	cc47;
54635	:douta	=	16'h	cc47;
54636	:douta	=	16'h	cc47;
54637	:douta	=	16'h	cc47;
54638	:douta	=	16'h	cc47;
54639	:douta	=	16'h	cc47;
54640	:douta	=	16'h	cc47;
54641	:douta	=	16'h	cc67;
54642	:douta	=	16'h	cc67;
54643	:douta	=	16'h	cc67;
54644	:douta	=	16'h	cc47;
54645	:douta	=	16'h	cc47;
54646	:douta	=	16'h	cc67;
54647	:douta	=	16'h	cc67;
54648	:douta	=	16'h	cc68;
54649	:douta	=	16'h	cc68;
54650	:douta	=	16'h	cc68;
54651	:douta	=	16'h	cc68;
54652	:douta	=	16'h	cc68;
54653	:douta	=	16'h	cc67;
54654	:douta	=	16'h	cc68;
54655	:douta	=	16'h	cc68;
54656	:douta	=	16'h	cc68;
54657	:douta	=	16'h	cc88;
54658	:douta	=	16'h	cc88;
54659	:douta	=	16'h	cc68;
54660	:douta	=	16'h	cc88;
54661	:douta	=	16'h	cc68;
54662	:douta	=	16'h	cc88;
54663	:douta	=	16'h	cc68;
54664	:douta	=	16'h	cc88;
54665	:douta	=	16'h	cc68;
54666	:douta	=	16'h	cc88;
54667	:douta	=	16'h	cc88;
54668	:douta	=	16'h	cc88;
54669	:douta	=	16'h	d488;
54670	:douta	=	16'h	d488;
54671	:douta	=	16'h	d488;
54672	:douta	=	16'h	cc88;
54673	:douta	=	16'h	cc88;
54674	:douta	=	16'h	cc88;
54675	:douta	=	16'h	d488;
54676	:douta	=	16'h	d4a9;
54677	:douta	=	16'h	cc88;
54678	:douta	=	16'h	d488;
54679	:douta	=	16'h	d489;
54680	:douta	=	16'h	d489;
54681	:douta	=	16'h	d488;
54682	:douta	=	16'h	cc88;
54683	:douta	=	16'h	d4a9;
54684	:douta	=	16'h	cc88;
54685	:douta	=	16'h	d4a9;
54686	:douta	=	16'h	d4a9;
54687	:douta	=	16'h	d489;
54688	:douta	=	16'h	cc88;
54689	:douta	=	16'h	cc88;
54690	:douta	=	16'h	d487;
54691	:douta	=	16'h	ad31;
54692	:douta	=	16'h	deb7;
54693	:douta	=	16'h	cc25;
54694	:douta	=	16'h	d488;
54695	:douta	=	16'h	cc88;
54696	:douta	=	16'h	cc88;
54697	:douta	=	16'h	cc88;
54698	:douta	=	16'h	cc88;
54699	:douta	=	16'h	cc88;
54700	:douta	=	16'h	cc68;
54701	:douta	=	16'h	cc88;
54702	:douta	=	16'h	cc88;
54703	:douta	=	16'h	cc68;
54704	:douta	=	16'h	cc89;
54705	:douta	=	16'h	cc69;
54706	:douta	=	16'h	8bef;
54707	:douta	=	16'h	9c4f;
54708	:douta	=	16'h	9c4f;
54709	:douta	=	16'h	a4b1;
54710	:douta	=	16'h	bd32;
54711	:douta	=	16'h	b533;
54712	:douta	=	16'h	bd33;
54713	:douta	=	16'h	c574;
54714	:douta	=	16'h	bd34;
54715	:douta	=	16'h	b534;
54716	:douta	=	16'h	b514;
54717	:douta	=	16'h	a4b3;
54718	:douta	=	16'h	9493;
54719	:douta	=	16'h	8c73;
54720	:douta	=	16'h	8c53;
54721	:douta	=	16'h	9453;
54722	:douta	=	16'h	9453;
54723	:douta	=	16'h	8c53;
54724	:douta	=	16'h	73d0;
54725	:douta	=	16'h	6b2f;
54726	:douta	=	16'h	6b2e;
54727	:douta	=	16'h	6b4f;
54728	:douta	=	16'h	6b2e;
54729	:douta	=	16'h	6b2e;
54730	:douta	=	16'h	632e;
54731	:douta	=	16'h	5acd;
54732	:douta	=	16'h	6b2e;
54733	:douta	=	16'h	630d;
54734	:douta	=	16'h	62ed;
54735	:douta	=	16'h	736f;
54736	:douta	=	16'h	62cd;
54737	:douta	=	16'h	5a8c;
54738	:douta	=	16'h	5a8b;
54739	:douta	=	16'h	522a;
54740	:douta	=	16'h	62cc;
54741	:douta	=	16'h	7b8f;
54742	:douta	=	16'h	8bf1;
54743	:douta	=	16'h	a4b3;
54744	:douta	=	16'h	9c72;
54745	:douta	=	16'h	83d1;
54746	:douta	=	16'h	6b6f;
54747	:douta	=	16'h	7390;
54748	:douta	=	16'h	6b4f;
54749	:douta	=	16'h	736f;
54750	:douta	=	16'h	6b2f;
54751	:douta	=	16'h	5aee;
54752	:douta	=	16'h	52cd;
54753	:douta	=	16'h	7c73;
54754	:douta	=	16'h	b69a;
54755	:douta	=	16'h	ffff;
54756	:douta	=	16'h	ffff;
54757	:douta	=	16'h	ffff;
54758	:douta	=	16'h	edd5;
54759	:douta	=	16'h	dcd0;
54760	:douta	=	16'h	b346;
54761	:douta	=	16'h	9aa3;
54762	:douta	=	16'h	a305;
54763	:douta	=	16'h	9b67;
54764	:douta	=	16'h	a388;
54765	:douta	=	16'h	a368;
54766	:douta	=	16'h	a368;
54767	:douta	=	16'h	a367;
54768	:douta	=	16'h	a368;
54769	:douta	=	16'h	a368;
54770	:douta	=	16'h	a368;
54771	:douta	=	16'h	a368;
54772	:douta	=	16'h	a368;
54773	:douta	=	16'h	a388;
54774	:douta	=	16'h	a368;
54775	:douta	=	16'h	a368;
54776	:douta	=	16'h	a368;
54777	:douta	=	16'h	a368;
54778	:douta	=	16'h	a368;
54779	:douta	=	16'h	a368;
54780	:douta	=	16'h	a349;
54781	:douta	=	16'h	a348;
54782	:douta	=	16'h	a349;
54783	:douta	=	16'h	a349;
54784	:douta	=	16'h	cdb5;
54785	:douta	=	16'h	bd95;
54786	:douta	=	16'h	ad15;
54787	:douta	=	16'h	9473;
54788	:douta	=	16'h	a515;
54789	:douta	=	16'h	acf5;
54790	:douta	=	16'h	a4d5;
54791	:douta	=	16'h	a4f5;
54792	:douta	=	16'h	94d5;
54793	:douta	=	16'h	9d58;
54794	:douta	=	16'h	6370;
54795	:douta	=	16'h	39e8;
54796	:douta	=	16'h	3166;
54797	:douta	=	16'h	20a3;
54798	:douta	=	16'h	20a2;
54799	:douta	=	16'h	28e3;
54800	:douta	=	16'h	28e3;
54801	:douta	=	16'h	20e3;
54802	:douta	=	16'h	20e3;
54803	:douta	=	16'h	20e3;
54804	:douta	=	16'h	20e3;
54805	:douta	=	16'h	20c3;
54806	:douta	=	16'h	20e3;
54807	:douta	=	16'h	20c3;
54808	:douta	=	16'h	20a2;
54809	:douta	=	16'h	18a2;
54810	:douta	=	16'h	20a2;
54811	:douta	=	16'h	20a2;
54812	:douta	=	16'h	20c2;
54813	:douta	=	16'h	20a2;
54814	:douta	=	16'h	20a2;
54815	:douta	=	16'h	20a2;
54816	:douta	=	16'h	20a2;
54817	:douta	=	16'h	28e3;
54818	:douta	=	16'h	28e3;
54819	:douta	=	16'h	28e3;
54820	:douta	=	16'h	28e2;
54821	:douta	=	16'h	3103;
54822	:douta	=	16'h	3103;
54823	:douta	=	16'h	3123;
54824	:douta	=	16'h	3923;
54825	:douta	=	16'h	3944;
54826	:douta	=	16'h	3923;
54827	:douta	=	16'h	4143;
54828	:douta	=	16'h	49e8;
54829	:douta	=	16'h	4a4a;
54830	:douta	=	16'h	10a5;
54831	:douta	=	16'h	3924;
54832	:douta	=	16'h	59a4;
54833	:douta	=	16'h	59c4;
54834	:douta	=	16'h	59c4;
54835	:douta	=	16'h	59c4;
54836	:douta	=	16'h	61c4;
54837	:douta	=	16'h	61c4;
54838	:douta	=	16'h	61c4;
54839	:douta	=	16'h	61c3;
54840	:douta	=	16'h	69c3;
54841	:douta	=	16'h	69c3;
54842	:douta	=	16'h	6a03;
54843	:douta	=	16'h	7223;
54844	:douta	=	16'h	7244;
54845	:douta	=	16'h	7aa6;
54846	:douta	=	16'h	82e7;
54847	:douta	=	16'h	8b49;
54848	:douta	=	16'h	9beb;
54849	:douta	=	16'h	9c2c;
54850	:douta	=	16'h	b4ce;
54851	:douta	=	16'h	b50f;
54852	:douta	=	16'h	c5b1;
54853	:douta	=	16'h	ce13;
54854	:douta	=	16'h	d633;
54855	:douta	=	16'h	d653;
54856	:douta	=	16'h	e6f5;
54857	:douta	=	16'h	93cb;
54858	:douta	=	16'h	cdf2;
54859	:douta	=	16'h	c5b1;
54860	:douta	=	16'h	bd4f;
54861	:douta	=	16'h	bd0f;
54862	:douta	=	16'h	b4ad;
54863	:douta	=	16'h	a40a;
54864	:douta	=	16'h	a3ca;
54865	:douta	=	16'h	9ba8;
54866	:douta	=	16'h	a387;
54867	:douta	=	16'h	a386;
54868	:douta	=	16'h	a345;
54869	:douta	=	16'h	ab45;
54870	:douta	=	16'h	ab65;
54871	:douta	=	16'h	ab65;
54872	:douta	=	16'h	b385;
54873	:douta	=	16'h	b3a5;
54874	:douta	=	16'h	b3a6;
54875	:douta	=	16'h	bbe6;
54876	:douta	=	16'h	bbe6;
54877	:douta	=	16'h	bbe7;
54878	:douta	=	16'h	bbe7;
54879	:douta	=	16'h	bc07;
54880	:douta	=	16'h	c407;
54881	:douta	=	16'h	c427;
54882	:douta	=	16'h	c426;
54883	:douta	=	16'h	c426;
54884	:douta	=	16'h	c428;
54885	:douta	=	16'h	c426;
54886	:douta	=	16'h	c447;
54887	:douta	=	16'h	c447;
54888	:douta	=	16'h	c447;
54889	:douta	=	16'h	c447;
54890	:douta	=	16'h	c447;
54891	:douta	=	16'h	c447;
54892	:douta	=	16'h	cc67;
54893	:douta	=	16'h	cc67;
54894	:douta	=	16'h	cc47;
54895	:douta	=	16'h	cc47;
54896	:douta	=	16'h	cc47;
54897	:douta	=	16'h	cc68;
54898	:douta	=	16'h	cc48;
54899	:douta	=	16'h	cc67;
54900	:douta	=	16'h	cc67;
54901	:douta	=	16'h	cc67;
54902	:douta	=	16'h	cc67;
54903	:douta	=	16'h	cc67;
54904	:douta	=	16'h	cc68;
54905	:douta	=	16'h	cc68;
54906	:douta	=	16'h	cc68;
54907	:douta	=	16'h	cc68;
54908	:douta	=	16'h	cc68;
54909	:douta	=	16'h	cc68;
54910	:douta	=	16'h	cc68;
54911	:douta	=	16'h	cc67;
54912	:douta	=	16'h	cc68;
54913	:douta	=	16'h	cc68;
54914	:douta	=	16'h	cc68;
54915	:douta	=	16'h	cc68;
54916	:douta	=	16'h	cc68;
54917	:douta	=	16'h	cc88;
54918	:douta	=	16'h	d488;
54919	:douta	=	16'h	cc68;
54920	:douta	=	16'h	cc88;
54921	:douta	=	16'h	cc68;
54922	:douta	=	16'h	cc88;
54923	:douta	=	16'h	cc88;
54924	:douta	=	16'h	cc68;
54925	:douta	=	16'h	cc88;
54926	:douta	=	16'h	cc88;
54927	:douta	=	16'h	d488;
54928	:douta	=	16'h	d489;
54929	:douta	=	16'h	cc88;
54930	:douta	=	16'h	cc88;
54931	:douta	=	16'h	d488;
54932	:douta	=	16'h	cc88;
54933	:douta	=	16'h	d4a9;
54934	:douta	=	16'h	d489;
54935	:douta	=	16'h	d489;
54936	:douta	=	16'h	d488;
54937	:douta	=	16'h	d4a9;
54938	:douta	=	16'h	d4a9;
54939	:douta	=	16'h	d4a9;
54940	:douta	=	16'h	d488;
54941	:douta	=	16'h	d4a9;
54942	:douta	=	16'h	cc88;
54943	:douta	=	16'h	cc88;
54944	:douta	=	16'h	cc88;
54945	:douta	=	16'h	cc88;
54946	:douta	=	16'h	d487;
54947	:douta	=	16'h	ad32;
54948	:douta	=	16'h	deb7;
54949	:douta	=	16'h	cc25;
54950	:douta	=	16'h	cc88;
54951	:douta	=	16'h	cc88;
54952	:douta	=	16'h	cc88;
54953	:douta	=	16'h	cc88;
54954	:douta	=	16'h	d489;
54955	:douta	=	16'h	cc89;
54956	:douta	=	16'h	cc88;
54957	:douta	=	16'h	cc88;
54958	:douta	=	16'h	cc88;
54959	:douta	=	16'h	cc88;
54960	:douta	=	16'h	cc69;
54961	:douta	=	16'h	d487;
54962	:douta	=	16'h	9430;
54963	:douta	=	16'h	940f;
54964	:douta	=	16'h	9c50;
54965	:douta	=	16'h	a491;
54966	:douta	=	16'h	b513;
54967	:douta	=	16'h	b533;
54968	:douta	=	16'h	acf3;
54969	:douta	=	16'h	bd34;
54970	:douta	=	16'h	b513;
54971	:douta	=	16'h	acd4;
54972	:douta	=	16'h	9c93;
54973	:douta	=	16'h	9473;
54974	:douta	=	16'h	8c53;
54975	:douta	=	16'h	8412;
54976	:douta	=	16'h	8432;
54977	:douta	=	16'h	7bd1;
54978	:douta	=	16'h	7bf2;
54979	:douta	=	16'h	8412;
54980	:douta	=	16'h	8433;
54981	:douta	=	16'h	6b4f;
54982	:douta	=	16'h	630e;
54983	:douta	=	16'h	6b2e;
54984	:douta	=	16'h	62ed;
54985	:douta	=	16'h	62ed;
54986	:douta	=	16'h	630d;
54987	:douta	=	16'h	62cd;
54988	:douta	=	16'h	62ed;
54989	:douta	=	16'h	7b6f;
54990	:douta	=	16'h	630e;
54991	:douta	=	16'h	62ed;
54992	:douta	=	16'h	62ed;
54993	:douta	=	16'h	62ed;
54994	:douta	=	16'h	7b8f;
54995	:douta	=	16'h	83d0;
54996	:douta	=	16'h	9c92;
54997	:douta	=	16'h	9452;
54998	:douta	=	16'h	a493;
54999	:douta	=	16'h	838f;
55000	:douta	=	16'h	734e;
55001	:douta	=	16'h	62ed;
55002	:douta	=	16'h	83f0;
55003	:douta	=	16'h	6b4f;
55004	:douta	=	16'h	4a2a;
55005	:douta	=	16'h	5acd;
55006	:douta	=	16'h	8473;
55007	:douta	=	16'h	ae18;
55008	:douta	=	16'h	c73d;
55009	:douta	=	16'h	ffff;
55010	:douta	=	16'h	ffff;
55011	:douta	=	16'h	f636;
55012	:douta	=	16'h	d44d;
55013	:douta	=	16'h	c389;
55014	:douta	=	16'h	aac4;
55015	:douta	=	16'h	9ac4;
55016	:douta	=	16'h	a388;
55017	:douta	=	16'h	a388;
55018	:douta	=	16'h	a388;
55019	:douta	=	16'h	ab88;
55020	:douta	=	16'h	a388;
55021	:douta	=	16'h	a388;
55022	:douta	=	16'h	a368;
55023	:douta	=	16'h	ab88;
55024	:douta	=	16'h	a368;
55025	:douta	=	16'h	a368;
55026	:douta	=	16'h	a368;
55027	:douta	=	16'h	ab88;
55028	:douta	=	16'h	ab68;
55029	:douta	=	16'h	a368;
55030	:douta	=	16'h	a368;
55031	:douta	=	16'h	a368;
55032	:douta	=	16'h	a368;
55033	:douta	=	16'h	a388;
55034	:douta	=	16'h	a368;
55035	:douta	=	16'h	a368;
55036	:douta	=	16'h	a368;
55037	:douta	=	16'h	a368;
55038	:douta	=	16'h	a368;
55039	:douta	=	16'h	a369;
55040	:douta	=	16'h	c5b6;
55041	:douta	=	16'h	ad56;
55042	:douta	=	16'h	9494;
55043	:douta	=	16'h	a515;
55044	:douta	=	16'h	a4f5;
55045	:douta	=	16'h	ad16;
55046	:douta	=	16'h	a4f5;
55047	:douta	=	16'h	a4f5;
55048	:douta	=	16'h	8475;
55049	:douta	=	16'h	634e;
55050	:douta	=	16'h	1020;
55051	:douta	=	16'h	3125;
55052	:douta	=	16'h	31a6;
55053	:douta	=	16'h	426c;
55054	:douta	=	16'h	4aac;
55055	:douta	=	16'h	424b;
55056	:douta	=	16'h	3165;
55057	:douta	=	16'h	28e3;
55058	:douta	=	16'h	2082;
55059	:douta	=	16'h	28c3;
55060	:douta	=	16'h	20c3;
55061	:douta	=	16'h	20e3;
55062	:douta	=	16'h	20c3;
55063	:douta	=	16'h	20e3;
55064	:douta	=	16'h	1882;
55065	:douta	=	16'h	20a2;
55066	:douta	=	16'h	20a2;
55067	:douta	=	16'h	20a2;
55068	:douta	=	16'h	20c2;
55069	:douta	=	16'h	20c2;
55070	:douta	=	16'h	20a2;
55071	:douta	=	16'h	20a2;
55072	:douta	=	16'h	20c2;
55073	:douta	=	16'h	28e3;
55074	:douta	=	16'h	28e3;
55075	:douta	=	16'h	28e2;
55076	:douta	=	16'h	28e2;
55077	:douta	=	16'h	28e2;
55078	:douta	=	16'h	30e2;
55079	:douta	=	16'h	3103;
55080	:douta	=	16'h	30e2;
55081	:douta	=	16'h	30c2;
55082	:douta	=	16'h	3902;
55083	:douta	=	16'h	3902;
55084	:douta	=	16'h	4a4a;
55085	:douta	=	16'h	39e9;
55086	:douta	=	16'h	18c4;
55087	:douta	=	16'h	51c5;
55088	:douta	=	16'h	6246;
55089	:douta	=	16'h	6ac8;
55090	:douta	=	16'h	7329;
55091	:douta	=	16'h	838b;
55092	:douta	=	16'h	8bcc;
55093	:douta	=	16'h	9c6e;
55094	:douta	=	16'h	acef;
55095	:douta	=	16'h	ad30;
55096	:douta	=	16'h	bdb2;
55097	:douta	=	16'h	bd92;
55098	:douta	=	16'h	d675;
55099	:douta	=	16'h	bd71;
55100	:douta	=	16'h	bd51;
55101	:douta	=	16'h	b50f;
55102	:douta	=	16'h	accd;
55103	:douta	=	16'h	a44c;
55104	:douta	=	16'h	9bca;
55105	:douta	=	16'h	9389;
55106	:douta	=	16'h	8b27;
55107	:douta	=	16'h	8b07;
55108	:douta	=	16'h	8ae6;
55109	:douta	=	16'h	8aa5;
55110	:douta	=	16'h	8285;
55111	:douta	=	16'h	8285;
55112	:douta	=	16'h	8aa5;
55113	:douta	=	16'h	51c5;
55114	:douta	=	16'h	92e5;
55115	:douta	=	16'h	92c5;
55116	:douta	=	16'h	9306;
55117	:douta	=	16'h	9305;
55118	:douta	=	16'h	9305;
55119	:douta	=	16'h	9306;
55120	:douta	=	16'h	9b27;
55121	:douta	=	16'h	9326;
55122	:douta	=	16'h	a366;
55123	:douta	=	16'h	ab86;
55124	:douta	=	16'h	aba7;
55125	:douta	=	16'h	aba6;
55126	:douta	=	16'h	b3c7;
55127	:douta	=	16'h	b3c7;
55128	:douta	=	16'h	bbc7;
55129	:douta	=	16'h	bbe7;
55130	:douta	=	16'h	bbe6;
55131	:douta	=	16'h	bbe7;
55132	:douta	=	16'h	c3e7;
55133	:douta	=	16'h	bbe7;
55134	:douta	=	16'h	bc07;
55135	:douta	=	16'h	bc06;
55136	:douta	=	16'h	c427;
55137	:douta	=	16'h	c407;
55138	:douta	=	16'h	c426;
55139	:douta	=	16'h	c447;
55140	:douta	=	16'h	c426;
55141	:douta	=	16'h	c447;
55142	:douta	=	16'h	c447;
55143	:douta	=	16'h	c448;
55144	:douta	=	16'h	c448;
55145	:douta	=	16'h	cc47;
55146	:douta	=	16'h	cc47;
55147	:douta	=	16'h	cc47;
55148	:douta	=	16'h	cc47;
55149	:douta	=	16'h	cc47;
55150	:douta	=	16'h	cc67;
55151	:douta	=	16'h	cc67;
55152	:douta	=	16'h	cc47;
55153	:douta	=	16'h	cc47;
55154	:douta	=	16'h	cc68;
55155	:douta	=	16'h	cc48;
55156	:douta	=	16'h	cc68;
55157	:douta	=	16'h	cc68;
55158	:douta	=	16'h	cc48;
55159	:douta	=	16'h	cc48;
55160	:douta	=	16'h	cc68;
55161	:douta	=	16'h	cc68;
55162	:douta	=	16'h	cc68;
55163	:douta	=	16'h	cc68;
55164	:douta	=	16'h	cc68;
55165	:douta	=	16'h	cc68;
55166	:douta	=	16'h	cc68;
55167	:douta	=	16'h	cc68;
55168	:douta	=	16'h	cc68;
55169	:douta	=	16'h	cc68;
55170	:douta	=	16'h	cc68;
55171	:douta	=	16'h	cc68;
55172	:douta	=	16'h	cc68;
55173	:douta	=	16'h	cc68;
55174	:douta	=	16'h	cc68;
55175	:douta	=	16'h	cc68;
55176	:douta	=	16'h	d488;
55177	:douta	=	16'h	cc88;
55178	:douta	=	16'h	d488;
55179	:douta	=	16'h	d488;
55180	:douta	=	16'h	cc88;
55181	:douta	=	16'h	cc68;
55182	:douta	=	16'h	cc69;
55183	:douta	=	16'h	cc88;
55184	:douta	=	16'h	cc88;
55185	:douta	=	16'h	d4a9;
55186	:douta	=	16'h	d4a9;
55187	:douta	=	16'h	d4a9;
55188	:douta	=	16'h	d488;
55189	:douta	=	16'h	cc89;
55190	:douta	=	16'h	d489;
55191	:douta	=	16'h	d489;
55192	:douta	=	16'h	d4a9;
55193	:douta	=	16'h	d488;
55194	:douta	=	16'h	d4a9;
55195	:douta	=	16'h	d488;
55196	:douta	=	16'h	d488;
55197	:douta	=	16'h	cc88;
55198	:douta	=	16'h	d4a9;
55199	:douta	=	16'h	d4a9;
55200	:douta	=	16'h	d488;
55201	:douta	=	16'h	d4a9;
55202	:douta	=	16'h	d488;
55203	:douta	=	16'h	ad32;
55204	:douta	=	16'h	deb7;
55205	:douta	=	16'h	cc25;
55206	:douta	=	16'h	cc88;
55207	:douta	=	16'h	d488;
55208	:douta	=	16'h	cc88;
55209	:douta	=	16'h	cc88;
55210	:douta	=	16'h	cc89;
55211	:douta	=	16'h	cc89;
55212	:douta	=	16'h	cc88;
55213	:douta	=	16'h	cc89;
55214	:douta	=	16'h	cc89;
55215	:douta	=	16'h	cc69;
55216	:douta	=	16'h	cc89;
55217	:douta	=	16'h	d488;
55218	:douta	=	16'h	9c0f;
55219	:douta	=	16'h	8bef;
55220	:douta	=	16'h	9c51;
55221	:douta	=	16'h	a492;
55222	:douta	=	16'h	9452;
55223	:douta	=	16'h	a4d4;
55224	:douta	=	16'h	a4d4;
55225	:douta	=	16'h	9cb3;
55226	:douta	=	16'h	9cb3;
55227	:douta	=	16'h	9452;
55228	:douta	=	16'h	8432;
55229	:douta	=	16'h	8412;
55230	:douta	=	16'h	73b0;
55231	:douta	=	16'h	6b90;
55232	:douta	=	16'h	6b6f;
55233	:douta	=	16'h	6b4f;
55234	:douta	=	16'h	6b70;
55235	:douta	=	16'h	630e;
55236	:douta	=	16'h	630e;
55237	:douta	=	16'h	632e;
55238	:douta	=	16'h	630e;
55239	:douta	=	16'h	630e;
55240	:douta	=	16'h	62cd;
55241	:douta	=	16'h	5aac;
55242	:douta	=	16'h	62cd;
55243	:douta	=	16'h	62ed;
55244	:douta	=	16'h	6b0d;
55245	:douta	=	16'h	83f0;
55246	:douta	=	16'h	8c11;
55247	:douta	=	16'h	8bf1;
55248	:douta	=	16'h	9452;
55249	:douta	=	16'h	8410;
55250	:douta	=	16'h	6b4e;
55251	:douta	=	16'h	7bb0;
55252	:douta	=	16'h	7bb0;
55253	:douta	=	16'h	6acd;
55254	:douta	=	16'h	6acd;
55255	:douta	=	16'h	6b0d;
55256	:douta	=	16'h	6b8f;
55257	:douta	=	16'h	add7;
55258	:douta	=	16'h	efff;
55259	:douta	=	16'h	ffff;
55260	:douta	=	16'h	ffff;
55261	:douta	=	16'h	ffbd;
55262	:douta	=	16'h	ed71;
55263	:douta	=	16'h	bb87;
55264	:douta	=	16'h	b305;
55265	:douta	=	16'h	a304;
55266	:douta	=	16'h	a367;
55267	:douta	=	16'h	aba8;
55268	:douta	=	16'h	aba8;
55269	:douta	=	16'h	aba7;
55270	:douta	=	16'h	a388;
55271	:douta	=	16'h	aba8;
55272	:douta	=	16'h	ab88;
55273	:douta	=	16'h	ab88;
55274	:douta	=	16'h	ab88;
55275	:douta	=	16'h	a388;
55276	:douta	=	16'h	a388;
55277	:douta	=	16'h	ab88;
55278	:douta	=	16'h	ab88;
55279	:douta	=	16'h	ab88;
55280	:douta	=	16'h	ab89;
55281	:douta	=	16'h	ab88;
55282	:douta	=	16'h	ab89;
55283	:douta	=	16'h	a388;
55284	:douta	=	16'h	aba8;
55285	:douta	=	16'h	ab88;
55286	:douta	=	16'h	ab88;
55287	:douta	=	16'h	a368;
55288	:douta	=	16'h	a368;
55289	:douta	=	16'h	a368;
55290	:douta	=	16'h	a368;
55291	:douta	=	16'h	a368;
55292	:douta	=	16'h	a368;
55293	:douta	=	16'h	ab68;
55294	:douta	=	16'h	ab68;
55295	:douta	=	16'h	a368;
55296	:douta	=	16'h	c596;
55297	:douta	=	16'h	a516;
55298	:douta	=	16'h	8c53;
55299	:douta	=	16'h	ad36;
55300	:douta	=	16'h	a4f5;
55301	:douta	=	16'h	ad16;
55302	:douta	=	16'h	a515;
55303	:douta	=	16'h	a4f5;
55304	:douta	=	16'h	8cd6;
55305	:douta	=	16'h	41e8;
55306	:douta	=	16'h	1861;
55307	:douta	=	16'h	20c2;
55308	:douta	=	16'h	28c3;
55309	:douta	=	16'h	3125;
55310	:douta	=	16'h	39c8;
55311	:douta	=	16'h	426b;
55312	:douta	=	16'h	42cd;
55313	:douta	=	16'h	428c;
55314	:douta	=	16'h	3187;
55315	:douta	=	16'h	2082;
55316	:douta	=	16'h	2082;
55317	:douta	=	16'h	20a2;
55318	:douta	=	16'h	20c3;
55319	:douta	=	16'h	20e3;
55320	:douta	=	16'h	2082;
55321	:douta	=	16'h	20a2;
55322	:douta	=	16'h	20a2;
55323	:douta	=	16'h	20a2;
55324	:douta	=	16'h	20a2;
55325	:douta	=	16'h	20a2;
55326	:douta	=	16'h	20a2;
55327	:douta	=	16'h	2082;
55328	:douta	=	16'h	20a2;
55329	:douta	=	16'h	20a2;
55330	:douta	=	16'h	20a1;
55331	:douta	=	16'h	20a1;
55332	:douta	=	16'h	28c2;
55333	:douta	=	16'h	28e2;
55334	:douta	=	16'h	3123;
55335	:douta	=	16'h	4165;
55336	:douta	=	16'h	41a5;
55337	:douta	=	16'h	51e6;
55338	:douta	=	16'h	5227;
55339	:douta	=	16'h	62a9;
55340	:douta	=	16'h	4a29;
55341	:douta	=	16'h	31c8;
55342	:douta	=	16'h	3146;
55343	:douta	=	16'h	942f;
55344	:douta	=	16'h	9c8f;
55345	:douta	=	16'h	9cd0;
55346	:douta	=	16'h	a4f1;
55347	:douta	=	16'h	a4f0;
55348	:douta	=	16'h	acf0;
55349	:douta	=	16'h	a4cf;
55350	:douta	=	16'h	9c8e;
55351	:douta	=	16'h	9c6d;
55352	:douta	=	16'h	940c;
55353	:douta	=	16'h	8bcb;
55354	:douta	=	16'h	b510;
55355	:douta	=	16'h	7aa6;
55356	:douta	=	16'h	7aa6;
55357	:douta	=	16'h	7a65;
55358	:douta	=	16'h	7a64;
55359	:douta	=	16'h	7a44;
55360	:douta	=	16'h	7a44;
55361	:douta	=	16'h	7a44;
55362	:douta	=	16'h	7a64;
55363	:douta	=	16'h	8284;
55364	:douta	=	16'h	8aa5;
55365	:douta	=	16'h	8aa5;
55366	:douta	=	16'h	8ac5;
55367	:douta	=	16'h	8ae6;
55368	:douta	=	16'h	92e6;
55369	:douta	=	16'h	59c4;
55370	:douta	=	16'h	9b27;
55371	:douta	=	16'h	9306;
55372	:douta	=	16'h	9326;
55373	:douta	=	16'h	9326;
55374	:douta	=	16'h	9307;
55375	:douta	=	16'h	9306;
55376	:douta	=	16'h	9b26;
55377	:douta	=	16'h	9b47;
55378	:douta	=	16'h	a367;
55379	:douta	=	16'h	ab86;
55380	:douta	=	16'h	ab87;
55381	:douta	=	16'h	b3a7;
55382	:douta	=	16'h	b3c7;
55383	:douta	=	16'h	b3c7;
55384	:douta	=	16'h	b3c6;
55385	:douta	=	16'h	bbe7;
55386	:douta	=	16'h	bbe6;
55387	:douta	=	16'h	bbe7;
55388	:douta	=	16'h	bc07;
55389	:douta	=	16'h	bc06;
55390	:douta	=	16'h	c406;
55391	:douta	=	16'h	bc06;
55392	:douta	=	16'h	bc07;
55393	:douta	=	16'h	c407;
55394	:douta	=	16'h	c407;
55395	:douta	=	16'h	c427;
55396	:douta	=	16'h	c427;
55397	:douta	=	16'h	c447;
55398	:douta	=	16'h	c447;
55399	:douta	=	16'h	c427;
55400	:douta	=	16'h	c448;
55401	:douta	=	16'h	c448;
55402	:douta	=	16'h	cc47;
55403	:douta	=	16'h	c447;
55404	:douta	=	16'h	c447;
55405	:douta	=	16'h	c447;
55406	:douta	=	16'h	cc47;
55407	:douta	=	16'h	cc47;
55408	:douta	=	16'h	cc47;
55409	:douta	=	16'h	cc47;
55410	:douta	=	16'h	cc47;
55411	:douta	=	16'h	cc68;
55412	:douta	=	16'h	cc67;
55413	:douta	=	16'h	cc68;
55414	:douta	=	16'h	cc68;
55415	:douta	=	16'h	cc68;
55416	:douta	=	16'h	cc48;
55417	:douta	=	16'h	cc48;
55418	:douta	=	16'h	cc47;
55419	:douta	=	16'h	cc88;
55420	:douta	=	16'h	cc68;
55421	:douta	=	16'h	cc68;
55422	:douta	=	16'h	cc68;
55423	:douta	=	16'h	cc68;
55424	:douta	=	16'h	cc68;
55425	:douta	=	16'h	cc68;
55426	:douta	=	16'h	cc68;
55427	:douta	=	16'h	cc68;
55428	:douta	=	16'h	cc68;
55429	:douta	=	16'h	cc68;
55430	:douta	=	16'h	d488;
55431	:douta	=	16'h	cc68;
55432	:douta	=	16'h	cc88;
55433	:douta	=	16'h	cc88;
55434	:douta	=	16'h	cc68;
55435	:douta	=	16'h	cc68;
55436	:douta	=	16'h	cc88;
55437	:douta	=	16'h	d489;
55438	:douta	=	16'h	d489;
55439	:douta	=	16'h	cc88;
55440	:douta	=	16'h	cc88;
55441	:douta	=	16'h	cc88;
55442	:douta	=	16'h	cc88;
55443	:douta	=	16'h	d488;
55444	:douta	=	16'h	cc88;
55445	:douta	=	16'h	cc88;
55446	:douta	=	16'h	d489;
55447	:douta	=	16'h	d489;
55448	:douta	=	16'h	d4a9;
55449	:douta	=	16'h	d488;
55450	:douta	=	16'h	cc88;
55451	:douta	=	16'h	cc88;
55452	:douta	=	16'h	d4a9;
55453	:douta	=	16'h	cc88;
55454	:douta	=	16'h	d488;
55455	:douta	=	16'h	d488;
55456	:douta	=	16'h	cc88;
55457	:douta	=	16'h	cc88;
55458	:douta	=	16'h	d488;
55459	:douta	=	16'h	ad32;
55460	:douta	=	16'h	deb8;
55461	:douta	=	16'h	cc25;
55462	:douta	=	16'h	cc88;
55463	:douta	=	16'h	cc89;
55464	:douta	=	16'h	cc88;
55465	:douta	=	16'h	cc88;
55466	:douta	=	16'h	cc89;
55467	:douta	=	16'h	cc89;
55468	:douta	=	16'h	cc88;
55469	:douta	=	16'h	cc69;
55470	:douta	=	16'h	cc89;
55471	:douta	=	16'h	cc69;
55472	:douta	=	16'h	cc69;
55473	:douta	=	16'h	cc69;
55474	:douta	=	16'h	a42d;
55475	:douta	=	16'h	83f0;
55476	:douta	=	16'h	9431;
55477	:douta	=	16'h	9451;
55478	:douta	=	16'h	9c73;
55479	:douta	=	16'h	9452;
55480	:douta	=	16'h	8c73;
55481	:douta	=	16'h	8412;
55482	:douta	=	16'h	8c53;
55483	:douta	=	16'h	7bf2;
55484	:douta	=	16'h	7bd1;
55485	:douta	=	16'h	73b0;
55486	:douta	=	16'h	6b6f;
55487	:douta	=	16'h	6b2e;
55488	:douta	=	16'h	6b4f;
55489	:douta	=	16'h	632e;
55490	:douta	=	16'h	6b4f;
55491	:douta	=	16'h	6b4f;
55492	:douta	=	16'h	5acd;
55493	:douta	=	16'h	6b4f;
55494	:douta	=	16'h	5aee;
55495	:douta	=	16'h	62ad;
55496	:douta	=	16'h	62cd;
55497	:douta	=	16'h	62ed;
55498	:douta	=	16'h	8c32;
55499	:douta	=	16'h	7bd0;
55500	:douta	=	16'h	8c11;
55501	:douta	=	16'h	9c72;
55502	:douta	=	16'h	9c72;
55503	:douta	=	16'h	422a;
55504	:douta	=	16'h	9432;
55505	:douta	=	16'h	7b6e;
55506	:douta	=	16'h	62ad;
55507	:douta	=	16'h	5aad;
55508	:douta	=	16'h	73b0;
55509	:douta	=	16'h	73f0;
55510	:douta	=	16'h	8c93;
55511	:douta	=	16'h	c71c;
55512	:douta	=	16'h	efff;
55513	:douta	=	16'h	ffff;
55514	:douta	=	16'h	ff1a;
55515	:douta	=	16'h	f5d4;
55516	:douta	=	16'h	cbca;
55517	:douta	=	16'h	bb47;
55518	:douta	=	16'h	a2e3;
55519	:douta	=	16'h	a3a7;
55520	:douta	=	16'h	abc8;
55521	:douta	=	16'h	b3a9;
55522	:douta	=	16'h	aba8;
55523	:douta	=	16'h	b3a8;
55524	:douta	=	16'h	b3c8;
55525	:douta	=	16'h	ab89;
55526	:douta	=	16'h	aba8;
55527	:douta	=	16'h	ab88;
55528	:douta	=	16'h	ab88;
55529	:douta	=	16'h	aba8;
55530	:douta	=	16'h	ab89;
55531	:douta	=	16'h	ab88;
55532	:douta	=	16'h	b3a8;
55533	:douta	=	16'h	ab88;
55534	:douta	=	16'h	aba9;
55535	:douta	=	16'h	ab89;
55536	:douta	=	16'h	aba8;
55537	:douta	=	16'h	ab89;
55538	:douta	=	16'h	ab88;
55539	:douta	=	16'h	ab88;
55540	:douta	=	16'h	ab88;
55541	:douta	=	16'h	ab88;
55542	:douta	=	16'h	ab88;
55543	:douta	=	16'h	ab88;
55544	:douta	=	16'h	ab89;
55545	:douta	=	16'h	ab88;
55546	:douta	=	16'h	a368;
55547	:douta	=	16'h	a368;
55548	:douta	=	16'h	a368;
55549	:douta	=	16'h	ab68;
55550	:douta	=	16'h	ab68;
55551	:douta	=	16'h	a368;
55552	:douta	=	16'h	b556;
55553	:douta	=	16'h	9494;
55554	:douta	=	16'h	8412;
55555	:douta	=	16'h	ad36;
55556	:douta	=	16'h	ad36;
55557	:douta	=	16'h	ad15;
55558	:douta	=	16'h	a515;
55559	:douta	=	16'h	94b5;
55560	:douta	=	16'h	a579;
55561	:douta	=	16'h	1040;
55562	:douta	=	16'h	28e3;
55563	:douta	=	16'h	28e3;
55564	:douta	=	16'h	28e3;
55565	:douta	=	16'h	28e3;
55566	:douta	=	16'h	28e3;
55567	:douta	=	16'h	28e3;
55568	:douta	=	16'h	20c2;
55569	:douta	=	16'h	20c2;
55570	:douta	=	16'h	31a7;
55571	:douta	=	16'h	428c;
55572	:douta	=	16'h	4acd;
55573	:douta	=	16'h	428c;
55574	:douta	=	16'h	3a2a;
55575	:douta	=	16'h	2925;
55576	:douta	=	16'h	2924;
55577	:douta	=	16'h	2945;
55578	:douta	=	16'h	2965;
55579	:douta	=	16'h	3186;
55580	:douta	=	16'h	3986;
55581	:douta	=	16'h	39a6;
55582	:douta	=	16'h	39c7;
55583	:douta	=	16'h	41e8;
55584	:douta	=	16'h	4a28;
55585	:douta	=	16'h	528a;
55586	:douta	=	16'h	52aa;
55587	:douta	=	16'h	5aaa;
55588	:douta	=	16'h	5aaa;
55589	:douta	=	16'h	5aca;
55590	:douta	=	16'h	62ca;
55591	:douta	=	16'h	62c9;
55592	:douta	=	16'h	6288;
55593	:douta	=	16'h	5a47;
55594	:douta	=	16'h	5a47;
55595	:douta	=	16'h	5226;
55596	:douta	=	16'h	4a4a;
55597	:douta	=	16'h	2167;
55598	:douta	=	16'h	3924;
55599	:douta	=	16'h	59a4;
55600	:douta	=	16'h	5184;
55601	:douta	=	16'h	5184;
55602	:douta	=	16'h	59a4;
55603	:douta	=	16'h	59a4;
55604	:douta	=	16'h	59a3;
55605	:douta	=	16'h	61c4;
55606	:douta	=	16'h	61e4;
55607	:douta	=	16'h	6a04;
55608	:douta	=	16'h	6a04;
55609	:douta	=	16'h	838c;
55610	:douta	=	16'h	8329;
55611	:douta	=	16'h	7a85;
55612	:douta	=	16'h	7a85;
55613	:douta	=	16'h	82a5;
55614	:douta	=	16'h	7a85;
55615	:douta	=	16'h	82a5;
55616	:douta	=	16'h	82a5;
55617	:douta	=	16'h	82c5;
55618	:douta	=	16'h	82c5;
55619	:douta	=	16'h	8aa5;
55620	:douta	=	16'h	8aa5;
55621	:douta	=	16'h	8ac6;
55622	:douta	=	16'h	8ac6;
55623	:douta	=	16'h	8ac6;
55624	:douta	=	16'h	92e6;
55625	:douta	=	16'h	59e5;
55626	:douta	=	16'h	9b47;
55627	:douta	=	16'h	9326;
55628	:douta	=	16'h	9326;
55629	:douta	=	16'h	9326;
55630	:douta	=	16'h	9326;
55631	:douta	=	16'h	9326;
55632	:douta	=	16'h	9306;
55633	:douta	=	16'h	9b26;
55634	:douta	=	16'h	a367;
55635	:douta	=	16'h	ab86;
55636	:douta	=	16'h	ab87;
55637	:douta	=	16'h	b3a7;
55638	:douta	=	16'h	b3c7;
55639	:douta	=	16'h	b3c7;
55640	:douta	=	16'h	b3e6;
55641	:douta	=	16'h	b3e6;
55642	:douta	=	16'h	bbc6;
55643	:douta	=	16'h	bbe6;
55644	:douta	=	16'h	bbe7;
55645	:douta	=	16'h	bbe7;
55646	:douta	=	16'h	bc07;
55647	:douta	=	16'h	c407;
55648	:douta	=	16'h	c407;
55649	:douta	=	16'h	c407;
55650	:douta	=	16'h	c427;
55651	:douta	=	16'h	c426;
55652	:douta	=	16'h	c427;
55653	:douta	=	16'h	c426;
55654	:douta	=	16'h	c426;
55655	:douta	=	16'h	c448;
55656	:douta	=	16'h	c428;
55657	:douta	=	16'h	c448;
55658	:douta	=	16'h	cc47;
55659	:douta	=	16'h	c447;
55660	:douta	=	16'h	cc47;
55661	:douta	=	16'h	cc47;
55662	:douta	=	16'h	cc68;
55663	:douta	=	16'h	cc47;
55664	:douta	=	16'h	cc47;
55665	:douta	=	16'h	cc47;
55666	:douta	=	16'h	cc67;
55667	:douta	=	16'h	cc48;
55668	:douta	=	16'h	cc68;
55669	:douta	=	16'h	cc68;
55670	:douta	=	16'h	cc68;
55671	:douta	=	16'h	cc68;
55672	:douta	=	16'h	cc68;
55673	:douta	=	16'h	cc68;
55674	:douta	=	16'h	cc68;
55675	:douta	=	16'h	cc48;
55676	:douta	=	16'h	cc68;
55677	:douta	=	16'h	cc68;
55678	:douta	=	16'h	cc68;
55679	:douta	=	16'h	cc68;
55680	:douta	=	16'h	cc68;
55681	:douta	=	16'h	cc68;
55682	:douta	=	16'h	cc88;
55683	:douta	=	16'h	cc68;
55684	:douta	=	16'h	cc68;
55685	:douta	=	16'h	cc88;
55686	:douta	=	16'h	cc68;
55687	:douta	=	16'h	cc88;
55688	:douta	=	16'h	cc88;
55689	:douta	=	16'h	cc68;
55690	:douta	=	16'h	cc88;
55691	:douta	=	16'h	cc88;
55692	:douta	=	16'h	cc88;
55693	:douta	=	16'h	d4a9;
55694	:douta	=	16'h	cc88;
55695	:douta	=	16'h	d4a9;
55696	:douta	=	16'h	d4a9;
55697	:douta	=	16'h	cc88;
55698	:douta	=	16'h	cc88;
55699	:douta	=	16'h	d488;
55700	:douta	=	16'h	cc89;
55701	:douta	=	16'h	d489;
55702	:douta	=	16'h	d489;
55703	:douta	=	16'h	cc89;
55704	:douta	=	16'h	cc89;
55705	:douta	=	16'h	d489;
55706	:douta	=	16'h	d488;
55707	:douta	=	16'h	d488;
55708	:douta	=	16'h	d4a9;
55709	:douta	=	16'h	cc88;
55710	:douta	=	16'h	d488;
55711	:douta	=	16'h	cc88;
55712	:douta	=	16'h	d4a9;
55713	:douta	=	16'h	cc89;
55714	:douta	=	16'h	d487;
55715	:douta	=	16'h	ad33;
55716	:douta	=	16'h	deb7;
55717	:douta	=	16'h	cc26;
55718	:douta	=	16'h	d488;
55719	:douta	=	16'h	cc89;
55720	:douta	=	16'h	cc89;
55721	:douta	=	16'h	cc88;
55722	:douta	=	16'h	cc89;
55723	:douta	=	16'h	cc69;
55724	:douta	=	16'h	d489;
55725	:douta	=	16'h	cc69;
55726	:douta	=	16'h	cc69;
55727	:douta	=	16'h	cc69;
55728	:douta	=	16'h	cc69;
55729	:douta	=	16'h	cc69;
55730	:douta	=	16'h	cc69;
55731	:douta	=	16'h	9c50;
55732	:douta	=	16'h	9451;
55733	:douta	=	16'h	9451;
55734	:douta	=	16'h	83f1;
55735	:douta	=	16'h	8c12;
55736	:douta	=	16'h	7bb0;
55737	:douta	=	16'h	7bd1;
55738	:douta	=	16'h	73b0;
55739	:douta	=	16'h	8432;
55740	:douta	=	16'h	632e;
55741	:douta	=	16'h	632e;
55742	:douta	=	16'h	6b2e;
55743	:douta	=	16'h	6b0e;
55744	:douta	=	16'h	62cd;
55745	:douta	=	16'h	5aab;
55746	:douta	=	16'h	528b;
55747	:douta	=	16'h	5aed;
55748	:douta	=	16'h	630e;
55749	:douta	=	16'h	83f1;
55750	:douta	=	16'h	9472;
55751	:douta	=	16'h	9472;
55752	:douta	=	16'h	6b0e;
55753	:douta	=	16'h	9432;
55754	:douta	=	16'h	7bb0;
55755	:douta	=	16'h	730e;
55756	:douta	=	16'h	6acc;
55757	:douta	=	16'h	7b8f;
55758	:douta	=	16'h	83ef;
55759	:douta	=	16'h	9d14;
55760	:douta	=	16'h	df5c;
55761	:douta	=	16'h	f7ff;
55762	:douta	=	16'h	ffff;
55763	:douta	=	16'h	ffff;
55764	:douta	=	16'h	ffff;
55765	:douta	=	16'h	fe15;
55766	:douta	=	16'h	e50f;
55767	:douta	=	16'h	bb46;
55768	:douta	=	16'h	b304;
55769	:douta	=	16'h	ab66;
55770	:douta	=	16'h	b3c8;
55771	:douta	=	16'h	b3c8;
55772	:douta	=	16'h	b3c8;
55773	:douta	=	16'h	b3a8;
55774	:douta	=	16'h	b3c8;
55775	:douta	=	16'h	b3c8;
55776	:douta	=	16'h	abc8;
55777	:douta	=	16'h	b3a8;
55778	:douta	=	16'h	b3a8;
55779	:douta	=	16'h	b3a8;
55780	:douta	=	16'h	aba8;
55781	:douta	=	16'h	aba8;
55782	:douta	=	16'h	b3a8;
55783	:douta	=	16'h	b3c8;
55784	:douta	=	16'h	b3a8;
55785	:douta	=	16'h	ab88;
55786	:douta	=	16'h	aba8;
55787	:douta	=	16'h	b3c8;
55788	:douta	=	16'h	aba8;
55789	:douta	=	16'h	b3a8;
55790	:douta	=	16'h	aba8;
55791	:douta	=	16'h	aba8;
55792	:douta	=	16'h	ab88;
55793	:douta	=	16'h	ab88;
55794	:douta	=	16'h	aba9;
55795	:douta	=	16'h	ab89;
55796	:douta	=	16'h	ab88;
55797	:douta	=	16'h	aba9;
55798	:douta	=	16'h	aba9;
55799	:douta	=	16'h	ab88;
55800	:douta	=	16'h	ab89;
55801	:douta	=	16'h	ab88;
55802	:douta	=	16'h	a368;
55803	:douta	=	16'h	ab68;
55804	:douta	=	16'h	ab68;
55805	:douta	=	16'h	a368;
55806	:douta	=	16'h	ab88;
55807	:douta	=	16'h	a368;
55808	:douta	=	16'h	b536;
55809	:douta	=	16'h	8c73;
55810	:douta	=	16'h	8c53;
55811	:douta	=	16'h	a4f5;
55812	:douta	=	16'h	ad36;
55813	:douta	=	16'h	a4f5;
55814	:douta	=	16'h	9cf5;
55815	:douta	=	16'h	8c95;
55816	:douta	=	16'h	8cf7;
55817	:douta	=	16'h	1861;
55818	:douta	=	16'h	28e3;
55819	:douta	=	16'h	2903;
55820	:douta	=	16'h	28e3;
55821	:douta	=	16'h	28e3;
55822	:douta	=	16'h	28e3;
55823	:douta	=	16'h	2903;
55824	:douta	=	16'h	20c3;
55825	:douta	=	16'h	28e3;
55826	:douta	=	16'h	20a2;
55827	:douta	=	16'h	2924;
55828	:douta	=	16'h	2966;
55829	:douta	=	16'h	426b;
55830	:douta	=	16'h	4aac;
55831	:douta	=	16'h	31a8;
55832	:douta	=	16'h	39c8;
55833	:douta	=	16'h	39e8;
55834	:douta	=	16'h	39e8;
55835	:douta	=	16'h	3a08;
55836	:douta	=	16'h	39c7;
55837	:douta	=	16'h	39c7;
55838	:douta	=	16'h	39c7;
55839	:douta	=	16'h	39c7;
55840	:douta	=	16'h	39a6;
55841	:douta	=	16'h	41a7;
55842	:douta	=	16'h	41a6;
55843	:douta	=	16'h	39a5;
55844	:douta	=	16'h	3985;
55845	:douta	=	16'h	3964;
55846	:douta	=	16'h	3944;
55847	:douta	=	16'h	3944;
55848	:douta	=	16'h	3943;
55849	:douta	=	16'h	3902;
55850	:douta	=	16'h	3922;
55851	:douta	=	16'h	3923;
55852	:douta	=	16'h	4a4a;
55853	:douta	=	16'h	2146;
55854	:douta	=	16'h	3944;
55855	:douta	=	16'h	59a3;
55856	:douta	=	16'h	59a4;
55857	:douta	=	16'h	59c4;
55858	:douta	=	16'h	61e4;
55859	:douta	=	16'h	59c4;
55860	:douta	=	16'h	61e4;
55861	:douta	=	16'h	6204;
55862	:douta	=	16'h	6204;
55863	:douta	=	16'h	6a04;
55864	:douta	=	16'h	7265;
55865	:douta	=	16'h	83ed;
55866	:douta	=	16'h	82e7;
55867	:douta	=	16'h	7a84;
55868	:douta	=	16'h	7a85;
55869	:douta	=	16'h	7a85;
55870	:douta	=	16'h	7a85;
55871	:douta	=	16'h	82a5;
55872	:douta	=	16'h	82a5;
55873	:douta	=	16'h	82c5;
55874	:douta	=	16'h	8aa5;
55875	:douta	=	16'h	8aa5;
55876	:douta	=	16'h	8ac6;
55877	:douta	=	16'h	8ae6;
55878	:douta	=	16'h	8ac6;
55879	:douta	=	16'h	8ae7;
55880	:douta	=	16'h	9307;
55881	:douta	=	16'h	6205;
55882	:douta	=	16'h	9b47;
55883	:douta	=	16'h	9306;
55884	:douta	=	16'h	9306;
55885	:douta	=	16'h	9306;
55886	:douta	=	16'h	9326;
55887	:douta	=	16'h	9326;
55888	:douta	=	16'h	9327;
55889	:douta	=	16'h	9b46;
55890	:douta	=	16'h	a367;
55891	:douta	=	16'h	ab86;
55892	:douta	=	16'h	aba7;
55893	:douta	=	16'h	b3a7;
55894	:douta	=	16'h	b3c6;
55895	:douta	=	16'h	b3c7;
55896	:douta	=	16'h	bbe7;
55897	:douta	=	16'h	b3c7;
55898	:douta	=	16'h	bbe7;
55899	:douta	=	16'h	bbe7;
55900	:douta	=	16'h	bc07;
55901	:douta	=	16'h	bbe6;
55902	:douta	=	16'h	bc07;
55903	:douta	=	16'h	c407;
55904	:douta	=	16'h	c407;
55905	:douta	=	16'h	c407;
55906	:douta	=	16'h	c447;
55907	:douta	=	16'h	c427;
55908	:douta	=	16'h	c427;
55909	:douta	=	16'h	c427;
55910	:douta	=	16'h	c428;
55911	:douta	=	16'h	c448;
55912	:douta	=	16'h	c428;
55913	:douta	=	16'h	c448;
55914	:douta	=	16'h	cc47;
55915	:douta	=	16'h	c447;
55916	:douta	=	16'h	cc47;
55917	:douta	=	16'h	cc47;
55918	:douta	=	16'h	cc67;
55919	:douta	=	16'h	cc68;
55920	:douta	=	16'h	cc67;
55921	:douta	=	16'h	cc67;
55922	:douta	=	16'h	cc47;
55923	:douta	=	16'h	cc68;
55924	:douta	=	16'h	cc48;
55925	:douta	=	16'h	cc48;
55926	:douta	=	16'h	cc68;
55927	:douta	=	16'h	cc68;
55928	:douta	=	16'h	cc68;
55929	:douta	=	16'h	cc68;
55930	:douta	=	16'h	cc68;
55931	:douta	=	16'h	cc68;
55932	:douta	=	16'h	cc68;
55933	:douta	=	16'h	cc68;
55934	:douta	=	16'h	cc68;
55935	:douta	=	16'h	cc68;
55936	:douta	=	16'h	cc68;
55937	:douta	=	16'h	cc68;
55938	:douta	=	16'h	cc68;
55939	:douta	=	16'h	cc68;
55940	:douta	=	16'h	cc68;
55941	:douta	=	16'h	cc88;
55942	:douta	=	16'h	cc88;
55943	:douta	=	16'h	cc88;
55944	:douta	=	16'h	cc88;
55945	:douta	=	16'h	cc68;
55946	:douta	=	16'h	cc88;
55947	:douta	=	16'h	cc88;
55948	:douta	=	16'h	cc89;
55949	:douta	=	16'h	d4aa;
55950	:douta	=	16'h	d4aa;
55951	:douta	=	16'h	d489;
55952	:douta	=	16'h	d489;
55953	:douta	=	16'h	d488;
55954	:douta	=	16'h	d488;
55955	:douta	=	16'h	cc88;
55956	:douta	=	16'h	cc89;
55957	:douta	=	16'h	d489;
55958	:douta	=	16'h	d489;
55959	:douta	=	16'h	cc89;
55960	:douta	=	16'h	cc88;
55961	:douta	=	16'h	d489;
55962	:douta	=	16'h	cc88;
55963	:douta	=	16'h	d488;
55964	:douta	=	16'h	cc89;
55965	:douta	=	16'h	cc88;
55966	:douta	=	16'h	d4a9;
55967	:douta	=	16'h	cc88;
55968	:douta	=	16'h	d489;
55969	:douta	=	16'h	cc89;
55970	:douta	=	16'h	d488;
55971	:douta	=	16'h	ad53;
55972	:douta	=	16'h	deb7;
55973	:douta	=	16'h	cc26;
55974	:douta	=	16'h	cc89;
55975	:douta	=	16'h	cc89;
55976	:douta	=	16'h	cc89;
55977	:douta	=	16'h	cc68;
55978	:douta	=	16'h	cc89;
55979	:douta	=	16'h	cc69;
55980	:douta	=	16'h	d489;
55981	:douta	=	16'h	cc69;
55982	:douta	=	16'h	cc69;
55983	:douta	=	16'h	cc69;
55984	:douta	=	16'h	cc69;
55985	:douta	=	16'h	cc69;
55986	:douta	=	16'h	d486;
55987	:douta	=	16'h	b44d;
55988	:douta	=	16'h	9430;
55989	:douta	=	16'h	8c31;
55990	:douta	=	16'h	83d0;
55991	:douta	=	16'h	7bd1;
55992	:douta	=	16'h	83f1;
55993	:douta	=	16'h	7bd1;
55994	:douta	=	16'h	73b0;
55995	:douta	=	16'h	7bb1;
55996	:douta	=	16'h	6b4f;
55997	:douta	=	16'h	632f;
55998	:douta	=	16'h	630e;
55999	:douta	=	16'h	62cd;
56000	:douta	=	16'h	62ed;
56001	:douta	=	16'h	5aac;
56002	:douta	=	16'h	734e;
56003	:douta	=	16'h	8411;
56004	:douta	=	16'h	9472;
56005	:douta	=	16'h	8c32;
56006	:douta	=	16'h	83d0;
56007	:douta	=	16'h	7baf;
56008	:douta	=	16'h	5a8c;
56009	:douta	=	16'h	736f;
56010	:douta	=	16'h	628c;
56011	:douta	=	16'h	630d;
56012	:douta	=	16'h	8431;
56013	:douta	=	16'h	be59;
56014	:douta	=	16'h	df5d;
56015	:douta	=	16'h	ffff;
56016	:douta	=	16'h	ffff;
56017	:douta	=	16'h	ffff;
56018	:douta	=	16'h	feb9;
56019	:douta	=	16'h	edf4;
56020	:douta	=	16'h	cba8;
56021	:douta	=	16'h	b322;
56022	:douta	=	16'h	b344;
56023	:douta	=	16'h	b3e8;
56024	:douta	=	16'h	b3e8;
56025	:douta	=	16'h	b3c8;
56026	:douta	=	16'h	b3c8;
56027	:douta	=	16'h	b3c8;
56028	:douta	=	16'h	b3a8;
56029	:douta	=	16'h	b3c9;
56030	:douta	=	16'h	b3a8;
56031	:douta	=	16'h	b3c8;
56032	:douta	=	16'h	b3c8;
56033	:douta	=	16'h	b3c8;
56034	:douta	=	16'h	b3c8;
56035	:douta	=	16'h	b3c8;
56036	:douta	=	16'h	b3c8;
56037	:douta	=	16'h	b3a8;
56038	:douta	=	16'h	aba8;
56039	:douta	=	16'h	aba8;
56040	:douta	=	16'h	b3c9;
56041	:douta	=	16'h	aba8;
56042	:douta	=	16'h	b3c8;
56043	:douta	=	16'h	b3a8;
56044	:douta	=	16'h	b3c8;
56045	:douta	=	16'h	b3a8;
56046	:douta	=	16'h	aba8;
56047	:douta	=	16'h	ab88;
56048	:douta	=	16'h	ab89;
56049	:douta	=	16'h	ab89;
56050	:douta	=	16'h	ab88;
56051	:douta	=	16'h	ab88;
56052	:douta	=	16'h	ab89;
56053	:douta	=	16'h	ab89;
56054	:douta	=	16'h	ab88;
56055	:douta	=	16'h	ab89;
56056	:douta	=	16'h	ab89;
56057	:douta	=	16'h	a368;
56058	:douta	=	16'h	a368;
56059	:douta	=	16'h	a368;
56060	:douta	=	16'h	a368;
56061	:douta	=	16'h	a368;
56062	:douta	=	16'h	ab88;
56063	:douta	=	16'h	ab68;
56064	:douta	=	16'h	a4f6;
56065	:douta	=	16'h	9c94;
56066	:douta	=	16'h	a4f5;
56067	:douta	=	16'h	9cb4;
56068	:douta	=	16'h	ad36;
56069	:douta	=	16'h	ad15;
56070	:douta	=	16'h	8cb6;
56071	:douta	=	16'h	8c96;
56072	:douta	=	16'h	634f;
56073	:douta	=	16'h	28e3;
56074	:douta	=	16'h	2903;
56075	:douta	=	16'h	28e3;
56076	:douta	=	16'h	28e3;
56077	:douta	=	16'h	28e3;
56078	:douta	=	16'h	28e3;
56079	:douta	=	16'h	28e3;
56080	:douta	=	16'h	28e3;
56081	:douta	=	16'h	28e3;
56082	:douta	=	16'h	28e3;
56083	:douta	=	16'h	20a3;
56084	:douta	=	16'h	20c3;
56085	:douta	=	16'h	2082;
56086	:douta	=	16'h	20a3;
56087	:douta	=	16'h	20c3;
56088	:douta	=	16'h	20a2;
56089	:douta	=	16'h	20a2;
56090	:douta	=	16'h	20a2;
56091	:douta	=	16'h	2082;
56092	:douta	=	16'h	20a2;
56093	:douta	=	16'h	20a2;
56094	:douta	=	16'h	20a2;
56095	:douta	=	16'h	20c2;
56096	:douta	=	16'h	20a2;
56097	:douta	=	16'h	28e2;
56098	:douta	=	16'h	30e2;
56099	:douta	=	16'h	30e2;
56100	:douta	=	16'h	3103;
56101	:douta	=	16'h	3123;
56102	:douta	=	16'h	3103;
56103	:douta	=	16'h	4143;
56104	:douta	=	16'h	3923;
56105	:douta	=	16'h	4143;
56106	:douta	=	16'h	4143;
56107	:douta	=	16'h	49a6;
56108	:douta	=	16'h	39e8;
56109	:douta	=	16'h	10e4;
56110	:douta	=	16'h	4985;
56111	:douta	=	16'h	59c4;
56112	:douta	=	16'h	59c4;
56113	:douta	=	16'h	59c4;
56114	:douta	=	16'h	59e4;
56115	:douta	=	16'h	61e4;
56116	:douta	=	16'h	6204;
56117	:douta	=	16'h	6a04;
56118	:douta	=	16'h	6a24;
56119	:douta	=	16'h	6a04;
56120	:douta	=	16'h	6a87;
56121	:douta	=	16'h	94b1;
56122	:douta	=	16'h	7244;
56123	:douta	=	16'h	7a84;
56124	:douta	=	16'h	7a64;
56125	:douta	=	16'h	7a85;
56126	:douta	=	16'h	7a85;
56127	:douta	=	16'h	82a5;
56128	:douta	=	16'h	82a5;
56129	:douta	=	16'h	82a5;
56130	:douta	=	16'h	8aa5;
56131	:douta	=	16'h	8ac6;
56132	:douta	=	16'h	8ac6;
56133	:douta	=	16'h	8ac6;
56134	:douta	=	16'h	8ae6;
56135	:douta	=	16'h	8ac6;
56136	:douta	=	16'h	8ac6;
56137	:douta	=	16'h	7265;
56138	:douta	=	16'h	9b26;
56139	:douta	=	16'h	9306;
56140	:douta	=	16'h	9b47;
56141	:douta	=	16'h	9326;
56142	:douta	=	16'h	9326;
56143	:douta	=	16'h	9326;
56144	:douta	=	16'h	9b27;
56145	:douta	=	16'h	9b26;
56146	:douta	=	16'h	a367;
56147	:douta	=	16'h	a386;
56148	:douta	=	16'h	aba7;
56149	:douta	=	16'h	b3a7;
56150	:douta	=	16'h	b3c6;
56151	:douta	=	16'h	b3c7;
56152	:douta	=	16'h	bbc7;
56153	:douta	=	16'h	bbe7;
56154	:douta	=	16'h	bbe7;
56155	:douta	=	16'h	bbe7;
56156	:douta	=	16'h	bbe7;
56157	:douta	=	16'h	bc07;
56158	:douta	=	16'h	bc07;
56159	:douta	=	16'h	c407;
56160	:douta	=	16'h	c407;
56161	:douta	=	16'h	c427;
56162	:douta	=	16'h	c427;
56163	:douta	=	16'h	c427;
56164	:douta	=	16'h	c427;
56165	:douta	=	16'h	c428;
56166	:douta	=	16'h	c427;
56167	:douta	=	16'h	c428;
56168	:douta	=	16'h	c428;
56169	:douta	=	16'h	c428;
56170	:douta	=	16'h	cc47;
56171	:douta	=	16'h	cc47;
56172	:douta	=	16'h	cc47;
56173	:douta	=	16'h	cc47;
56174	:douta	=	16'h	cc47;
56175	:douta	=	16'h	cc47;
56176	:douta	=	16'h	cc68;
56177	:douta	=	16'h	cc67;
56178	:douta	=	16'h	cc67;
56179	:douta	=	16'h	cc68;
56180	:douta	=	16'h	cc68;
56181	:douta	=	16'h	cc68;
56182	:douta	=	16'h	cc48;
56183	:douta	=	16'h	cc48;
56184	:douta	=	16'h	cc68;
56185	:douta	=	16'h	cc68;
56186	:douta	=	16'h	cc68;
56187	:douta	=	16'h	cc68;
56188	:douta	=	16'h	cc68;
56189	:douta	=	16'h	cc68;
56190	:douta	=	16'h	cc68;
56191	:douta	=	16'h	cc68;
56192	:douta	=	16'h	cc68;
56193	:douta	=	16'h	cc68;
56194	:douta	=	16'h	cc69;
56195	:douta	=	16'h	cc69;
56196	:douta	=	16'h	cc88;
56197	:douta	=	16'h	cc88;
56198	:douta	=	16'h	cc88;
56199	:douta	=	16'h	cc88;
56200	:douta	=	16'h	cc88;
56201	:douta	=	16'h	cc88;
56202	:douta	=	16'h	cc89;
56203	:douta	=	16'h	cc89;
56204	:douta	=	16'h	cc88;
56205	:douta	=	16'h	cc88;
56206	:douta	=	16'h	cc68;
56207	:douta	=	16'h	cc88;
56208	:douta	=	16'h	cc88;
56209	:douta	=	16'h	d488;
56210	:douta	=	16'h	d488;
56211	:douta	=	16'h	d488;
56212	:douta	=	16'h	cc89;
56213	:douta	=	16'h	cc89;
56214	:douta	=	16'h	cc89;
56215	:douta	=	16'h	cc89;
56216	:douta	=	16'h	d488;
56217	:douta	=	16'h	d489;
56218	:douta	=	16'h	d488;
56219	:douta	=	16'h	cc88;
56220	:douta	=	16'h	d489;
56221	:douta	=	16'h	d489;
56222	:douta	=	16'h	cc89;
56223	:douta	=	16'h	cc89;
56224	:douta	=	16'h	cc89;
56225	:douta	=	16'h	cc89;
56226	:douta	=	16'h	d488;
56227	:douta	=	16'h	ad33;
56228	:douta	=	16'h	deb7;
56229	:douta	=	16'h	cc26;
56230	:douta	=	16'h	cc89;
56231	:douta	=	16'h	cc89;
56232	:douta	=	16'h	cc69;
56233	:douta	=	16'h	cc89;
56234	:douta	=	16'h	cc89;
56235	:douta	=	16'h	cc89;
56236	:douta	=	16'h	cc69;
56237	:douta	=	16'h	cc89;
56238	:douta	=	16'h	cc69;
56239	:douta	=	16'h	cc68;
56240	:douta	=	16'h	cc49;
56241	:douta	=	16'h	cc69;
56242	:douta	=	16'h	cc69;
56243	:douta	=	16'h	dc86;
56244	:douta	=	16'h	7bf1;
56245	:douta	=	16'h	9431;
56246	:douta	=	16'h	8411;
56247	:douta	=	16'h	7390;
56248	:douta	=	16'h	738f;
56249	:douta	=	16'h	6b6f;
56250	:douta	=	16'h	6b4f;
56251	:douta	=	16'h	6b4f;
56252	:douta	=	16'h	5aed;
56253	:douta	=	16'h	4a6b;
56254	:douta	=	16'h	422b;
56255	:douta	=	16'h	62ee;
56256	:douta	=	16'h	528d;
56257	:douta	=	16'h	acd4;
56258	:douta	=	16'h	7bb0;
56259	:douta	=	16'h	7b90;
56260	:douta	=	16'h	7b90;
56261	:douta	=	16'h	62cd;
56262	:douta	=	16'h	6b4f;
56263	:douta	=	16'h	8431;
56264	:douta	=	16'h	add7;
56265	:douta	=	16'h	d71d;
56266	:douta	=	16'h	ffff;
56267	:douta	=	16'h	ffff;
56268	:douta	=	16'h	ff9c;
56269	:douta	=	16'h	e5d3;
56270	:douta	=	16'h	dd0e;
56271	:douta	=	16'h	cbc7;
56272	:douta	=	16'h	bb64;
56273	:douta	=	16'h	bba5;
56274	:douta	=	16'h	bc08;
56275	:douta	=	16'h	bc08;
56276	:douta	=	16'h	bc09;
56277	:douta	=	16'h	bbe8;
56278	:douta	=	16'h	bbe9;
56279	:douta	=	16'h	b3c9;
56280	:douta	=	16'h	bbe9;
56281	:douta	=	16'h	b3e9;
56282	:douta	=	16'h	b3c8;
56283	:douta	=	16'h	bbc9;
56284	:douta	=	16'h	b3e9;
56285	:douta	=	16'h	b3e9;
56286	:douta	=	16'h	b3e9;
56287	:douta	=	16'h	b3c8;
56288	:douta	=	16'h	b3c8;
56289	:douta	=	16'h	b3c8;
56290	:douta	=	16'h	b3c8;
56291	:douta	=	16'h	b3a8;
56292	:douta	=	16'h	b3c8;
56293	:douta	=	16'h	b3a8;
56294	:douta	=	16'h	b3c8;
56295	:douta	=	16'h	b3a8;
56296	:douta	=	16'h	b3a8;
56297	:douta	=	16'h	b3c8;
56298	:douta	=	16'h	b3c8;
56299	:douta	=	16'h	b3c8;
56300	:douta	=	16'h	b3a8;
56301	:douta	=	16'h	b3c8;
56302	:douta	=	16'h	b3c8;
56303	:douta	=	16'h	aba8;
56304	:douta	=	16'h	b3a8;
56305	:douta	=	16'h	b3a8;
56306	:douta	=	16'h	ab88;
56307	:douta	=	16'h	ab88;
56308	:douta	=	16'h	ab89;
56309	:douta	=	16'h	ab88;
56310	:douta	=	16'h	ab88;
56311	:douta	=	16'h	ab88;
56312	:douta	=	16'h	ab89;
56313	:douta	=	16'h	ab89;
56314	:douta	=	16'h	a368;
56315	:douta	=	16'h	ab88;
56316	:douta	=	16'h	a368;
56317	:douta	=	16'h	ab88;
56318	:douta	=	16'h	ab68;
56319	:douta	=	16'h	a368;
56320	:douta	=	16'h	9cb5;
56321	:douta	=	16'h	9c94;
56322	:douta	=	16'h	a516;
56323	:douta	=	16'h	a4f4;
56324	:douta	=	16'h	ad16;
56325	:douta	=	16'h	ad15;
56326	:douta	=	16'h	8cb6;
56327	:douta	=	16'h	94d6;
56328	:douta	=	16'h	422a;
56329	:douta	=	16'h	2903;
56330	:douta	=	16'h	2903;
56331	:douta	=	16'h	28e3;
56332	:douta	=	16'h	28e3;
56333	:douta	=	16'h	28e3;
56334	:douta	=	16'h	28e3;
56335	:douta	=	16'h	28e3;
56336	:douta	=	16'h	20e3;
56337	:douta	=	16'h	28e3;
56338	:douta	=	16'h	28e3;
56339	:douta	=	16'h	20c3;
56340	:douta	=	16'h	20c3;
56341	:douta	=	16'h	18c3;
56342	:douta	=	16'h	20c3;
56343	:douta	=	16'h	2082;
56344	:douta	=	16'h	20a2;
56345	:douta	=	16'h	20a3;
56346	:douta	=	16'h	20a3;
56347	:douta	=	16'h	20a3;
56348	:douta	=	16'h	20c2;
56349	:douta	=	16'h	20c2;
56350	:douta	=	16'h	20c2;
56351	:douta	=	16'h	20c2;
56352	:douta	=	16'h	20c2;
56353	:douta	=	16'h	28e3;
56354	:douta	=	16'h	30e3;
56355	:douta	=	16'h	3103;
56356	:douta	=	16'h	3103;
56357	:douta	=	16'h	3103;
56358	:douta	=	16'h	3923;
56359	:douta	=	16'h	4124;
56360	:douta	=	16'h	4123;
56361	:douta	=	16'h	4143;
56362	:douta	=	16'h	4163;
56363	:douta	=	16'h	49c7;
56364	:douta	=	16'h	31a8;
56365	:douta	=	16'h	10c4;
56366	:douta	=	16'h	51a5;
56367	:douta	=	16'h	59c4;
56368	:douta	=	16'h	59c4;
56369	:douta	=	16'h	61c4;
56370	:douta	=	16'h	61e4;
56371	:douta	=	16'h	61e4;
56372	:douta	=	16'h	6204;
56373	:douta	=	16'h	6a04;
56374	:douta	=	16'h	6a04;
56375	:douta	=	16'h	7224;
56376	:douta	=	16'h	72c9;
56377	:douta	=	16'h	a533;
56378	:douta	=	16'h	7203;
56379	:douta	=	16'h	7a64;
56380	:douta	=	16'h	7a84;
56381	:douta	=	16'h	7a85;
56382	:douta	=	16'h	7a85;
56383	:douta	=	16'h	82c6;
56384	:douta	=	16'h	82a5;
56385	:douta	=	16'h	82c5;
56386	:douta	=	16'h	8aa5;
56387	:douta	=	16'h	8aa5;
56388	:douta	=	16'h	8aa5;
56389	:douta	=	16'h	8ac6;
56390	:douta	=	16'h	8ae6;
56391	:douta	=	16'h	8ac6;
56392	:douta	=	16'h	8ae6;
56393	:douta	=	16'h	7264;
56394	:douta	=	16'h	9b26;
56395	:douta	=	16'h	9326;
56396	:douta	=	16'h	9b47;
56397	:douta	=	16'h	9b47;
56398	:douta	=	16'h	9306;
56399	:douta	=	16'h	9326;
56400	:douta	=	16'h	9327;
56401	:douta	=	16'h	9b26;
56402	:douta	=	16'h	a367;
56403	:douta	=	16'h	ab87;
56404	:douta	=	16'h	ab87;
56405	:douta	=	16'h	b3c7;
56406	:douta	=	16'h	b3c6;
56407	:douta	=	16'h	b3c7;
56408	:douta	=	16'h	bbe8;
56409	:douta	=	16'h	bbe8;
56410	:douta	=	16'h	bbe7;
56411	:douta	=	16'h	bbe7;
56412	:douta	=	16'h	bbe7;
56413	:douta	=	16'h	bbe7;
56414	:douta	=	16'h	bbe7;
56415	:douta	=	16'h	c407;
56416	:douta	=	16'h	c427;
56417	:douta	=	16'h	c427;
56418	:douta	=	16'h	c427;
56419	:douta	=	16'h	c428;
56420	:douta	=	16'h	c427;
56421	:douta	=	16'h	c428;
56422	:douta	=	16'h	c427;
56423	:douta	=	16'h	c428;
56424	:douta	=	16'h	c428;
56425	:douta	=	16'h	c448;
56426	:douta	=	16'h	cc47;
56427	:douta	=	16'h	cc47;
56428	:douta	=	16'h	cc47;
56429	:douta	=	16'h	cc47;
56430	:douta	=	16'h	cc47;
56431	:douta	=	16'h	cc67;
56432	:douta	=	16'h	cc67;
56433	:douta	=	16'h	cc67;
56434	:douta	=	16'h	cc68;
56435	:douta	=	16'h	cc67;
56436	:douta	=	16'h	cc67;
56437	:douta	=	16'h	cc68;
56438	:douta	=	16'h	cc68;
56439	:douta	=	16'h	cc48;
56440	:douta	=	16'h	cc68;
56441	:douta	=	16'h	cc68;
56442	:douta	=	16'h	cc68;
56443	:douta	=	16'h	cc68;
56444	:douta	=	16'h	cc68;
56445	:douta	=	16'h	cc68;
56446	:douta	=	16'h	cc48;
56447	:douta	=	16'h	cc68;
56448	:douta	=	16'h	cc68;
56449	:douta	=	16'h	cc69;
56450	:douta	=	16'h	cc69;
56451	:douta	=	16'h	cc69;
56452	:douta	=	16'h	cc89;
56453	:douta	=	16'h	d488;
56454	:douta	=	16'h	cc88;
56455	:douta	=	16'h	cc88;
56456	:douta	=	16'h	cc88;
56457	:douta	=	16'h	cc88;
56458	:douta	=	16'h	cc89;
56459	:douta	=	16'h	cc89;
56460	:douta	=	16'h	cc89;
56461	:douta	=	16'h	cc89;
56462	:douta	=	16'h	cc89;
56463	:douta	=	16'h	d489;
56464	:douta	=	16'h	cc89;
56465	:douta	=	16'h	cc89;
56466	:douta	=	16'h	d489;
56467	:douta	=	16'h	d489;
56468	:douta	=	16'h	cc89;
56469	:douta	=	16'h	d489;
56470	:douta	=	16'h	cc89;
56471	:douta	=	16'h	d489;
56472	:douta	=	16'h	d488;
56473	:douta	=	16'h	cc89;
56474	:douta	=	16'h	cc89;
56475	:douta	=	16'h	d489;
56476	:douta	=	16'h	d489;
56477	:douta	=	16'h	d489;
56478	:douta	=	16'h	cc89;
56479	:douta	=	16'h	cc69;
56480	:douta	=	16'h	cc89;
56481	:douta	=	16'h	cc89;
56482	:douta	=	16'h	d488;
56483	:douta	=	16'h	ad53;
56484	:douta	=	16'h	e6b7;
56485	:douta	=	16'h	cc27;
56486	:douta	=	16'h	cc89;
56487	:douta	=	16'h	cc89;
56488	:douta	=	16'h	cc69;
56489	:douta	=	16'h	cc69;
56490	:douta	=	16'h	cc89;
56491	:douta	=	16'h	cc89;
56492	:douta	=	16'h	cc89;
56493	:douta	=	16'h	cc89;
56494	:douta	=	16'h	cc89;
56495	:douta	=	16'h	cc89;
56496	:douta	=	16'h	cc69;
56497	:douta	=	16'h	cc69;
56498	:douta	=	16'h	cc69;
56499	:douta	=	16'h	d487;
56500	:douta	=	16'h	7bd0;
56501	:douta	=	16'h	7bcf;
56502	:douta	=	16'h	83f0;
56503	:douta	=	16'h	7390;
56504	:douta	=	16'h	6b6e;
56505	:douta	=	16'h	6b2f;
56506	:douta	=	16'h	6b2e;
56507	:douta	=	16'h	528c;
56508	:douta	=	16'h	528c;
56509	:douta	=	16'h	632e;
56510	:douta	=	16'h	83f1;
56511	:douta	=	16'h	9473;
56512	:douta	=	16'h	31cb;
56513	:douta	=	16'h	9411;
56514	:douta	=	16'h	62ed;
56515	:douta	=	16'h	62cd;
56516	:douta	=	16'h	630e;
56517	:douta	=	16'h	7c13;
56518	:douta	=	16'h	c69b;
56519	:douta	=	16'h	ef9f;
56520	:douta	=	16'h	ffff;
56521	:douta	=	16'h	ff9e;
56522	:douta	=	16'h	e615;
56523	:douta	=	16'h	d48c;
56524	:douta	=	16'h	cc09;
56525	:douta	=	16'h	bb85;
56526	:douta	=	16'h	bb85;
56527	:douta	=	16'h	bc28;
56528	:douta	=	16'h	c429;
56529	:douta	=	16'h	bc09;
56530	:douta	=	16'h	bc09;
56531	:douta	=	16'h	bc08;
56532	:douta	=	16'h	bbe8;
56533	:douta	=	16'h	bc08;
56534	:douta	=	16'h	bc09;
56535	:douta	=	16'h	bbe9;
56536	:douta	=	16'h	bbe9;
56537	:douta	=	16'h	bbe9;
56538	:douta	=	16'h	bbe9;
56539	:douta	=	16'h	b3e9;
56540	:douta	=	16'h	b3e8;
56541	:douta	=	16'h	b3c9;
56542	:douta	=	16'h	bbe9;
56543	:douta	=	16'h	b3e9;
56544	:douta	=	16'h	b3c9;
56545	:douta	=	16'h	b3c8;
56546	:douta	=	16'h	b3c8;
56547	:douta	=	16'h	b3e9;
56548	:douta	=	16'h	b3a8;
56549	:douta	=	16'h	b3c8;
56550	:douta	=	16'h	b3c8;
56551	:douta	=	16'h	b3a8;
56552	:douta	=	16'h	b3a8;
56553	:douta	=	16'h	b3a9;
56554	:douta	=	16'h	b3a9;
56555	:douta	=	16'h	b3c9;
56556	:douta	=	16'h	b3c8;
56557	:douta	=	16'h	b3a8;
56558	:douta	=	16'h	b3c8;
56559	:douta	=	16'h	aba8;
56560	:douta	=	16'h	ab88;
56561	:douta	=	16'h	b3a8;
56562	:douta	=	16'h	ab88;
56563	:douta	=	16'h	aba9;
56564	:douta	=	16'h	ab89;
56565	:douta	=	16'h	aba9;
56566	:douta	=	16'h	ab88;
56567	:douta	=	16'h	ab88;
56568	:douta	=	16'h	ab88;
56569	:douta	=	16'h	ab88;
56570	:douta	=	16'h	ab88;
56571	:douta	=	16'h	a368;
56572	:douta	=	16'h	ab68;
56573	:douta	=	16'h	ab89;
56574	:douta	=	16'h	a368;
56575	:douta	=	16'h	a368;
56576	:douta	=	16'h	9474;
56577	:douta	=	16'h	9cb4;
56578	:douta	=	16'h	a516;
56579	:douta	=	16'h	b534;
56580	:douta	=	16'h	ad15;
56581	:douta	=	16'h	9cd6;
56582	:douta	=	16'h	94d6;
56583	:douta	=	16'h	8cd7;
56584	:douta	=	16'h	2104;
56585	:douta	=	16'h	28e3;
56586	:douta	=	16'h	2903;
56587	:douta	=	16'h	28e3;
56588	:douta	=	16'h	28e3;
56589	:douta	=	16'h	28e3;
56590	:douta	=	16'h	28e3;
56591	:douta	=	16'h	28e3;
56592	:douta	=	16'h	28e3;
56593	:douta	=	16'h	20c3;
56594	:douta	=	16'h	20c3;
56595	:douta	=	16'h	28e3;
56596	:douta	=	16'h	20c3;
56597	:douta	=	16'h	20a3;
56598	:douta	=	16'h	20e3;
56599	:douta	=	16'h	18a1;
56600	:douta	=	16'h	20c2;
56601	:douta	=	16'h	20a2;
56602	:douta	=	16'h	20e3;
56603	:douta	=	16'h	20c2;
56604	:douta	=	16'h	20a2;
56605	:douta	=	16'h	28c3;
56606	:douta	=	16'h	20a2;
56607	:douta	=	16'h	28e3;
56608	:douta	=	16'h	28e3;
56609	:douta	=	16'h	30e3;
56610	:douta	=	16'h	30e3;
56611	:douta	=	16'h	3103;
56612	:douta	=	16'h	3103;
56613	:douta	=	16'h	3923;
56614	:douta	=	16'h	3923;
56615	:douta	=	16'h	3943;
56616	:douta	=	16'h	4124;
56617	:douta	=	16'h	4163;
56618	:douta	=	16'h	4143;
56619	:douta	=	16'h	4a08;
56620	:douta	=	16'h	2146;
56621	:douta	=	16'h	0884;
56622	:douta	=	16'h	59c4;
56623	:douta	=	16'h	51a4;
56624	:douta	=	16'h	59e5;
56625	:douta	=	16'h	61c4;
56626	:douta	=	16'h	61c4;
56627	:douta	=	16'h	6204;
56628	:douta	=	16'h	6a04;
56629	:douta	=	16'h	6a04;
56630	:douta	=	16'h	6a04;
56631	:douta	=	16'h	6a24;
56632	:douta	=	16'h	734b;
56633	:douta	=	16'h	ad53;
56634	:douta	=	16'h	71e3;
56635	:douta	=	16'h	7a64;
56636	:douta	=	16'h	7a84;
56637	:douta	=	16'h	7a85;
56638	:douta	=	16'h	7a85;
56639	:douta	=	16'h	82a5;
56640	:douta	=	16'h	82c5;
56641	:douta	=	16'h	82a5;
56642	:douta	=	16'h	8ac6;
56643	:douta	=	16'h	8ac6;
56644	:douta	=	16'h	8ae6;
56645	:douta	=	16'h	8ac6;
56646	:douta	=	16'h	92e7;
56647	:douta	=	16'h	9307;
56648	:douta	=	16'h	9307;
56649	:douta	=	16'h	7244;
56650	:douta	=	16'h	9b47;
56651	:douta	=	16'h	9326;
56652	:douta	=	16'h	9326;
56653	:douta	=	16'h	9b47;
56654	:douta	=	16'h	9306;
56655	:douta	=	16'h	9326;
56656	:douta	=	16'h	9327;
56657	:douta	=	16'h	9b67;
56658	:douta	=	16'h	a367;
56659	:douta	=	16'h	ab87;
56660	:douta	=	16'h	b3a7;
56661	:douta	=	16'h	b3c6;
56662	:douta	=	16'h	b3c7;
56663	:douta	=	16'h	b3c7;
56664	:douta	=	16'h	b3c7;
56665	:douta	=	16'h	bbe7;
56666	:douta	=	16'h	bbe7;
56667	:douta	=	16'h	bbe7;
56668	:douta	=	16'h	bc07;
56669	:douta	=	16'h	bc07;
56670	:douta	=	16'h	bc07;
56671	:douta	=	16'h	bc07;
56672	:douta	=	16'h	c407;
56673	:douta	=	16'h	c427;
56674	:douta	=	16'h	c428;
56675	:douta	=	16'h	c428;
56676	:douta	=	16'h	c428;
56677	:douta	=	16'h	c427;
56678	:douta	=	16'h	c428;
56679	:douta	=	16'h	c448;
56680	:douta	=	16'h	c448;
56681	:douta	=	16'h	c448;
56682	:douta	=	16'h	c428;
56683	:douta	=	16'h	c448;
56684	:douta	=	16'h	cc48;
56685	:douta	=	16'h	c448;
56686	:douta	=	16'h	cc47;
56687	:douta	=	16'h	cc47;
56688	:douta	=	16'h	cc47;
56689	:douta	=	16'h	cc68;
56690	:douta	=	16'h	cc68;
56691	:douta	=	16'h	cc68;
56692	:douta	=	16'h	cc68;
56693	:douta	=	16'h	cc68;
56694	:douta	=	16'h	cc67;
56695	:douta	=	16'h	cc67;
56696	:douta	=	16'h	cc68;
56697	:douta	=	16'h	cc68;
56698	:douta	=	16'h	cc68;
56699	:douta	=	16'h	cc68;
56700	:douta	=	16'h	cc68;
56701	:douta	=	16'h	cc68;
56702	:douta	=	16'h	cc68;
56703	:douta	=	16'h	cc68;
56704	:douta	=	16'h	cc69;
56705	:douta	=	16'h	cc69;
56706	:douta	=	16'h	cc48;
56707	:douta	=	16'h	cc69;
56708	:douta	=	16'h	cc68;
56709	:douta	=	16'h	cc88;
56710	:douta	=	16'h	cc88;
56711	:douta	=	16'h	cc88;
56712	:douta	=	16'h	d488;
56713	:douta	=	16'h	d4a9;
56714	:douta	=	16'h	cc69;
56715	:douta	=	16'h	cc89;
56716	:douta	=	16'h	d489;
56717	:douta	=	16'h	cc89;
56718	:douta	=	16'h	d489;
56719	:douta	=	16'h	cc89;
56720	:douta	=	16'h	d4a9;
56721	:douta	=	16'h	d489;
56722	:douta	=	16'h	d489;
56723	:douta	=	16'h	d489;
56724	:douta	=	16'h	d489;
56725	:douta	=	16'h	cc89;
56726	:douta	=	16'h	cc89;
56727	:douta	=	16'h	cc89;
56728	:douta	=	16'h	d488;
56729	:douta	=	16'h	cc89;
56730	:douta	=	16'h	cc89;
56731	:douta	=	16'h	d489;
56732	:douta	=	16'h	d489;
56733	:douta	=	16'h	cc89;
56734	:douta	=	16'h	cc89;
56735	:douta	=	16'h	cc89;
56736	:douta	=	16'h	cc89;
56737	:douta	=	16'h	cc89;
56738	:douta	=	16'h	d468;
56739	:douta	=	16'h	ad53;
56740	:douta	=	16'h	deb7;
56741	:douta	=	16'h	cc27;
56742	:douta	=	16'h	cc69;
56743	:douta	=	16'h	cc89;
56744	:douta	=	16'h	cc69;
56745	:douta	=	16'h	cc69;
56746	:douta	=	16'h	cc69;
56747	:douta	=	16'h	cc89;
56748	:douta	=	16'h	cc69;
56749	:douta	=	16'h	cc89;
56750	:douta	=	16'h	cc69;
56751	:douta	=	16'h	cc69;
56752	:douta	=	16'h	cc69;
56753	:douta	=	16'h	cc69;
56754	:douta	=	16'h	cc68;
56755	:douta	=	16'h	cc6a;
56756	:douta	=	16'h	c469;
56757	:douta	=	16'h	8bef;
56758	:douta	=	16'h	732f;
56759	:douta	=	16'h	528c;
56760	:douta	=	16'h	62ed;
56761	:douta	=	16'h	7bf1;
56762	:douta	=	16'h	8c32;
56763	:douta	=	16'h	9493;
56764	:douta	=	16'h	8c53;
56765	:douta	=	16'h	5acd;
56766	:douta	=	16'h	8c53;
56767	:douta	=	16'h	9d17;
56768	:douta	=	16'h	953a;
56769	:douta	=	16'h	b6bf;
56770	:douta	=	16'h	c73f;
56771	:douta	=	16'h	e7bf;
56772	:douta	=	16'h	e75e;
56773	:douta	=	16'h	d593;
56774	:douta	=	16'h	c46b;
56775	:douta	=	16'h	c3e7;
56776	:douta	=	16'h	bba4;
56777	:douta	=	16'h	c3e6;
56778	:douta	=	16'h	c449;
56779	:douta	=	16'h	c428;
56780	:douta	=	16'h	c428;
56781	:douta	=	16'h	c429;
56782	:douta	=	16'h	c429;
56783	:douta	=	16'h	c429;
56784	:douta	=	16'h	bc28;
56785	:douta	=	16'h	bc09;
56786	:douta	=	16'h	bc08;
56787	:douta	=	16'h	bc09;
56788	:douta	=	16'h	bbe9;
56789	:douta	=	16'h	bc08;
56790	:douta	=	16'h	bc09;
56791	:douta	=	16'h	bc09;
56792	:douta	=	16'h	bbe9;
56793	:douta	=	16'h	bbe9;
56794	:douta	=	16'h	bbe9;
56795	:douta	=	16'h	bbe9;
56796	:douta	=	16'h	bbe9;
56797	:douta	=	16'h	bbe9;
56798	:douta	=	16'h	b3c8;
56799	:douta	=	16'h	b3e8;
56800	:douta	=	16'h	b3e8;
56801	:douta	=	16'h	b3e9;
56802	:douta	=	16'h	b3c9;
56803	:douta	=	16'h	b3c9;
56804	:douta	=	16'h	b3c9;
56805	:douta	=	16'h	b3c9;
56806	:douta	=	16'h	b3a8;
56807	:douta	=	16'h	b3a8;
56808	:douta	=	16'h	b3c8;
56809	:douta	=	16'h	b3a9;
56810	:douta	=	16'h	b3a9;
56811	:douta	=	16'h	b3c8;
56812	:douta	=	16'h	b3c8;
56813	:douta	=	16'h	b3c8;
56814	:douta	=	16'h	b3a8;
56815	:douta	=	16'h	b3c8;
56816	:douta	=	16'h	b3a8;
56817	:douta	=	16'h	b3a8;
56818	:douta	=	16'h	aba9;
56819	:douta	=	16'h	aba9;
56820	:douta	=	16'h	aba9;
56821	:douta	=	16'h	ab88;
56822	:douta	=	16'h	aba9;
56823	:douta	=	16'h	a388;
56824	:douta	=	16'h	aba9;
56825	:douta	=	16'h	ab89;
56826	:douta	=	16'h	ab88;
56827	:douta	=	16'h	ab89;
56828	:douta	=	16'h	ab88;
56829	:douta	=	16'h	a368;
56830	:douta	=	16'h	ab68;
56831	:douta	=	16'h	a388;
56832	:douta	=	16'h	9c94;
56833	:douta	=	16'h	9cd4;
56834	:douta	=	16'h	a516;
56835	:douta	=	16'h	b555;
56836	:douta	=	16'h	a516;
56837	:douta	=	16'h	8cb5;
56838	:douta	=	16'h	94f6;
56839	:douta	=	16'h	9518;
56840	:douta	=	16'h	1861;
56841	:douta	=	16'h	2924;
56842	:douta	=	16'h	28e3;
56843	:douta	=	16'h	28e3;
56844	:douta	=	16'h	28e3;
56845	:douta	=	16'h	28e3;
56846	:douta	=	16'h	20c2;
56847	:douta	=	16'h	28e3;
56848	:douta	=	16'h	28e3;
56849	:douta	=	16'h	28e3;
56850	:douta	=	16'h	28e3;
56851	:douta	=	16'h	20c3;
56852	:douta	=	16'h	20c3;
56853	:douta	=	16'h	20c3;
56854	:douta	=	16'h	20e3;
56855	:douta	=	16'h	20a2;
56856	:douta	=	16'h	20c2;
56857	:douta	=	16'h	20c2;
56858	:douta	=	16'h	20a2;
56859	:douta	=	16'h	20c2;
56860	:douta	=	16'h	20c2;
56861	:douta	=	16'h	28e3;
56862	:douta	=	16'h	28c3;
56863	:douta	=	16'h	28e2;
56864	:douta	=	16'h	28c2;
56865	:douta	=	16'h	3103;
56866	:douta	=	16'h	3103;
56867	:douta	=	16'h	3103;
56868	:douta	=	16'h	3103;
56869	:douta	=	16'h	3123;
56870	:douta	=	16'h	3923;
56871	:douta	=	16'h	4143;
56872	:douta	=	16'h	4144;
56873	:douta	=	16'h	4163;
56874	:douta	=	16'h	4964;
56875	:douta	=	16'h	4a49;
56876	:douta	=	16'h	1906;
56877	:douta	=	16'h	10a4;
56878	:douta	=	16'h	61c4;
56879	:douta	=	16'h	59c4;
56880	:douta	=	16'h	59c4;
56881	:douta	=	16'h	61e4;
56882	:douta	=	16'h	61e4;
56883	:douta	=	16'h	6204;
56884	:douta	=	16'h	6a04;
56885	:douta	=	16'h	6a04;
56886	:douta	=	16'h	7224;
56887	:douta	=	16'h	69e4;
56888	:douta	=	16'h	7bad;
56889	:douta	=	16'h	ad31;
56890	:douta	=	16'h	7a04;
56891	:douta	=	16'h	7a84;
56892	:douta	=	16'h	7a64;
56893	:douta	=	16'h	8285;
56894	:douta	=	16'h	7a85;
56895	:douta	=	16'h	82a5;
56896	:douta	=	16'h	8aa5;
56897	:douta	=	16'h	8aa5;
56898	:douta	=	16'h	8ac6;
56899	:douta	=	16'h	8aa5;
56900	:douta	=	16'h	8aa5;
56901	:douta	=	16'h	8ac6;
56902	:douta	=	16'h	8ac6;
56903	:douta	=	16'h	8ae6;
56904	:douta	=	16'h	9307;
56905	:douta	=	16'h	7265;
56906	:douta	=	16'h	9b47;
56907	:douta	=	16'h	9327;
56908	:douta	=	16'h	9b26;
56909	:douta	=	16'h	9b27;
56910	:douta	=	16'h	92e6;
56911	:douta	=	16'h	9327;
56912	:douta	=	16'h	9326;
56913	:douta	=	16'h	a346;
56914	:douta	=	16'h	ab87;
56915	:douta	=	16'h	ab86;
56916	:douta	=	16'h	aba7;
56917	:douta	=	16'h	aba6;
56918	:douta	=	16'h	b3e7;
56919	:douta	=	16'h	b3e6;
56920	:douta	=	16'h	b3e6;
56921	:douta	=	16'h	b3e6;
56922	:douta	=	16'h	bbe7;
56923	:douta	=	16'h	bc07;
56924	:douta	=	16'h	bbe7;
56925	:douta	=	16'h	bc07;
56926	:douta	=	16'h	bc07;
56927	:douta	=	16'h	bc07;
56928	:douta	=	16'h	c407;
56929	:douta	=	16'h	c407;
56930	:douta	=	16'h	c428;
56931	:douta	=	16'h	c427;
56932	:douta	=	16'h	c428;
56933	:douta	=	16'h	c448;
56934	:douta	=	16'h	c448;
56935	:douta	=	16'h	c448;
56936	:douta	=	16'h	c448;
56937	:douta	=	16'h	c448;
56938	:douta	=	16'h	cc47;
56939	:douta	=	16'h	cc47;
56940	:douta	=	16'h	c448;
56941	:douta	=	16'h	cc48;
56942	:douta	=	16'h	cc48;
56943	:douta	=	16'h	cc67;
56944	:douta	=	16'h	cc68;
56945	:douta	=	16'h	cc47;
56946	:douta	=	16'h	cc68;
56947	:douta	=	16'h	cc47;
56948	:douta	=	16'h	cc68;
56949	:douta	=	16'h	cc68;
56950	:douta	=	16'h	cc68;
56951	:douta	=	16'h	cc68;
56952	:douta	=	16'h	cc88;
56953	:douta	=	16'h	cc68;
56954	:douta	=	16'h	cc68;
56955	:douta	=	16'h	cc68;
56956	:douta	=	16'h	cc48;
56957	:douta	=	16'h	cc68;
56958	:douta	=	16'h	cc68;
56959	:douta	=	16'h	cc69;
56960	:douta	=	16'h	cc69;
56961	:douta	=	16'h	cc69;
56962	:douta	=	16'h	cc68;
56963	:douta	=	16'h	cc68;
56964	:douta	=	16'h	cc68;
56965	:douta	=	16'h	cc68;
56966	:douta	=	16'h	cc68;
56967	:douta	=	16'h	cc88;
56968	:douta	=	16'h	cc89;
56969	:douta	=	16'h	cc89;
56970	:douta	=	16'h	cc89;
56971	:douta	=	16'h	cc89;
56972	:douta	=	16'h	cc89;
56973	:douta	=	16'h	d489;
56974	:douta	=	16'h	cc69;
56975	:douta	=	16'h	d489;
56976	:douta	=	16'h	cc89;
56977	:douta	=	16'h	cc89;
56978	:douta	=	16'h	d489;
56979	:douta	=	16'h	cc89;
56980	:douta	=	16'h	d489;
56981	:douta	=	16'h	d489;
56982	:douta	=	16'h	d489;
56983	:douta	=	16'h	d489;
56984	:douta	=	16'h	d489;
56985	:douta	=	16'h	cc89;
56986	:douta	=	16'h	cc89;
56987	:douta	=	16'h	d489;
56988	:douta	=	16'h	d489;
56989	:douta	=	16'h	cc89;
56990	:douta	=	16'h	d4a9;
56991	:douta	=	16'h	cc89;
56992	:douta	=	16'h	cc88;
56993	:douta	=	16'h	cc89;
56994	:douta	=	16'h	d468;
56995	:douta	=	16'h	ad53;
56996	:douta	=	16'h	e6b7;
56997	:douta	=	16'h	cc47;
56998	:douta	=	16'h	cc69;
56999	:douta	=	16'h	cc89;
57000	:douta	=	16'h	cc69;
57001	:douta	=	16'h	cc69;
57002	:douta	=	16'h	cc89;
57003	:douta	=	16'h	cc89;
57004	:douta	=	16'h	cc69;
57005	:douta	=	16'h	cc69;
57006	:douta	=	16'h	cc89;
57007	:douta	=	16'h	cc69;
57008	:douta	=	16'h	cc69;
57009	:douta	=	16'h	cc69;
57010	:douta	=	16'h	cc68;
57011	:douta	=	16'h	cc69;
57012	:douta	=	16'h	d487;
57013	:douta	=	16'h	cc69;
57014	:douta	=	16'h	7bf1;
57015	:douta	=	16'h	630e;
57016	:douta	=	16'h	8c74;
57017	:douta	=	16'h	8c95;
57018	:douta	=	16'h	94f6;
57019	:douta	=	16'h	7bd3;
57020	:douta	=	16'h	7bf1;
57021	:douta	=	16'h	9518;
57022	:douta	=	16'h	df7f;
57023	:douta	=	16'h	e7ff;
57024	:douta	=	16'h	dfff;
57025	:douta	=	16'h	d6de;
57026	:douta	=	16'h	ce18;
57027	:douta	=	16'h	c48e;
57028	:douta	=	16'h	c40a;
57029	:douta	=	16'h	bba4;
57030	:douta	=	16'h	c407;
57031	:douta	=	16'h	cc28;
57032	:douta	=	16'h	c449;
57033	:douta	=	16'h	c449;
57034	:douta	=	16'h	c428;
57035	:douta	=	16'h	c429;
57036	:douta	=	16'h	c429;
57037	:douta	=	16'h	c429;
57038	:douta	=	16'h	c429;
57039	:douta	=	16'h	c429;
57040	:douta	=	16'h	bc08;
57041	:douta	=	16'h	bc08;
57042	:douta	=	16'h	c429;
57043	:douta	=	16'h	bc09;
57044	:douta	=	16'h	bc09;
57045	:douta	=	16'h	bc09;
57046	:douta	=	16'h	bc09;
57047	:douta	=	16'h	bc09;
57048	:douta	=	16'h	bc09;
57049	:douta	=	16'h	bbe9;
57050	:douta	=	16'h	bbe9;
57051	:douta	=	16'h	bc09;
57052	:douta	=	16'h	bbe9;
57053	:douta	=	16'h	bbe9;
57054	:douta	=	16'h	bbe9;
57055	:douta	=	16'h	b3e8;
57056	:douta	=	16'h	b3e8;
57057	:douta	=	16'h	b3e8;
57058	:douta	=	16'h	b3e8;
57059	:douta	=	16'h	b3e8;
57060	:douta	=	16'h	b3c8;
57061	:douta	=	16'h	b3e8;
57062	:douta	=	16'h	b3a8;
57063	:douta	=	16'h	b3a8;
57064	:douta	=	16'h	b3c8;
57065	:douta	=	16'h	b3a9;
57066	:douta	=	16'h	b3a9;
57067	:douta	=	16'h	b3a9;
57068	:douta	=	16'h	b3a8;
57069	:douta	=	16'h	b3c8;
57070	:douta	=	16'h	b3c8;
57071	:douta	=	16'h	aba8;
57072	:douta	=	16'h	b3a8;
57073	:douta	=	16'h	aba9;
57074	:douta	=	16'h	aba9;
57075	:douta	=	16'h	ab88;
57076	:douta	=	16'h	ab89;
57077	:douta	=	16'h	ab88;
57078	:douta	=	16'h	ab89;
57079	:douta	=	16'h	ab88;
57080	:douta	=	16'h	ab89;
57081	:douta	=	16'h	ab88;
57082	:douta	=	16'h	ab89;
57083	:douta	=	16'h	ab88;
57084	:douta	=	16'h	a389;
57085	:douta	=	16'h	a368;
57086	:douta	=	16'h	a388;
57087	:douta	=	16'h	a388;
57088	:douta	=	16'h	a4f5;
57089	:douta	=	16'h	a4f5;
57090	:douta	=	16'h	9cb4;
57091	:douta	=	16'h	bd75;
57092	:douta	=	16'h	94b5;
57093	:douta	=	16'h	8c95;
57094	:douta	=	16'h	8cb7;
57095	:douta	=	16'h	7c53;
57096	:douta	=	16'h	28e2;
57097	:douta	=	16'h	28e3;
57098	:douta	=	16'h	28e3;
57099	:douta	=	16'h	28e3;
57100	:douta	=	16'h	28e3;
57101	:douta	=	16'h	28e3;
57102	:douta	=	16'h	28e3;
57103	:douta	=	16'h	28e3;
57104	:douta	=	16'h	28e3;
57105	:douta	=	16'h	20c3;
57106	:douta	=	16'h	20c3;
57107	:douta	=	16'h	20c3;
57108	:douta	=	16'h	20a3;
57109	:douta	=	16'h	20c3;
57110	:douta	=	16'h	20c3;
57111	:douta	=	16'h	20a2;
57112	:douta	=	16'h	20a2;
57113	:douta	=	16'h	20a2;
57114	:douta	=	16'h	20c2;
57115	:douta	=	16'h	20c2;
57116	:douta	=	16'h	20c2;
57117	:douta	=	16'h	28c3;
57118	:douta	=	16'h	28e3;
57119	:douta	=	16'h	28e3;
57120	:douta	=	16'h	30e3;
57121	:douta	=	16'h	28e2;
57122	:douta	=	16'h	30e2;
57123	:douta	=	16'h	3103;
57124	:douta	=	16'h	3103;
57125	:douta	=	16'h	3923;
57126	:douta	=	16'h	3923;
57127	:douta	=	16'h	4144;
57128	:douta	=	16'h	4143;
57129	:douta	=	16'h	4984;
57130	:douta	=	16'h	4143;
57131	:douta	=	16'h	528b;
57132	:douta	=	16'h	10c5;
57133	:douta	=	16'h	18c4;
57134	:douta	=	16'h	59c4;
57135	:douta	=	16'h	59c4;
57136	:douta	=	16'h	59c4;
57137	:douta	=	16'h	61e4;
57138	:douta	=	16'h	61e4;
57139	:douta	=	16'h	6204;
57140	:douta	=	16'h	6a04;
57141	:douta	=	16'h	6a25;
57142	:douta	=	16'h	6a24;
57143	:douta	=	16'h	7203;
57144	:douta	=	16'h	9cb0;
57145	:douta	=	16'h	accf;
57146	:douta	=	16'h	7a44;
57147	:douta	=	16'h	7a84;
57148	:douta	=	16'h	7a85;
57149	:douta	=	16'h	8285;
57150	:douta	=	16'h	7a85;
57151	:douta	=	16'h	8aa6;
57152	:douta	=	16'h	8aa5;
57153	:douta	=	16'h	8aa5;
57154	:douta	=	16'h	8ac6;
57155	:douta	=	16'h	8ac6;
57156	:douta	=	16'h	8ac6;
57157	:douta	=	16'h	8ac6;
57158	:douta	=	16'h	8ac6;
57159	:douta	=	16'h	9307;
57160	:douta	=	16'h	9306;
57161	:douta	=	16'h	82a6;
57162	:douta	=	16'h	9b26;
57163	:douta	=	16'h	9b47;
57164	:douta	=	16'h	9b27;
57165	:douta	=	16'h	9b47;
57166	:douta	=	16'h	92e5;
57167	:douta	=	16'h	9326;
57168	:douta	=	16'h	9327;
57169	:douta	=	16'h	a367;
57170	:douta	=	16'h	ab87;
57171	:douta	=	16'h	ab86;
57172	:douta	=	16'h	b3a7;
57173	:douta	=	16'h	b3c7;
57174	:douta	=	16'h	b3c6;
57175	:douta	=	16'h	b3c7;
57176	:douta	=	16'h	b3c7;
57177	:douta	=	16'h	bbe7;
57178	:douta	=	16'h	bbe7;
57179	:douta	=	16'h	bbe7;
57180	:douta	=	16'h	bc07;
57181	:douta	=	16'h	bc07;
57182	:douta	=	16'h	c407;
57183	:douta	=	16'h	bc07;
57184	:douta	=	16'h	c407;
57185	:douta	=	16'h	c428;
57186	:douta	=	16'h	c428;
57187	:douta	=	16'h	c427;
57188	:douta	=	16'h	c428;
57189	:douta	=	16'h	c428;
57190	:douta	=	16'h	c428;
57191	:douta	=	16'h	c448;
57192	:douta	=	16'h	c448;
57193	:douta	=	16'h	cc48;
57194	:douta	=	16'h	cc47;
57195	:douta	=	16'h	c447;
57196	:douta	=	16'h	cc67;
57197	:douta	=	16'h	cc48;
57198	:douta	=	16'h	cc48;
57199	:douta	=	16'h	cc67;
57200	:douta	=	16'h	cc47;
57201	:douta	=	16'h	cc68;
57202	:douta	=	16'h	cc67;
57203	:douta	=	16'h	cc68;
57204	:douta	=	16'h	cc47;
57205	:douta	=	16'h	cc68;
57206	:douta	=	16'h	cc67;
57207	:douta	=	16'h	cc68;
57208	:douta	=	16'h	cc68;
57209	:douta	=	16'h	cc68;
57210	:douta	=	16'h	cc68;
57211	:douta	=	16'h	cc68;
57212	:douta	=	16'h	cc68;
57213	:douta	=	16'h	cc68;
57214	:douta	=	16'h	cc68;
57215	:douta	=	16'h	cc68;
57216	:douta	=	16'h	cc68;
57217	:douta	=	16'h	cc68;
57218	:douta	=	16'h	cc88;
57219	:douta	=	16'h	cc68;
57220	:douta	=	16'h	cc68;
57221	:douta	=	16'h	cc89;
57222	:douta	=	16'h	cc69;
57223	:douta	=	16'h	d489;
57224	:douta	=	16'h	cc89;
57225	:douta	=	16'h	cc89;
57226	:douta	=	16'h	cc89;
57227	:douta	=	16'h	d489;
57228	:douta	=	16'h	d489;
57229	:douta	=	16'h	cc89;
57230	:douta	=	16'h	cc89;
57231	:douta	=	16'h	d48a;
57232	:douta	=	16'h	d489;
57233	:douta	=	16'h	d489;
57234	:douta	=	16'h	cc89;
57235	:douta	=	16'h	d489;
57236	:douta	=	16'h	d489;
57237	:douta	=	16'h	cc89;
57238	:douta	=	16'h	cc89;
57239	:douta	=	16'h	cc69;
57240	:douta	=	16'h	cc89;
57241	:douta	=	16'h	d48a;
57242	:douta	=	16'h	cc8a;
57243	:douta	=	16'h	cc89;
57244	:douta	=	16'h	d489;
57245	:douta	=	16'h	cc89;
57246	:douta	=	16'h	cc89;
57247	:douta	=	16'h	cc89;
57248	:douta	=	16'h	d489;
57249	:douta	=	16'h	cc69;
57250	:douta	=	16'h	d468;
57251	:douta	=	16'h	ad33;
57252	:douta	=	16'h	e6b7;
57253	:douta	=	16'h	cc47;
57254	:douta	=	16'h	cc69;
57255	:douta	=	16'h	cc89;
57256	:douta	=	16'h	cc69;
57257	:douta	=	16'h	cc69;
57258	:douta	=	16'h	cc69;
57259	:douta	=	16'h	cc69;
57260	:douta	=	16'h	cc89;
57261	:douta	=	16'h	cc89;
57262	:douta	=	16'h	cc69;
57263	:douta	=	16'h	cc69;
57264	:douta	=	16'h	cc69;
57265	:douta	=	16'h	cc69;
57266	:douta	=	16'h	cc69;
57267	:douta	=	16'h	cc69;
57268	:douta	=	16'h	c468;
57269	:douta	=	16'h	cc69;
57270	:douta	=	16'h	d447;
57271	:douta	=	16'h	c449;
57272	:douta	=	16'h	cc48;
57273	:douta	=	16'h	cc49;
57274	:douta	=	16'h	d468;
57275	:douta	=	16'h	d485;
57276	:douta	=	16'h	cc6b;
57277	:douta	=	16'h	d618;
57278	:douta	=	16'h	bc4b;
57279	:douta	=	16'h	c428;
57280	:douta	=	16'h	c3a3;
57281	:douta	=	16'h	c448;
57282	:douta	=	16'h	cc49;
57283	:douta	=	16'h	cc4a;
57284	:douta	=	16'h	c449;
57285	:douta	=	16'h	cc49;
57286	:douta	=	16'h	c449;
57287	:douta	=	16'h	c448;
57288	:douta	=	16'h	c428;
57289	:douta	=	16'h	c428;
57290	:douta	=	16'h	c428;
57291	:douta	=	16'h	c449;
57292	:douta	=	16'h	c449;
57293	:douta	=	16'h	c429;
57294	:douta	=	16'h	c429;
57295	:douta	=	16'h	bc08;
57296	:douta	=	16'h	c429;
57297	:douta	=	16'h	c429;
57298	:douta	=	16'h	c429;
57299	:douta	=	16'h	bc09;
57300	:douta	=	16'h	bc09;
57301	:douta	=	16'h	bc09;
57302	:douta	=	16'h	bc09;
57303	:douta	=	16'h	bc09;
57304	:douta	=	16'h	bc09;
57305	:douta	=	16'h	bc09;
57306	:douta	=	16'h	bc09;
57307	:douta	=	16'h	bbe9;
57308	:douta	=	16'h	bbe9;
57309	:douta	=	16'h	b3c8;
57310	:douta	=	16'h	bbe9;
57311	:douta	=	16'h	b3e9;
57312	:douta	=	16'h	b3e9;
57313	:douta	=	16'h	b3c9;
57314	:douta	=	16'h	b3c9;
57315	:douta	=	16'h	b3c8;
57316	:douta	=	16'h	b3c9;
57317	:douta	=	16'h	b3c8;
57318	:douta	=	16'h	b3c9;
57319	:douta	=	16'h	b3c8;
57320	:douta	=	16'h	b3a8;
57321	:douta	=	16'h	b3c8;
57322	:douta	=	16'h	b3a8;
57323	:douta	=	16'h	b3c8;
57324	:douta	=	16'h	b3c9;
57325	:douta	=	16'h	b3c8;
57326	:douta	=	16'h	b3c8;
57327	:douta	=	16'h	b3a8;
57328	:douta	=	16'h	b3a8;
57329	:douta	=	16'h	ab89;
57330	:douta	=	16'h	ab89;
57331	:douta	=	16'h	aba9;
57332	:douta	=	16'h	ab89;
57333	:douta	=	16'h	aba9;
57334	:douta	=	16'h	aba9;
57335	:douta	=	16'h	aba8;
57336	:douta	=	16'h	aba8;
57337	:douta	=	16'h	aba8;
57338	:douta	=	16'h	aba8;
57339	:douta	=	16'h	a388;
57340	:douta	=	16'h	a388;
57341	:douta	=	16'h	a389;
57342	:douta	=	16'h	a388;
57343	:douta	=	16'h	a389;
57344	:douta	=	16'h	a4d5;
57345	:douta	=	16'h	a4f5;
57346	:douta	=	16'h	9cd4;
57347	:douta	=	16'h	b555;
57348	:douta	=	16'h	8c95;
57349	:douta	=	16'h	8c95;
57350	:douta	=	16'h	94f7;
57351	:douta	=	16'h	636f;
57352	:douta	=	16'h	28e3;
57353	:douta	=	16'h	28e3;
57354	:douta	=	16'h	28e3;
57355	:douta	=	16'h	28e3;
57356	:douta	=	16'h	28e3;
57357	:douta	=	16'h	28e3;
57358	:douta	=	16'h	28e3;
57359	:douta	=	16'h	28e3;
57360	:douta	=	16'h	28e3;
57361	:douta	=	16'h	28e3;
57362	:douta	=	16'h	20c3;
57363	:douta	=	16'h	20c3;
57364	:douta	=	16'h	20a3;
57365	:douta	=	16'h	20e3;
57366	:douta	=	16'h	20c3;
57367	:douta	=	16'h	20a2;
57368	:douta	=	16'h	20c2;
57369	:douta	=	16'h	20a2;
57370	:douta	=	16'h	20c2;
57371	:douta	=	16'h	20c2;
57372	:douta	=	16'h	28c3;
57373	:douta	=	16'h	28e3;
57374	:douta	=	16'h	28e2;
57375	:douta	=	16'h	28e3;
57376	:douta	=	16'h	30e3;
57377	:douta	=	16'h	28e3;
57378	:douta	=	16'h	3103;
57379	:douta	=	16'h	3103;
57380	:douta	=	16'h	3123;
57381	:douta	=	16'h	3103;
57382	:douta	=	16'h	3944;
57383	:douta	=	16'h	4124;
57384	:douta	=	16'h	4164;
57385	:douta	=	16'h	4984;
57386	:douta	=	16'h	4964;
57387	:douta	=	16'h	528b;
57388	:douta	=	16'h	10c5;
57389	:douta	=	16'h	20e4;
57390	:douta	=	16'h	59c4;
57391	:douta	=	16'h	59c4;
57392	:douta	=	16'h	61c4;
57393	:douta	=	16'h	61e4;
57394	:douta	=	16'h	61e4;
57395	:douta	=	16'h	6204;
57396	:douta	=	16'h	6a24;
57397	:douta	=	16'h	6a24;
57398	:douta	=	16'h	7224;
57399	:douta	=	16'h	6a03;
57400	:douta	=	16'h	a511;
57401	:douta	=	16'h	a48d;
57402	:douta	=	16'h	7a64;
57403	:douta	=	16'h	7a84;
57404	:douta	=	16'h	7a85;
57405	:douta	=	16'h	82a5;
57406	:douta	=	16'h	82a5;
57407	:douta	=	16'h	8aa6;
57408	:douta	=	16'h	8aa5;
57409	:douta	=	16'h	8ac6;
57410	:douta	=	16'h	8ac6;
57411	:douta	=	16'h	8ac5;
57412	:douta	=	16'h	8ac6;
57413	:douta	=	16'h	8ae6;
57414	:douta	=	16'h	8ac6;
57415	:douta	=	16'h	9306;
57416	:douta	=	16'h	9306;
57417	:douta	=	16'h	8ac6;
57418	:douta	=	16'h	9306;
57419	:douta	=	16'h	9b46;
57420	:douta	=	16'h	9326;
57421	:douta	=	16'h	9b47;
57422	:douta	=	16'h	9306;
57423	:douta	=	16'h	9307;
57424	:douta	=	16'h	9326;
57425	:douta	=	16'h	a367;
57426	:douta	=	16'h	ab87;
57427	:douta	=	16'h	aba7;
57428	:douta	=	16'h	aba7;
57429	:douta	=	16'h	b3c7;
57430	:douta	=	16'h	b3c6;
57431	:douta	=	16'h	b3c7;
57432	:douta	=	16'h	b3e6;
57433	:douta	=	16'h	bbe7;
57434	:douta	=	16'h	bbe7;
57435	:douta	=	16'h	bc07;
57436	:douta	=	16'h	bbe7;
57437	:douta	=	16'h	bbe7;
57438	:douta	=	16'h	bc07;
57439	:douta	=	16'h	bc07;
57440	:douta	=	16'h	bc07;
57441	:douta	=	16'h	bc07;
57442	:douta	=	16'h	c448;
57443	:douta	=	16'h	c427;
57444	:douta	=	16'h	c428;
57445	:douta	=	16'h	c448;
57446	:douta	=	16'h	c448;
57447	:douta	=	16'h	c448;
57448	:douta	=	16'h	c428;
57449	:douta	=	16'h	cc48;
57450	:douta	=	16'h	c447;
57451	:douta	=	16'h	cc47;
57452	:douta	=	16'h	cc48;
57453	:douta	=	16'h	cc48;
57454	:douta	=	16'h	cc48;
57455	:douta	=	16'h	cc68;
57456	:douta	=	16'h	cc67;
57457	:douta	=	16'h	cc67;
57458	:douta	=	16'h	cc47;
57459	:douta	=	16'h	cc67;
57460	:douta	=	16'h	cc68;
57461	:douta	=	16'h	cc67;
57462	:douta	=	16'h	cc68;
57463	:douta	=	16'h	cc68;
57464	:douta	=	16'h	cc68;
57465	:douta	=	16'h	cc68;
57466	:douta	=	16'h	cc68;
57467	:douta	=	16'h	cc68;
57468	:douta	=	16'h	cc68;
57469	:douta	=	16'h	cc68;
57470	:douta	=	16'h	cc88;
57471	:douta	=	16'h	cc88;
57472	:douta	=	16'h	cc68;
57473	:douta	=	16'h	cc68;
57474	:douta	=	16'h	cc68;
57475	:douta	=	16'h	cc88;
57476	:douta	=	16'h	cc88;
57477	:douta	=	16'h	cc89;
57478	:douta	=	16'h	cc68;
57479	:douta	=	16'h	cc89;
57480	:douta	=	16'h	cc89;
57481	:douta	=	16'h	cc89;
57482	:douta	=	16'h	cc89;
57483	:douta	=	16'h	d489;
57484	:douta	=	16'h	cc89;
57485	:douta	=	16'h	cc69;
57486	:douta	=	16'h	cc89;
57487	:douta	=	16'h	d489;
57488	:douta	=	16'h	cc69;
57489	:douta	=	16'h	d489;
57490	:douta	=	16'h	cc89;
57491	:douta	=	16'h	cc69;
57492	:douta	=	16'h	cc89;
57493	:douta	=	16'h	cc89;
57494	:douta	=	16'h	cc89;
57495	:douta	=	16'h	cc89;
57496	:douta	=	16'h	cc89;
57497	:douta	=	16'h	cc89;
57498	:douta	=	16'h	cc8a;
57499	:douta	=	16'h	cc69;
57500	:douta	=	16'h	d489;
57501	:douta	=	16'h	cc69;
57502	:douta	=	16'h	cc89;
57503	:douta	=	16'h	cc89;
57504	:douta	=	16'h	cc88;
57505	:douta	=	16'h	cc69;
57506	:douta	=	16'h	d468;
57507	:douta	=	16'h	ad53;
57508	:douta	=	16'h	de96;
57509	:douta	=	16'h	cc47;
57510	:douta	=	16'h	cc68;
57511	:douta	=	16'h	cc69;
57512	:douta	=	16'h	cc69;
57513	:douta	=	16'h	cc69;
57514	:douta	=	16'h	cc69;
57515	:douta	=	16'h	cc69;
57516	:douta	=	16'h	cc69;
57517	:douta	=	16'h	cc69;
57518	:douta	=	16'h	cc69;
57519	:douta	=	16'h	cc89;
57520	:douta	=	16'h	cc69;
57521	:douta	=	16'h	cc69;
57522	:douta	=	16'h	cc69;
57523	:douta	=	16'h	cc69;
57524	:douta	=	16'h	cc69;
57525	:douta	=	16'h	cc68;
57526	:douta	=	16'h	cc69;
57527	:douta	=	16'h	cc48;
57528	:douta	=	16'h	cc69;
57529	:douta	=	16'h	cc69;
57530	:douta	=	16'h	cc69;
57531	:douta	=	16'h	cc49;
57532	:douta	=	16'h	cc68;
57533	:douta	=	16'h	c3c3;
57534	:douta	=	16'h	d447;
57535	:douta	=	16'h	cc68;
57536	:douta	=	16'h	cc49;
57537	:douta	=	16'h	c449;
57538	:douta	=	16'h	c449;
57539	:douta	=	16'h	c448;
57540	:douta	=	16'h	c448;
57541	:douta	=	16'h	c449;
57542	:douta	=	16'h	cc29;
57543	:douta	=	16'h	c448;
57544	:douta	=	16'h	c428;
57545	:douta	=	16'h	c428;
57546	:douta	=	16'h	c428;
57547	:douta	=	16'h	c429;
57548	:douta	=	16'h	c429;
57549	:douta	=	16'h	c429;
57550	:douta	=	16'h	c429;
57551	:douta	=	16'h	bc08;
57552	:douta	=	16'h	c429;
57553	:douta	=	16'h	c429;
57554	:douta	=	16'h	c429;
57555	:douta	=	16'h	bc09;
57556	:douta	=	16'h	bc08;
57557	:douta	=	16'h	bc09;
57558	:douta	=	16'h	bc09;
57559	:douta	=	16'h	bc09;
57560	:douta	=	16'h	bc09;
57561	:douta	=	16'h	bc09;
57562	:douta	=	16'h	bbe9;
57563	:douta	=	16'h	bbe9;
57564	:douta	=	16'h	b3c9;
57565	:douta	=	16'h	bbe9;
57566	:douta	=	16'h	b3e8;
57567	:douta	=	16'h	b3e9;
57568	:douta	=	16'h	b3e9;
57569	:douta	=	16'h	b3c9;
57570	:douta	=	16'h	b3e9;
57571	:douta	=	16'h	b3c9;
57572	:douta	=	16'h	b3c8;
57573	:douta	=	16'h	b3c8;
57574	:douta	=	16'h	b3c8;
57575	:douta	=	16'h	b3c8;
57576	:douta	=	16'h	b3a8;
57577	:douta	=	16'h	b3c9;
57578	:douta	=	16'h	b3a8;
57579	:douta	=	16'h	b3a8;
57580	:douta	=	16'h	b3c8;
57581	:douta	=	16'h	b3a8;
57582	:douta	=	16'h	aba9;
57583	:douta	=	16'h	b3a8;
57584	:douta	=	16'h	b3c8;
57585	:douta	=	16'h	aba9;
57586	:douta	=	16'h	aba9;
57587	:douta	=	16'h	aba9;
57588	:douta	=	16'h	aba9;
57589	:douta	=	16'h	ab88;
57590	:douta	=	16'h	aba9;
57591	:douta	=	16'h	aba8;
57592	:douta	=	16'h	aba8;
57593	:douta	=	16'h	a388;
57594	:douta	=	16'h	a388;
57595	:douta	=	16'h	a388;
57596	:douta	=	16'h	a388;
57597	:douta	=	16'h	a388;
57598	:douta	=	16'h	a368;
57599	:douta	=	16'h	a368;
57600	:douta	=	16'h	a4f5;
57601	:douta	=	16'h	a4d5;
57602	:douta	=	16'h	a4d4;
57603	:douta	=	16'h	a515;
57604	:douta	=	16'h	8cb6;
57605	:douta	=	16'h	94b6;
57606	:douta	=	16'h	8495;
57607	:douta	=	16'h	3186;
57608	:douta	=	16'h	2903;
57609	:douta	=	16'h	28e3;
57610	:douta	=	16'h	28e3;
57611	:douta	=	16'h	28e3;
57612	:douta	=	16'h	28e3;
57613	:douta	=	16'h	28e3;
57614	:douta	=	16'h	20c3;
57615	:douta	=	16'h	28e3;
57616	:douta	=	16'h	28e3;
57617	:douta	=	16'h	28e3;
57618	:douta	=	16'h	20c3;
57619	:douta	=	16'h	20a3;
57620	:douta	=	16'h	20c3;
57621	:douta	=	16'h	20e3;
57622	:douta	=	16'h	20e3;
57623	:douta	=	16'h	20a2;
57624	:douta	=	16'h	1881;
57625	:douta	=	16'h	20c2;
57626	:douta	=	16'h	20a2;
57627	:douta	=	16'h	20a2;
57628	:douta	=	16'h	28e3;
57629	:douta	=	16'h	28e3;
57630	:douta	=	16'h	28e3;
57631	:douta	=	16'h	30e3;
57632	:douta	=	16'h	28e3;
57633	:douta	=	16'h	30e3;
57634	:douta	=	16'h	3103;
57635	:douta	=	16'h	3103;
57636	:douta	=	16'h	3923;
57637	:douta	=	16'h	3923;
57638	:douta	=	16'h	4123;
57639	:douta	=	16'h	4144;
57640	:douta	=	16'h	4143;
57641	:douta	=	16'h	4963;
57642	:douta	=	16'h	4964;
57643	:douta	=	16'h	4a49;
57644	:douta	=	16'h	10a5;
57645	:douta	=	16'h	3924;
57646	:douta	=	16'h	51a4;
57647	:douta	=	16'h	59c4;
57648	:douta	=	16'h	59c4;
57649	:douta	=	16'h	61e4;
57650	:douta	=	16'h	61e4;
57651	:douta	=	16'h	6a24;
57652	:douta	=	16'h	6a04;
57653	:douta	=	16'h	6a24;
57654	:douta	=	16'h	7224;
57655	:douta	=	16'h	7245;
57656	:douta	=	16'h	b592;
57657	:douta	=	16'h	93aa;
57658	:douta	=	16'h	7a64;
57659	:douta	=	16'h	7a85;
57660	:douta	=	16'h	7a85;
57661	:douta	=	16'h	7a85;
57662	:douta	=	16'h	8285;
57663	:douta	=	16'h	8aa6;
57664	:douta	=	16'h	82c5;
57665	:douta	=	16'h	8ac6;
57666	:douta	=	16'h	8ac6;
57667	:douta	=	16'h	8ac6;
57668	:douta	=	16'h	8ac6;
57669	:douta	=	16'h	8ac6;
57670	:douta	=	16'h	8ac6;
57671	:douta	=	16'h	9306;
57672	:douta	=	16'h	9306;
57673	:douta	=	16'h	9b47;
57674	:douta	=	16'h	7a85;
57675	:douta	=	16'h	a347;
57676	:douta	=	16'h	9b47;
57677	:douta	=	16'h	9b47;
57678	:douta	=	16'h	9306;
57679	:douta	=	16'h	9b47;
57680	:douta	=	16'h	9b47;
57681	:douta	=	16'h	a367;
57682	:douta	=	16'h	ab87;
57683	:douta	=	16'h	aba7;
57684	:douta	=	16'h	b3a7;
57685	:douta	=	16'h	b3c7;
57686	:douta	=	16'h	b3c7;
57687	:douta	=	16'h	bbe7;
57688	:douta	=	16'h	bbe7;
57689	:douta	=	16'h	bbe7;
57690	:douta	=	16'h	bbe7;
57691	:douta	=	16'h	bbe7;
57692	:douta	=	16'h	bbe7;
57693	:douta	=	16'h	bc07;
57694	:douta	=	16'h	bc08;
57695	:douta	=	16'h	c407;
57696	:douta	=	16'h	bc07;
57697	:douta	=	16'h	c428;
57698	:douta	=	16'h	c428;
57699	:douta	=	16'h	c428;
57700	:douta	=	16'h	c428;
57701	:douta	=	16'h	c428;
57702	:douta	=	16'h	c448;
57703	:douta	=	16'h	c448;
57704	:douta	=	16'h	c448;
57705	:douta	=	16'h	cc67;
57706	:douta	=	16'h	cc47;
57707	:douta	=	16'h	cc47;
57708	:douta	=	16'h	cc48;
57709	:douta	=	16'h	cc48;
57710	:douta	=	16'h	cc67;
57711	:douta	=	16'h	cc68;
57712	:douta	=	16'h	cc67;
57713	:douta	=	16'h	cc68;
57714	:douta	=	16'h	cc67;
57715	:douta	=	16'h	cc68;
57716	:douta	=	16'h	cc47;
57717	:douta	=	16'h	cc68;
57718	:douta	=	16'h	cc67;
57719	:douta	=	16'h	cc68;
57720	:douta	=	16'h	cc68;
57721	:douta	=	16'h	cc68;
57722	:douta	=	16'h	cc68;
57723	:douta	=	16'h	cc88;
57724	:douta	=	16'h	cc68;
57725	:douta	=	16'h	cc88;
57726	:douta	=	16'h	cc68;
57727	:douta	=	16'h	cc68;
57728	:douta	=	16'h	cc88;
57729	:douta	=	16'h	cc88;
57730	:douta	=	16'h	cc88;
57731	:douta	=	16'h	cc68;
57732	:douta	=	16'h	cc68;
57733	:douta	=	16'h	cc69;
57734	:douta	=	16'h	cc68;
57735	:douta	=	16'h	cc69;
57736	:douta	=	16'h	cc89;
57737	:douta	=	16'h	cc89;
57738	:douta	=	16'h	cc89;
57739	:douta	=	16'h	cc89;
57740	:douta	=	16'h	d489;
57741	:douta	=	16'h	cc69;
57742	:douta	=	16'h	cc69;
57743	:douta	=	16'h	cc69;
57744	:douta	=	16'h	d489;
57745	:douta	=	16'h	cc89;
57746	:douta	=	16'h	d489;
57747	:douta	=	16'h	cc89;
57748	:douta	=	16'h	d489;
57749	:douta	=	16'h	d489;
57750	:douta	=	16'h	cc89;
57751	:douta	=	16'h	cc69;
57752	:douta	=	16'h	cc89;
57753	:douta	=	16'h	d48a;
57754	:douta	=	16'h	cc89;
57755	:douta	=	16'h	cc89;
57756	:douta	=	16'h	cc8a;
57757	:douta	=	16'h	cc89;
57758	:douta	=	16'h	cc89;
57759	:douta	=	16'h	cc69;
57760	:douta	=	16'h	cc88;
57761	:douta	=	16'h	cc89;
57762	:douta	=	16'h	d468;
57763	:douta	=	16'h	ad53;
57764	:douta	=	16'h	e6b7;
57765	:douta	=	16'h	cc27;
57766	:douta	=	16'h	cc89;
57767	:douta	=	16'h	cc69;
57768	:douta	=	16'h	cc69;
57769	:douta	=	16'h	cc89;
57770	:douta	=	16'h	cc69;
57771	:douta	=	16'h	cc69;
57772	:douta	=	16'h	cc69;
57773	:douta	=	16'h	cc69;
57774	:douta	=	16'h	cc69;
57775	:douta	=	16'h	cc69;
57776	:douta	=	16'h	cc69;
57777	:douta	=	16'h	cc69;
57778	:douta	=	16'h	cc69;
57779	:douta	=	16'h	cc49;
57780	:douta	=	16'h	cc48;
57781	:douta	=	16'h	cc69;
57782	:douta	=	16'h	cc69;
57783	:douta	=	16'h	cc49;
57784	:douta	=	16'h	cc68;
57785	:douta	=	16'h	cc69;
57786	:douta	=	16'h	cc49;
57787	:douta	=	16'h	cc69;
57788	:douta	=	16'h	cc48;
57789	:douta	=	16'h	cc69;
57790	:douta	=	16'h	cc49;
57791	:douta	=	16'h	cc49;
57792	:douta	=	16'h	cc49;
57793	:douta	=	16'h	c449;
57794	:douta	=	16'h	c429;
57795	:douta	=	16'h	cc49;
57796	:douta	=	16'h	cc49;
57797	:douta	=	16'h	cc49;
57798	:douta	=	16'h	c448;
57799	:douta	=	16'h	c428;
57800	:douta	=	16'h	c428;
57801	:douta	=	16'h	c449;
57802	:douta	=	16'h	c449;
57803	:douta	=	16'h	c429;
57804	:douta	=	16'h	c449;
57805	:douta	=	16'h	c429;
57806	:douta	=	16'h	c429;
57807	:douta	=	16'h	c429;
57808	:douta	=	16'h	c429;
57809	:douta	=	16'h	c429;
57810	:douta	=	16'h	bc09;
57811	:douta	=	16'h	c429;
57812	:douta	=	16'h	bc08;
57813	:douta	=	16'h	bc09;
57814	:douta	=	16'h	bc09;
57815	:douta	=	16'h	bc09;
57816	:douta	=	16'h	bbe8;
57817	:douta	=	16'h	bc09;
57818	:douta	=	16'h	b3e8;
57819	:douta	=	16'h	b3e8;
57820	:douta	=	16'h	bbe9;
57821	:douta	=	16'h	bbe9;
57822	:douta	=	16'h	bbe9;
57823	:douta	=	16'h	bbe9;
57824	:douta	=	16'h	b3c9;
57825	:douta	=	16'h	b3e9;
57826	:douta	=	16'h	b3e9;
57827	:douta	=	16'h	b3c8;
57828	:douta	=	16'h	b3c8;
57829	:douta	=	16'h	b3c8;
57830	:douta	=	16'h	b3c8;
57831	:douta	=	16'h	b3c8;
57832	:douta	=	16'h	b3c8;
57833	:douta	=	16'h	b3c8;
57834	:douta	=	16'h	b3c8;
57835	:douta	=	16'h	b3c9;
57836	:douta	=	16'h	b3c9;
57837	:douta	=	16'h	b3c8;
57838	:douta	=	16'h	aba9;
57839	:douta	=	16'h	b3a9;
57840	:douta	=	16'h	aba9;
57841	:douta	=	16'h	aba9;
57842	:douta	=	16'h	aba9;
57843	:douta	=	16'h	aba9;
57844	:douta	=	16'h	ab89;
57845	:douta	=	16'h	abc9;
57846	:douta	=	16'h	aba9;
57847	:douta	=	16'h	ab88;
57848	:douta	=	16'h	ab89;
57849	:douta	=	16'h	ab89;
57850	:douta	=	16'h	a389;
57851	:douta	=	16'h	a368;
57852	:douta	=	16'h	a368;
57853	:douta	=	16'h	a389;
57854	:douta	=	16'h	a368;
57855	:douta	=	16'h	a388;
57856	:douta	=	16'h	a4f5;
57857	:douta	=	16'h	a4d5;
57858	:douta	=	16'h	a4d4;
57859	:douta	=	16'h	9cf5;
57860	:douta	=	16'h	94d6;
57861	:douta	=	16'h	8cb5;
57862	:douta	=	16'h	73b1;
57863	:douta	=	16'h	1881;
57864	:douta	=	16'h	2903;
57865	:douta	=	16'h	28e3;
57866	:douta	=	16'h	28e3;
57867	:douta	=	16'h	28e3;
57868	:douta	=	16'h	28e3;
57869	:douta	=	16'h	28e3;
57870	:douta	=	16'h	28e3;
57871	:douta	=	16'h	20c3;
57872	:douta	=	16'h	20c3;
57873	:douta	=	16'h	20c3;
57874	:douta	=	16'h	20c3;
57875	:douta	=	16'h	20c3;
57876	:douta	=	16'h	20c3;
57877	:douta	=	16'h	20e3;
57878	:douta	=	16'h	20a2;
57879	:douta	=	16'h	20a2;
57880	:douta	=	16'h	20c2;
57881	:douta	=	16'h	20c2;
57882	:douta	=	16'h	20a2;
57883	:douta	=	16'h	20a2;
57884	:douta	=	16'h	28c3;
57885	:douta	=	16'h	28e3;
57886	:douta	=	16'h	28e3;
57887	:douta	=	16'h	3103;
57888	:douta	=	16'h	3103;
57889	:douta	=	16'h	30e3;
57890	:douta	=	16'h	3103;
57891	:douta	=	16'h	3103;
57892	:douta	=	16'h	3923;
57893	:douta	=	16'h	4144;
57894	:douta	=	16'h	4144;
57895	:douta	=	16'h	4163;
57896	:douta	=	16'h	4964;
57897	:douta	=	16'h	4963;
57898	:douta	=	16'h	4985;
57899	:douta	=	16'h	4209;
57900	:douta	=	16'h	10c5;
57901	:douta	=	16'h	4964;
57902	:douta	=	16'h	59a4;
57903	:douta	=	16'h	59c4;
57904	:douta	=	16'h	61e4;
57905	:douta	=	16'h	6204;
57906	:douta	=	16'h	6204;
57907	:douta	=	16'h	6a04;
57908	:douta	=	16'h	6a04;
57909	:douta	=	16'h	6a24;
57910	:douta	=	16'h	6a24;
57911	:douta	=	16'h	7246;
57912	:douta	=	16'h	b572;
57913	:douta	=	16'h	8b28;
57914	:douta	=	16'h	7a64;
57915	:douta	=	16'h	7a85;
57916	:douta	=	16'h	7a85;
57917	:douta	=	16'h	7a85;
57918	:douta	=	16'h	82a5;
57919	:douta	=	16'h	82a6;
57920	:douta	=	16'h	8ac6;
57921	:douta	=	16'h	8ac6;
57922	:douta	=	16'h	8ac6;
57923	:douta	=	16'h	8ac6;
57924	:douta	=	16'h	8ac6;
57925	:douta	=	16'h	8ae6;
57926	:douta	=	16'h	8ac6;
57927	:douta	=	16'h	9306;
57928	:douta	=	16'h	9306;
57929	:douta	=	16'h	9b46;
57930	:douta	=	16'h	7266;
57931	:douta	=	16'h	a367;
57932	:douta	=	16'h	9326;
57933	:douta	=	16'h	9b26;
57934	:douta	=	16'h	9305;
57935	:douta	=	16'h	9305;
57936	:douta	=	16'h	9305;
57937	:douta	=	16'h	a346;
57938	:douta	=	16'h	a366;
57939	:douta	=	16'h	aba7;
57940	:douta	=	16'h	ab87;
57941	:douta	=	16'h	abc7;
57942	:douta	=	16'h	b3c7;
57943	:douta	=	16'h	b3c7;
57944	:douta	=	16'h	bbe7;
57945	:douta	=	16'h	bbe7;
57946	:douta	=	16'h	bbe7;
57947	:douta	=	16'h	bc07;
57948	:douta	=	16'h	bbe7;
57949	:douta	=	16'h	bc07;
57950	:douta	=	16'h	bc07;
57951	:douta	=	16'h	bc07;
57952	:douta	=	16'h	c428;
57953	:douta	=	16'h	c428;
57954	:douta	=	16'h	c427;
57955	:douta	=	16'h	c427;
57956	:douta	=	16'h	c427;
57957	:douta	=	16'h	c448;
57958	:douta	=	16'h	c427;
57959	:douta	=	16'h	c448;
57960	:douta	=	16'h	c448;
57961	:douta	=	16'h	cc47;
57962	:douta	=	16'h	cc47;
57963	:douta	=	16'h	c447;
57964	:douta	=	16'h	cc48;
57965	:douta	=	16'h	cc48;
57966	:douta	=	16'h	cc67;
57967	:douta	=	16'h	cc68;
57968	:douta	=	16'h	cc48;
57969	:douta	=	16'h	cc68;
57970	:douta	=	16'h	cc67;
57971	:douta	=	16'h	cc47;
57972	:douta	=	16'h	cc67;
57973	:douta	=	16'h	cc67;
57974	:douta	=	16'h	cc68;
57975	:douta	=	16'h	cc68;
57976	:douta	=	16'h	cc68;
57977	:douta	=	16'h	cc68;
57978	:douta	=	16'h	cc68;
57979	:douta	=	16'h	cc68;
57980	:douta	=	16'h	cc68;
57981	:douta	=	16'h	cc68;
57982	:douta	=	16'h	cc88;
57983	:douta	=	16'h	cc88;
57984	:douta	=	16'h	cc68;
57985	:douta	=	16'h	cc88;
57986	:douta	=	16'h	cc88;
57987	:douta	=	16'h	cc69;
57988	:douta	=	16'h	cc68;
57989	:douta	=	16'h	cc89;
57990	:douta	=	16'h	cc89;
57991	:douta	=	16'h	cc69;
57992	:douta	=	16'h	cc69;
57993	:douta	=	16'h	d489;
57994	:douta	=	16'h	cc89;
57995	:douta	=	16'h	cc69;
57996	:douta	=	16'h	d489;
57997	:douta	=	16'h	cc69;
57998	:douta	=	16'h	cc69;
57999	:douta	=	16'h	d489;
58000	:douta	=	16'h	cc69;
58001	:douta	=	16'h	cc89;
58002	:douta	=	16'h	d48a;
58003	:douta	=	16'h	cc89;
58004	:douta	=	16'h	cc89;
58005	:douta	=	16'h	cc69;
58006	:douta	=	16'h	cc89;
58007	:douta	=	16'h	cc69;
58008	:douta	=	16'h	cc69;
58009	:douta	=	16'h	cc8a;
58010	:douta	=	16'h	cc8a;
58011	:douta	=	16'h	cc89;
58012	:douta	=	16'h	cc8a;
58013	:douta	=	16'h	cc89;
58014	:douta	=	16'h	cc89;
58015	:douta	=	16'h	cc69;
58016	:douta	=	16'h	cc69;
58017	:douta	=	16'h	cc89;
58018	:douta	=	16'h	d468;
58019	:douta	=	16'h	ad73;
58020	:douta	=	16'h	e696;
58021	:douta	=	16'h	cc27;
58022	:douta	=	16'h	cc69;
58023	:douta	=	16'h	cc69;
58024	:douta	=	16'h	cc69;
58025	:douta	=	16'h	cc89;
58026	:douta	=	16'h	cc89;
58027	:douta	=	16'h	cc69;
58028	:douta	=	16'h	cc69;
58029	:douta	=	16'h	cc69;
58030	:douta	=	16'h	cc69;
58031	:douta	=	16'h	cc69;
58032	:douta	=	16'h	cc69;
58033	:douta	=	16'h	cc69;
58034	:douta	=	16'h	cc69;
58035	:douta	=	16'h	cc69;
58036	:douta	=	16'h	cc69;
58037	:douta	=	16'h	cc69;
58038	:douta	=	16'h	cc68;
58039	:douta	=	16'h	cc6a;
58040	:douta	=	16'h	cc69;
58041	:douta	=	16'h	cc49;
58042	:douta	=	16'h	cc49;
58043	:douta	=	16'h	cc69;
58044	:douta	=	16'h	c468;
58045	:douta	=	16'h	cc68;
58046	:douta	=	16'h	c449;
58047	:douta	=	16'h	cc69;
58048	:douta	=	16'h	cc49;
58049	:douta	=	16'h	c468;
58050	:douta	=	16'h	cc49;
58051	:douta	=	16'h	c449;
58052	:douta	=	16'h	c449;
58053	:douta	=	16'h	c449;
58054	:douta	=	16'h	c449;
58055	:douta	=	16'h	c428;
58056	:douta	=	16'h	c428;
58057	:douta	=	16'h	c449;
58058	:douta	=	16'h	c429;
58059	:douta	=	16'h	c429;
58060	:douta	=	16'h	c429;
58061	:douta	=	16'h	c429;
58062	:douta	=	16'h	c429;
58063	:douta	=	16'h	c429;
58064	:douta	=	16'h	bc09;
58065	:douta	=	16'h	bc09;
58066	:douta	=	16'h	c429;
58067	:douta	=	16'h	c429;
58068	:douta	=	16'h	bc08;
58069	:douta	=	16'h	bc09;
58070	:douta	=	16'h	bc09;
58071	:douta	=	16'h	bc29;
58072	:douta	=	16'h	bc09;
58073	:douta	=	16'h	bc09;
58074	:douta	=	16'h	bbe9;
58075	:douta	=	16'h	bc09;
58076	:douta	=	16'h	bbe9;
58077	:douta	=	16'h	bbe9;
58078	:douta	=	16'h	b3e8;
58079	:douta	=	16'h	bc09;
58080	:douta	=	16'h	b3e9;
58081	:douta	=	16'h	b3e9;
58082	:douta	=	16'h	b3e9;
58083	:douta	=	16'h	b3e9;
58084	:douta	=	16'h	b3c8;
58085	:douta	=	16'h	b3c8;
58086	:douta	=	16'h	b3c8;
58087	:douta	=	16'h	b3c9;
58088	:douta	=	16'h	b3c8;
58089	:douta	=	16'h	b3c8;
58090	:douta	=	16'h	b3c8;
58091	:douta	=	16'h	b3c9;
58092	:douta	=	16'h	b3c8;
58093	:douta	=	16'h	b3c8;
58094	:douta	=	16'h	b3c9;
58095	:douta	=	16'h	aba9;
58096	:douta	=	16'h	aba9;
58097	:douta	=	16'h	aba9;
58098	:douta	=	16'h	aba9;
58099	:douta	=	16'h	aba9;
58100	:douta	=	16'h	aba9;
58101	:douta	=	16'h	aba9;
58102	:douta	=	16'h	aba9;
58103	:douta	=	16'h	aba9;
58104	:douta	=	16'h	ab89;
58105	:douta	=	16'h	aba8;
58106	:douta	=	16'h	a388;
58107	:douta	=	16'h	ab89;
58108	:douta	=	16'h	a388;
58109	:douta	=	16'h	a388;
58110	:douta	=	16'h	a389;
58111	:douta	=	16'h	a368;
58112	:douta	=	16'h	a4d5;
58113	:douta	=	16'h	a4f5;
58114	:douta	=	16'h	acf4;
58115	:douta	=	16'h	8c95;
58116	:douta	=	16'h	94d6;
58117	:douta	=	16'h	8c96;
58118	:douta	=	16'h	39a7;
58119	:douta	=	16'h	2082;
58120	:douta	=	16'h	2904;
58121	:douta	=	16'h	28e3;
58122	:douta	=	16'h	28e3;
58123	:douta	=	16'h	28e3;
58124	:douta	=	16'h	28e3;
58125	:douta	=	16'h	28e3;
58126	:douta	=	16'h	28e3;
58127	:douta	=	16'h	28e3;
58128	:douta	=	16'h	28e3;
58129	:douta	=	16'h	28e3;
58130	:douta	=	16'h	28e3;
58131	:douta	=	16'h	20c3;
58132	:douta	=	16'h	20a2;
58133	:douta	=	16'h	20e3;
58134	:douta	=	16'h	2082;
58135	:douta	=	16'h	20c2;
58136	:douta	=	16'h	20a2;
58137	:douta	=	16'h	20a2;
58138	:douta	=	16'h	20c2;
58139	:douta	=	16'h	28c3;
58140	:douta	=	16'h	28c3;
58141	:douta	=	16'h	28e3;
58142	:douta	=	16'h	28e3;
58143	:douta	=	16'h	28e2;
58144	:douta	=	16'h	28e2;
58145	:douta	=	16'h	30e3;
58146	:douta	=	16'h	3103;
58147	:douta	=	16'h	3103;
58148	:douta	=	16'h	3923;
58149	:douta	=	16'h	4123;
58150	:douta	=	16'h	4123;
58151	:douta	=	16'h	4143;
58152	:douta	=	16'h	4143;
58153	:douta	=	16'h	4963;
58154	:douta	=	16'h	41c7;
58155	:douta	=	16'h	31a7;
58156	:douta	=	16'h	20c4;
58157	:douta	=	16'h	5184;
58158	:douta	=	16'h	59c4;
58159	:douta	=	16'h	59c4;
58160	:douta	=	16'h	61c4;
58161	:douta	=	16'h	6204;
58162	:douta	=	16'h	6a24;
58163	:douta	=	16'h	6204;
58164	:douta	=	16'h	6a04;
58165	:douta	=	16'h	6a24;
58166	:douta	=	16'h	7223;
58167	:douta	=	16'h	6a46;
58168	:douta	=	16'h	b550;
58169	:douta	=	16'h	7245;
58170	:douta	=	16'h	7a85;
58171	:douta	=	16'h	7a85;
58172	:douta	=	16'h	7a85;
58173	:douta	=	16'h	8285;
58174	:douta	=	16'h	82a6;
58175	:douta	=	16'h	8aa6;
58176	:douta	=	16'h	8aa6;
58177	:douta	=	16'h	8ac6;
58178	:douta	=	16'h	8ac6;
58179	:douta	=	16'h	8ac6;
58180	:douta	=	16'h	8ac6;
58181	:douta	=	16'h	92e7;
58182	:douta	=	16'h	9307;
58183	:douta	=	16'h	9306;
58184	:douta	=	16'h	9327;
58185	:douta	=	16'h	9b47;
58186	:douta	=	16'h	51e5;
58187	:douta	=	16'h	7265;
58188	:douta	=	16'h	92e4;
58189	:douta	=	16'h	8a82;
58190	:douta	=	16'h	8243;
58191	:douta	=	16'h	7a23;
58192	:douta	=	16'h	7202;
58193	:douta	=	16'h	8aa2;
58194	:douta	=	16'h	92c4;
58195	:douta	=	16'h	aba6;
58196	:douta	=	16'h	b3a7;
58197	:douta	=	16'h	b3c7;
58198	:douta	=	16'h	b3c7;
58199	:douta	=	16'h	b3e7;
58200	:douta	=	16'h	bbe7;
58201	:douta	=	16'h	bbe7;
58202	:douta	=	16'h	bc07;
58203	:douta	=	16'h	bc07;
58204	:douta	=	16'h	bc07;
58205	:douta	=	16'h	bc08;
58206	:douta	=	16'h	bc08;
58207	:douta	=	16'h	c428;
58208	:douta	=	16'h	bc07;
58209	:douta	=	16'h	c428;
58210	:douta	=	16'h	c428;
58211	:douta	=	16'h	c427;
58212	:douta	=	16'h	c448;
58213	:douta	=	16'h	c428;
58214	:douta	=	16'h	c448;
58215	:douta	=	16'h	c448;
58216	:douta	=	16'h	cc48;
58217	:douta	=	16'h	c448;
58218	:douta	=	16'h	c448;
58219	:douta	=	16'h	c448;
58220	:douta	=	16'h	cc48;
58221	:douta	=	16'h	cc48;
58222	:douta	=	16'h	c448;
58223	:douta	=	16'h	cc68;
58224	:douta	=	16'h	cc68;
58225	:douta	=	16'h	cc68;
58226	:douta	=	16'h	cc67;
58227	:douta	=	16'h	cc68;
58228	:douta	=	16'h	cc67;
58229	:douta	=	16'h	cc68;
58230	:douta	=	16'h	cc67;
58231	:douta	=	16'h	cc68;
58232	:douta	=	16'h	cc68;
58233	:douta	=	16'h	cc68;
58234	:douta	=	16'h	cc67;
58235	:douta	=	16'h	cc68;
58236	:douta	=	16'h	cc68;
58237	:douta	=	16'h	cc68;
58238	:douta	=	16'h	cc68;
58239	:douta	=	16'h	cc68;
58240	:douta	=	16'h	cc88;
58241	:douta	=	16'h	cc69;
58242	:douta	=	16'h	cc68;
58243	:douta	=	16'h	cc89;
58244	:douta	=	16'h	cc68;
58245	:douta	=	16'h	cc89;
58246	:douta	=	16'h	cc69;
58247	:douta	=	16'h	cc89;
58248	:douta	=	16'h	cc69;
58249	:douta	=	16'h	cc89;
58250	:douta	=	16'h	cc69;
58251	:douta	=	16'h	cc89;
58252	:douta	=	16'h	cc89;
58253	:douta	=	16'h	cc69;
58254	:douta	=	16'h	cc69;
58255	:douta	=	16'h	cc89;
58256	:douta	=	16'h	cc89;
58257	:douta	=	16'h	cc69;
58258	:douta	=	16'h	cc89;
58259	:douta	=	16'h	cc69;
58260	:douta	=	16'h	cc89;
58261	:douta	=	16'h	d489;
58262	:douta	=	16'h	cc89;
58263	:douta	=	16'h	cc89;
58264	:douta	=	16'h	cc89;
58265	:douta	=	16'h	d48a;
58266	:douta	=	16'h	d489;
58267	:douta	=	16'h	cc69;
58268	:douta	=	16'h	cc89;
58269	:douta	=	16'h	cc89;
58270	:douta	=	16'h	cc89;
58271	:douta	=	16'h	cc89;
58272	:douta	=	16'h	cc69;
58273	:douta	=	16'h	cc89;
58274	:douta	=	16'h	d468;
58275	:douta	=	16'h	ad73;
58276	:douta	=	16'h	e6b7;
58277	:douta	=	16'h	cc47;
58278	:douta	=	16'h	cc69;
58279	:douta	=	16'h	cc69;
58280	:douta	=	16'h	cc69;
58281	:douta	=	16'h	cc69;
58282	:douta	=	16'h	cc69;
58283	:douta	=	16'h	cc69;
58284	:douta	=	16'h	cc69;
58285	:douta	=	16'h	cc69;
58286	:douta	=	16'h	cc69;
58287	:douta	=	16'h	cc69;
58288	:douta	=	16'h	cc69;
58289	:douta	=	16'h	cc69;
58290	:douta	=	16'h	cc69;
58291	:douta	=	16'h	cc69;
58292	:douta	=	16'h	cc69;
58293	:douta	=	16'h	cc69;
58294	:douta	=	16'h	cc69;
58295	:douta	=	16'h	cc69;
58296	:douta	=	16'h	cc49;
58297	:douta	=	16'h	cc69;
58298	:douta	=	16'h	cc69;
58299	:douta	=	16'h	cc69;
58300	:douta	=	16'h	cc49;
58301	:douta	=	16'h	cc69;
58302	:douta	=	16'h	cc69;
58303	:douta	=	16'h	cc69;
58304	:douta	=	16'h	c449;
58305	:douta	=	16'h	c449;
58306	:douta	=	16'h	cc69;
58307	:douta	=	16'h	cc49;
58308	:douta	=	16'h	cc49;
58309	:douta	=	16'h	c449;
58310	:douta	=	16'h	c449;
58311	:douta	=	16'h	c449;
58312	:douta	=	16'h	c428;
58313	:douta	=	16'h	c449;
58314	:douta	=	16'h	c429;
58315	:douta	=	16'h	c429;
58316	:douta	=	16'h	c429;
58317	:douta	=	16'h	c429;
58318	:douta	=	16'h	c429;
58319	:douta	=	16'h	c429;
58320	:douta	=	16'h	c429;
58321	:douta	=	16'h	bc08;
58322	:douta	=	16'h	c429;
58323	:douta	=	16'h	bc09;
58324	:douta	=	16'h	bc29;
58325	:douta	=	16'h	bc09;
58326	:douta	=	16'h	bc09;
58327	:douta	=	16'h	bc09;
58328	:douta	=	16'h	bc09;
58329	:douta	=	16'h	bc09;
58330	:douta	=	16'h	bbe9;
58331	:douta	=	16'h	bbe9;
58332	:douta	=	16'h	bbe9;
58333	:douta	=	16'h	bbe9;
58334	:douta	=	16'h	b3e8;
58335	:douta	=	16'h	bbe9;
58336	:douta	=	16'h	b3e8;
58337	:douta	=	16'h	bbe9;
58338	:douta	=	16'h	b3c8;
58339	:douta	=	16'h	b3e9;
58340	:douta	=	16'h	b3c8;
58341	:douta	=	16'h	b3c9;
58342	:douta	=	16'h	b3c9;
58343	:douta	=	16'h	b3c8;
58344	:douta	=	16'h	b3c9;
58345	:douta	=	16'h	b3c9;
58346	:douta	=	16'h	b3c9;
58347	:douta	=	16'h	b3c8;
58348	:douta	=	16'h	b3c8;
58349	:douta	=	16'h	b3c8;
58350	:douta	=	16'h	aba9;
58351	:douta	=	16'h	aba9;
58352	:douta	=	16'h	aba9;
58353	:douta	=	16'h	aba8;
58354	:douta	=	16'h	aba9;
58355	:douta	=	16'h	aba9;
58356	:douta	=	16'h	aba9;
58357	:douta	=	16'h	aba9;
58358	:douta	=	16'h	aba9;
58359	:douta	=	16'h	ab88;
58360	:douta	=	16'h	ab88;
58361	:douta	=	16'h	ab88;
58362	:douta	=	16'h	ab89;
58363	:douta	=	16'h	a389;
58364	:douta	=	16'h	a389;
58365	:douta	=	16'h	ab89;
58366	:douta	=	16'h	a389;
58367	:douta	=	16'h	a368;
58368	:douta	=	16'h	a4f5;
58369	:douta	=	16'h	a4b4;
58370	:douta	=	16'h	a4f5;
58371	:douta	=	16'h	8cb6;
58372	:douta	=	16'h	8c95;
58373	:douta	=	16'h	94f8;
58374	:douta	=	16'h	20c3;
58375	:douta	=	16'h	28c3;
58376	:douta	=	16'h	28e3;
58377	:douta	=	16'h	2904;
58378	:douta	=	16'h	28e3;
58379	:douta	=	16'h	28e3;
58380	:douta	=	16'h	28e3;
58381	:douta	=	16'h	20c2;
58382	:douta	=	16'h	28e3;
58383	:douta	=	16'h	28e3;
58384	:douta	=	16'h	20c3;
58385	:douta	=	16'h	28e3;
58386	:douta	=	16'h	20a3;
58387	:douta	=	16'h	20e3;
58388	:douta	=	16'h	20c2;
58389	:douta	=	16'h	20c2;
58390	:douta	=	16'h	20a2;
58391	:douta	=	16'h	20a2;
58392	:douta	=	16'h	20a2;
58393	:douta	=	16'h	20c2;
58394	:douta	=	16'h	28e3;
58395	:douta	=	16'h	28c3;
58396	:douta	=	16'h	28c2;
58397	:douta	=	16'h	28e3;
58398	:douta	=	16'h	28e3;
58399	:douta	=	16'h	28e3;
58400	:douta	=	16'h	3103;
58401	:douta	=	16'h	3103;
58402	:douta	=	16'h	3103;
58403	:douta	=	16'h	3103;
58404	:douta	=	16'h	3923;
58405	:douta	=	16'h	4124;
58406	:douta	=	16'h	4124;
58407	:douta	=	16'h	4163;
58408	:douta	=	16'h	4964;
58409	:douta	=	16'h	4963;
58410	:douta	=	16'h	4a08;
58411	:douta	=	16'h	2967;
58412	:douta	=	16'h	28e4;
58413	:douta	=	16'h	59a4;
58414	:douta	=	16'h	59c4;
58415	:douta	=	16'h	61c4;
58416	:douta	=	16'h	61c4;
58417	:douta	=	16'h	6204;
58418	:douta	=	16'h	6204;
58419	:douta	=	16'h	6a24;
58420	:douta	=	16'h	6a24;
58421	:douta	=	16'h	7244;
58422	:douta	=	16'h	7224;
58423	:douta	=	16'h	6aa8;
58424	:douta	=	16'h	accf;
58425	:douta	=	16'h	7224;
58426	:douta	=	16'h	7a85;
58427	:douta	=	16'h	7a85;
58428	:douta	=	16'h	7a85;
58429	:douta	=	16'h	82a5;
58430	:douta	=	16'h	82a6;
58431	:douta	=	16'h	82c6;
58432	:douta	=	16'h	8ac6;
58433	:douta	=	16'h	8ae7;
58434	:douta	=	16'h	82c6;
58435	:douta	=	16'h	8ac6;
58436	:douta	=	16'h	8ae6;
58437	:douta	=	16'h	8ae7;
58438	:douta	=	16'h	8ae6;
58439	:douta	=	16'h	9306;
58440	:douta	=	16'h	9b27;
58441	:douta	=	16'h	9b26;
58442	:douta	=	16'h	7285;
58443	:douta	=	16'h	51c5;
58444	:douta	=	16'h	a3c9;
58445	:douta	=	16'h	9baa;
58446	:douta	=	16'h	93aa;
58447	:douta	=	16'h	940c;
58448	:douta	=	16'h	a46d;
58449	:douta	=	16'h	c572;
58450	:douta	=	16'h	7329;
58451	:douta	=	16'h	bbe7;
58452	:douta	=	16'h	b3a7;
58453	:douta	=	16'h	b3c7;
58454	:douta	=	16'h	b3c6;
58455	:douta	=	16'h	b3e7;
58456	:douta	=	16'h	bbe7;
58457	:douta	=	16'h	bbe7;
58458	:douta	=	16'h	bbe7;
58459	:douta	=	16'h	bc07;
58460	:douta	=	16'h	bc08;
58461	:douta	=	16'h	c408;
58462	:douta	=	16'h	c428;
58463	:douta	=	16'h	c428;
58464	:douta	=	16'h	c428;
58465	:douta	=	16'h	c428;
58466	:douta	=	16'h	c428;
58467	:douta	=	16'h	c428;
58468	:douta	=	16'h	c428;
58469	:douta	=	16'h	c427;
58470	:douta	=	16'h	c448;
58471	:douta	=	16'h	c448;
58472	:douta	=	16'h	cc48;
58473	:douta	=	16'h	cc48;
58474	:douta	=	16'h	c448;
58475	:douta	=	16'h	cc48;
58476	:douta	=	16'h	cc48;
58477	:douta	=	16'h	cc48;
58478	:douta	=	16'h	cc68;
58479	:douta	=	16'h	cc69;
58480	:douta	=	16'h	cc69;
58481	:douta	=	16'h	cc68;
58482	:douta	=	16'h	cc68;
58483	:douta	=	16'h	cc68;
58484	:douta	=	16'h	cc68;
58485	:douta	=	16'h	cc68;
58486	:douta	=	16'h	cc68;
58487	:douta	=	16'h	cc68;
58488	:douta	=	16'h	cc69;
58489	:douta	=	16'h	cc68;
58490	:douta	=	16'h	cc68;
58491	:douta	=	16'h	cc68;
58492	:douta	=	16'h	cc68;
58493	:douta	=	16'h	cc88;
58494	:douta	=	16'h	cc88;
58495	:douta	=	16'h	cc68;
58496	:douta	=	16'h	cc88;
58497	:douta	=	16'h	cc68;
58498	:douta	=	16'h	cc89;
58499	:douta	=	16'h	cc89;
58500	:douta	=	16'h	cc89;
58501	:douta	=	16'h	cc89;
58502	:douta	=	16'h	cc89;
58503	:douta	=	16'h	cc69;
58504	:douta	=	16'h	cc8a;
58505	:douta	=	16'h	cc69;
58506	:douta	=	16'h	cc89;
58507	:douta	=	16'h	cc69;
58508	:douta	=	16'h	cc69;
58509	:douta	=	16'h	cc69;
58510	:douta	=	16'h	cc69;
58511	:douta	=	16'h	cc69;
58512	:douta	=	16'h	cc89;
58513	:douta	=	16'h	cc89;
58514	:douta	=	16'h	cc69;
58515	:douta	=	16'h	cc89;
58516	:douta	=	16'h	cc89;
58517	:douta	=	16'h	d489;
58518	:douta	=	16'h	cc8a;
58519	:douta	=	16'h	cc89;
58520	:douta	=	16'h	cc89;
58521	:douta	=	16'h	cc89;
58522	:douta	=	16'h	d489;
58523	:douta	=	16'h	d489;
58524	:douta	=	16'h	cc69;
58525	:douta	=	16'h	cc89;
58526	:douta	=	16'h	cc89;
58527	:douta	=	16'h	cc89;
58528	:douta	=	16'h	cc89;
58529	:douta	=	16'h	cc69;
58530	:douta	=	16'h	d468;
58531	:douta	=	16'h	ad73;
58532	:douta	=	16'h	e696;
58533	:douta	=	16'h	cc47;
58534	:douta	=	16'h	cc69;
58535	:douta	=	16'h	cc68;
58536	:douta	=	16'h	cc69;
58537	:douta	=	16'h	cc69;
58538	:douta	=	16'h	cc69;
58539	:douta	=	16'h	cc69;
58540	:douta	=	16'h	cc69;
58541	:douta	=	16'h	cc69;
58542	:douta	=	16'h	cc69;
58543	:douta	=	16'h	cc69;
58544	:douta	=	16'h	cc69;
58545	:douta	=	16'h	cc69;
58546	:douta	=	16'h	cc69;
58547	:douta	=	16'h	cc69;
58548	:douta	=	16'h	cc69;
58549	:douta	=	16'h	cc69;
58550	:douta	=	16'h	cc69;
58551	:douta	=	16'h	cc69;
58552	:douta	=	16'h	cc69;
58553	:douta	=	16'h	c449;
58554	:douta	=	16'h	cc69;
58555	:douta	=	16'h	cc69;
58556	:douta	=	16'h	cc69;
58557	:douta	=	16'h	cc49;
58558	:douta	=	16'h	c449;
58559	:douta	=	16'h	cc69;
58560	:douta	=	16'h	c449;
58561	:douta	=	16'h	c449;
58562	:douta	=	16'h	cc49;
58563	:douta	=	16'h	cc49;
58564	:douta	=	16'h	cc49;
58565	:douta	=	16'h	cc49;
58566	:douta	=	16'h	c449;
58567	:douta	=	16'h	c449;
58568	:douta	=	16'h	c449;
58569	:douta	=	16'h	c428;
58570	:douta	=	16'h	c429;
58571	:douta	=	16'h	c429;
58572	:douta	=	16'h	c429;
58573	:douta	=	16'h	c429;
58574	:douta	=	16'h	c429;
58575	:douta	=	16'h	c429;
58576	:douta	=	16'h	c429;
58577	:douta	=	16'h	c409;
58578	:douta	=	16'h	bc29;
58579	:douta	=	16'h	bc09;
58580	:douta	=	16'h	bc29;
58581	:douta	=	16'h	bc09;
58582	:douta	=	16'h	bc09;
58583	:douta	=	16'h	bc09;
58584	:douta	=	16'h	bbe9;
58585	:douta	=	16'h	bc09;
58586	:douta	=	16'h	bbe9;
58587	:douta	=	16'h	bbe9;
58588	:douta	=	16'h	bc09;
58589	:douta	=	16'h	bbe9;
58590	:douta	=	16'h	bc09;
58591	:douta	=	16'h	b3e8;
58592	:douta	=	16'h	bbe9;
58593	:douta	=	16'h	b3c9;
58594	:douta	=	16'h	b3e9;
58595	:douta	=	16'h	b3e9;
58596	:douta	=	16'h	b3c8;
58597	:douta	=	16'h	b3c9;
58598	:douta	=	16'h	b3c9;
58599	:douta	=	16'h	b3c9;
58600	:douta	=	16'h	b3c9;
58601	:douta	=	16'h	b3c9;
58602	:douta	=	16'h	b3c9;
58603	:douta	=	16'h	b3c9;
58604	:douta	=	16'h	b3c8;
58605	:douta	=	16'h	b3c9;
58606	:douta	=	16'h	abc9;
58607	:douta	=	16'h	aba9;
58608	:douta	=	16'h	b3c8;
58609	:douta	=	16'h	b3c8;
58610	:douta	=	16'h	aba9;
58611	:douta	=	16'h	aba9;
58612	:douta	=	16'h	ab89;
58613	:douta	=	16'h	aba9;
58614	:douta	=	16'h	aba9;
58615	:douta	=	16'h	ab89;
58616	:douta	=	16'h	aba9;
58617	:douta	=	16'h	aba9;
58618	:douta	=	16'h	a389;
58619	:douta	=	16'h	ab89;
58620	:douta	=	16'h	a389;
58621	:douta	=	16'h	a389;
58622	:douta	=	16'h	ab89;
58623	:douta	=	16'h	a368;
58624	:douta	=	16'h	b535;
58625	:douta	=	16'h	94b4;
58626	:douta	=	16'h	9cd5;
58627	:douta	=	16'h	94d6;
58628	:douta	=	16'h	8495;
58629	:douta	=	16'h	8475;
58630	:douta	=	16'h	2081;
58631	:douta	=	16'h	2904;
58632	:douta	=	16'h	2903;
58633	:douta	=	16'h	2904;
58634	:douta	=	16'h	2904;
58635	:douta	=	16'h	28e3;
58636	:douta	=	16'h	28e3;
58637	:douta	=	16'h	28e3;
58638	:douta	=	16'h	28e3;
58639	:douta	=	16'h	28e3;
58640	:douta	=	16'h	20e3;
58641	:douta	=	16'h	20e3;
58642	:douta	=	16'h	20e3;
58643	:douta	=	16'h	20e3;
58644	:douta	=	16'h	20e3;
58645	:douta	=	16'h	20a2;
58646	:douta	=	16'h	20a2;
58647	:douta	=	16'h	20a2;
58648	:douta	=	16'h	20c2;
58649	:douta	=	16'h	20c2;
58650	:douta	=	16'h	28c3;
58651	:douta	=	16'h	20c2;
58652	:douta	=	16'h	28e3;
58653	:douta	=	16'h	28e3;
58654	:douta	=	16'h	28e3;
58655	:douta	=	16'h	28e2;
58656	:douta	=	16'h	3103;
58657	:douta	=	16'h	30e2;
58658	:douta	=	16'h	3123;
58659	:douta	=	16'h	3103;
58660	:douta	=	16'h	3944;
58661	:douta	=	16'h	4124;
58662	:douta	=	16'h	4143;
58663	:douta	=	16'h	4163;
58664	:douta	=	16'h	4163;
58665	:douta	=	16'h	4984;
58666	:douta	=	16'h	526a;
58667	:douta	=	16'h	1905;
58668	:douta	=	16'h	3924;
58669	:douta	=	16'h	61c3;
58670	:douta	=	16'h	59c4;
58671	:douta	=	16'h	59c4;
58672	:douta	=	16'h	61e4;
58673	:douta	=	16'h	6204;
58674	:douta	=	16'h	6204;
58675	:douta	=	16'h	6a04;
58676	:douta	=	16'h	6a24;
58677	:douta	=	16'h	7224;
58678	:douta	=	16'h	7224;
58679	:douta	=	16'h	7b6c;
58680	:douta	=	16'h	8baa;
58681	:douta	=	16'h	7223;
58682	:douta	=	16'h	7a85;
58683	:douta	=	16'h	7a85;
58684	:douta	=	16'h	7a85;
58685	:douta	=	16'h	82a5;
58686	:douta	=	16'h	82a5;
58687	:douta	=	16'h	82a6;
58688	:douta	=	16'h	8ac6;
58689	:douta	=	16'h	8ac6;
58690	:douta	=	16'h	8ac6;
58691	:douta	=	16'h	8ae7;
58692	:douta	=	16'h	8ac6;
58693	:douta	=	16'h	8ac6;
58694	:douta	=	16'h	9307;
58695	:douta	=	16'h	9306;
58696	:douta	=	16'h	9326;
58697	:douta	=	16'h	9326;
58698	:douta	=	16'h	ab87;
58699	:douta	=	16'h	6a24;
58700	:douta	=	16'h	e676;
58701	:douta	=	16'h	de97;
58702	:douta	=	16'h	cdf4;
58703	:douta	=	16'h	d635;
58704	:douta	=	16'h	d635;
58705	:douta	=	16'h	de97;
58706	:douta	=	16'h	6ae7;
58707	:douta	=	16'h	b3e7;
58708	:douta	=	16'h	b3c7;
58709	:douta	=	16'h	b3c7;
58710	:douta	=	16'h	b3e7;
58711	:douta	=	16'h	b3e7;
58712	:douta	=	16'h	bbe8;
58713	:douta	=	16'h	bbe7;
58714	:douta	=	16'h	bc07;
58715	:douta	=	16'h	bc07;
58716	:douta	=	16'h	bc07;
58717	:douta	=	16'h	bc07;
58718	:douta	=	16'h	bc07;
58719	:douta	=	16'h	bc07;
58720	:douta	=	16'h	c407;
58721	:douta	=	16'h	c428;
58722	:douta	=	16'h	c428;
58723	:douta	=	16'h	c428;
58724	:douta	=	16'h	c428;
58725	:douta	=	16'h	c448;
58726	:douta	=	16'h	c448;
58727	:douta	=	16'h	c448;
58728	:douta	=	16'h	c428;
58729	:douta	=	16'h	c448;
58730	:douta	=	16'h	c448;
58731	:douta	=	16'h	c448;
58732	:douta	=	16'h	cc49;
58733	:douta	=	16'h	cc49;
58734	:douta	=	16'h	c448;
58735	:douta	=	16'h	c448;
58736	:douta	=	16'h	c448;
58737	:douta	=	16'h	cc68;
58738	:douta	=	16'h	cc68;
58739	:douta	=	16'h	cc68;
58740	:douta	=	16'h	cc68;
58741	:douta	=	16'h	cc68;
58742	:douta	=	16'h	cc68;
58743	:douta	=	16'h	cc68;
58744	:douta	=	16'h	cc68;
58745	:douta	=	16'h	cc68;
58746	:douta	=	16'h	cc68;
58747	:douta	=	16'h	cc68;
58748	:douta	=	16'h	cc68;
58749	:douta	=	16'h	cc68;
58750	:douta	=	16'h	cc68;
58751	:douta	=	16'h	cc89;
58752	:douta	=	16'h	cc69;
58753	:douta	=	16'h	cc89;
58754	:douta	=	16'h	cc68;
58755	:douta	=	16'h	cc69;
58756	:douta	=	16'h	cc69;
58757	:douta	=	16'h	cc69;
58758	:douta	=	16'h	cc69;
58759	:douta	=	16'h	cc89;
58760	:douta	=	16'h	cc89;
58761	:douta	=	16'h	cc89;
58762	:douta	=	16'h	cc89;
58763	:douta	=	16'h	cc89;
58764	:douta	=	16'h	cc69;
58765	:douta	=	16'h	cc89;
58766	:douta	=	16'h	cc69;
58767	:douta	=	16'h	cc89;
58768	:douta	=	16'h	cc69;
58769	:douta	=	16'h	cc89;
58770	:douta	=	16'h	cc89;
58771	:douta	=	16'h	cc8a;
58772	:douta	=	16'h	cc89;
58773	:douta	=	16'h	cc89;
58774	:douta	=	16'h	cc89;
58775	:douta	=	16'h	d48a;
58776	:douta	=	16'h	cc8a;
58777	:douta	=	16'h	cc8a;
58778	:douta	=	16'h	cc89;
58779	:douta	=	16'h	cc89;
58780	:douta	=	16'h	cc89;
58781	:douta	=	16'h	cc89;
58782	:douta	=	16'h	cc89;
58783	:douta	=	16'h	cc89;
58784	:douta	=	16'h	cc89;
58785	:douta	=	16'h	cc89;
58786	:douta	=	16'h	d468;
58787	:douta	=	16'h	ad73;
58788	:douta	=	16'h	e696;
58789	:douta	=	16'h	cc47;
58790	:douta	=	16'h	cc89;
58791	:douta	=	16'h	cc69;
58792	:douta	=	16'h	cc69;
58793	:douta	=	16'h	cc89;
58794	:douta	=	16'h	cc69;
58795	:douta	=	16'h	cc69;
58796	:douta	=	16'h	cc89;
58797	:douta	=	16'h	cc69;
58798	:douta	=	16'h	cc69;
58799	:douta	=	16'h	cc69;
58800	:douta	=	16'h	cc69;
58801	:douta	=	16'h	cc69;
58802	:douta	=	16'h	cc69;
58803	:douta	=	16'h	cc69;
58804	:douta	=	16'h	cc69;
58805	:douta	=	16'h	cc69;
58806	:douta	=	16'h	cc69;
58807	:douta	=	16'h	cc69;
58808	:douta	=	16'h	cc49;
58809	:douta	=	16'h	cc69;
58810	:douta	=	16'h	cc69;
58811	:douta	=	16'h	cc69;
58812	:douta	=	16'h	cc49;
58813	:douta	=	16'h	cc69;
58814	:douta	=	16'h	c468;
58815	:douta	=	16'h	c448;
58816	:douta	=	16'h	c449;
58817	:douta	=	16'h	cc69;
58818	:douta	=	16'h	cc49;
58819	:douta	=	16'h	c449;
58820	:douta	=	16'h	c449;
58821	:douta	=	16'h	c449;
58822	:douta	=	16'h	c449;
58823	:douta	=	16'h	c449;
58824	:douta	=	16'h	c429;
58825	:douta	=	16'h	c429;
58826	:douta	=	16'h	c429;
58827	:douta	=	16'h	c429;
58828	:douta	=	16'h	c449;
58829	:douta	=	16'h	bc09;
58830	:douta	=	16'h	c429;
58831	:douta	=	16'h	c429;
58832	:douta	=	16'h	c429;
58833	:douta	=	16'h	c429;
58834	:douta	=	16'h	bc29;
58835	:douta	=	16'h	bc29;
58836	:douta	=	16'h	bc09;
58837	:douta	=	16'h	bc29;
58838	:douta	=	16'h	bc09;
58839	:douta	=	16'h	bc09;
58840	:douta	=	16'h	bc09;
58841	:douta	=	16'h	bc09;
58842	:douta	=	16'h	bbe9;
58843	:douta	=	16'h	bc09;
58844	:douta	=	16'h	bbe9;
58845	:douta	=	16'h	bbe9;
58846	:douta	=	16'h	bc09;
58847	:douta	=	16'h	bbe9;
58848	:douta	=	16'h	b3e9;
58849	:douta	=	16'h	bbe9;
58850	:douta	=	16'h	b3e9;
58851	:douta	=	16'h	b3e9;
58852	:douta	=	16'h	b3c8;
58853	:douta	=	16'h	b3c8;
58854	:douta	=	16'h	b3c9;
58855	:douta	=	16'h	b3e9;
58856	:douta	=	16'h	b3c9;
58857	:douta	=	16'h	b3c9;
58858	:douta	=	16'h	b3c9;
58859	:douta	=	16'h	b3c9;
58860	:douta	=	16'h	b3c9;
58861	:douta	=	16'h	b3c9;
58862	:douta	=	16'h	aba9;
58863	:douta	=	16'h	abc9;
58864	:douta	=	16'h	aba9;
58865	:douta	=	16'h	aba9;
58866	:douta	=	16'h	b3c8;
58867	:douta	=	16'h	aba8;
58868	:douta	=	16'h	aba9;
58869	:douta	=	16'h	aba9;
58870	:douta	=	16'h	aba9;
58871	:douta	=	16'h	aba9;
58872	:douta	=	16'h	ab89;
58873	:douta	=	16'h	ab89;
58874	:douta	=	16'h	a389;
58875	:douta	=	16'h	ab89;
58876	:douta	=	16'h	a389;
58877	:douta	=	16'h	a388;
58878	:douta	=	16'h	a388;
58879	:douta	=	16'h	a368;
58880	:douta	=	16'h	b556;
58881	:douta	=	16'h	9cb5;
58882	:douta	=	16'h	94b5;
58883	:douta	=	16'h	94f6;
58884	:douta	=	16'h	94f7;
58885	:douta	=	16'h	6b90;
58886	:douta	=	16'h	2904;
58887	:douta	=	16'h	2904;
58888	:douta	=	16'h	20e3;
58889	:douta	=	16'h	2904;
58890	:douta	=	16'h	2904;
58891	:douta	=	16'h	28e3;
58892	:douta	=	16'h	2903;
58893	:douta	=	16'h	28e3;
58894	:douta	=	16'h	28e3;
58895	:douta	=	16'h	28e3;
58896	:douta	=	16'h	20e3;
58897	:douta	=	16'h	20e3;
58898	:douta	=	16'h	20e3;
58899	:douta	=	16'h	20c3;
58900	:douta	=	16'h	20e3;
58901	:douta	=	16'h	18a2;
58902	:douta	=	16'h	20a2;
58903	:douta	=	16'h	20a2;
58904	:douta	=	16'h	20a2;
58905	:douta	=	16'h	20c2;
58906	:douta	=	16'h	20a2;
58907	:douta	=	16'h	20a2;
58908	:douta	=	16'h	28e3;
58909	:douta	=	16'h	28e3;
58910	:douta	=	16'h	28e3;
58911	:douta	=	16'h	28e3;
58912	:douta	=	16'h	3103;
58913	:douta	=	16'h	3103;
58914	:douta	=	16'h	3123;
58915	:douta	=	16'h	3923;
58916	:douta	=	16'h	3943;
58917	:douta	=	16'h	4124;
58918	:douta	=	16'h	4143;
58919	:douta	=	16'h	4964;
58920	:douta	=	16'h	4964;
58921	:douta	=	16'h	49a5;
58922	:douta	=	16'h	528b;
58923	:douta	=	16'h	10e5;
58924	:douta	=	16'h	4985;
58925	:douta	=	16'h	61e4;
58926	:douta	=	16'h	59c4;
58927	:douta	=	16'h	59c4;
58928	:douta	=	16'h	61e4;
58929	:douta	=	16'h	6204;
58930	:douta	=	16'h	6a24;
58931	:douta	=	16'h	6a04;
58932	:douta	=	16'h	6a24;
58933	:douta	=	16'h	7224;
58934	:douta	=	16'h	7265;
58935	:douta	=	16'h	83ee;
58936	:douta	=	16'h	8327;
58937	:douta	=	16'h	7224;
58938	:douta	=	16'h	8286;
58939	:douta	=	16'h	8285;
58940	:douta	=	16'h	8285;
58941	:douta	=	16'h	82a5;
58942	:douta	=	16'h	82c6;
58943	:douta	=	16'h	82c6;
58944	:douta	=	16'h	82c6;
58945	:douta	=	16'h	8ac6;
58946	:douta	=	16'h	8ac6;
58947	:douta	=	16'h	8b07;
58948	:douta	=	16'h	8ac6;
58949	:douta	=	16'h	8ac6;
58950	:douta	=	16'h	9307;
58951	:douta	=	16'h	9306;
58952	:douta	=	16'h	9326;
58953	:douta	=	16'h	9b27;
58954	:douta	=	16'h	9b27;
58955	:douta	=	16'h	a347;
58956	:douta	=	16'h	93ee;
58957	:douta	=	16'h	f6d8;
58958	:douta	=	16'h	de76;
58959	:douta	=	16'h	c551;
58960	:douta	=	16'h	e696;
58961	:douta	=	16'h	d656;
58962	:douta	=	16'h	6267;
58963	:douta	=	16'h	b3e7;
58964	:douta	=	16'h	aba7;
58965	:douta	=	16'h	b3c7;
58966	:douta	=	16'h	b3e7;
58967	:douta	=	16'h	b3e7;
58968	:douta	=	16'h	b3e7;
58969	:douta	=	16'h	bbe8;
58970	:douta	=	16'h	bbe7;
58971	:douta	=	16'h	bc07;
58972	:douta	=	16'h	bc07;
58973	:douta	=	16'h	bc07;
58974	:douta	=	16'h	bc07;
58975	:douta	=	16'h	c407;
58976	:douta	=	16'h	c407;
58977	:douta	=	16'h	c428;
58978	:douta	=	16'h	c428;
58979	:douta	=	16'h	c428;
58980	:douta	=	16'h	c428;
58981	:douta	=	16'h	c428;
58982	:douta	=	16'h	c448;
58983	:douta	=	16'h	c448;
58984	:douta	=	16'h	c448;
58985	:douta	=	16'h	c448;
58986	:douta	=	16'h	cc48;
58987	:douta	=	16'h	cc48;
58988	:douta	=	16'h	cc48;
58989	:douta	=	16'h	c449;
58990	:douta	=	16'h	cc68;
58991	:douta	=	16'h	cc68;
58992	:douta	=	16'h	cc68;
58993	:douta	=	16'h	cc67;
58994	:douta	=	16'h	cc67;
58995	:douta	=	16'h	cc68;
58996	:douta	=	16'h	cc68;
58997	:douta	=	16'h	cc68;
58998	:douta	=	16'h	cc68;
58999	:douta	=	16'h	cc68;
59000	:douta	=	16'h	cc68;
59001	:douta	=	16'h	cc68;
59002	:douta	=	16'h	cc68;
59003	:douta	=	16'h	cc88;
59004	:douta	=	16'h	cc68;
59005	:douta	=	16'h	cc69;
59006	:douta	=	16'h	cc68;
59007	:douta	=	16'h	cc69;
59008	:douta	=	16'h	cc69;
59009	:douta	=	16'h	cc69;
59010	:douta	=	16'h	cc68;
59011	:douta	=	16'h	cc69;
59012	:douta	=	16'h	cc89;
59013	:douta	=	16'h	cc69;
59014	:douta	=	16'h	d489;
59015	:douta	=	16'h	cc69;
59016	:douta	=	16'h	cc89;
59017	:douta	=	16'h	cc89;
59018	:douta	=	16'h	cc89;
59019	:douta	=	16'h	cc69;
59020	:douta	=	16'h	cc89;
59021	:douta	=	16'h	cc69;
59022	:douta	=	16'h	cc89;
59023	:douta	=	16'h	cc8a;
59024	:douta	=	16'h	cc69;
59025	:douta	=	16'h	cc89;
59026	:douta	=	16'h	cc89;
59027	:douta	=	16'h	cc8a;
59028	:douta	=	16'h	cc89;
59029	:douta	=	16'h	d489;
59030	:douta	=	16'h	cc89;
59031	:douta	=	16'h	cc8a;
59032	:douta	=	16'h	cc89;
59033	:douta	=	16'h	cc89;
59034	:douta	=	16'h	cc89;
59035	:douta	=	16'h	cc89;
59036	:douta	=	16'h	cc89;
59037	:douta	=	16'h	cc89;
59038	:douta	=	16'h	cc89;
59039	:douta	=	16'h	cc89;
59040	:douta	=	16'h	cc89;
59041	:douta	=	16'h	cc89;
59042	:douta	=	16'h	d488;
59043	:douta	=	16'h	ad74;
59044	:douta	=	16'h	e696;
59045	:douta	=	16'h	cc47;
59046	:douta	=	16'h	cc89;
59047	:douta	=	16'h	cc89;
59048	:douta	=	16'h	cc69;
59049	:douta	=	16'h	cc89;
59050	:douta	=	16'h	cc69;
59051	:douta	=	16'h	cc69;
59052	:douta	=	16'h	cc69;
59053	:douta	=	16'h	cc69;
59054	:douta	=	16'h	cc69;
59055	:douta	=	16'h	cc69;
59056	:douta	=	16'h	cc69;
59057	:douta	=	16'h	cc69;
59058	:douta	=	16'h	cc69;
59059	:douta	=	16'h	cc69;
59060	:douta	=	16'h	cc69;
59061	:douta	=	16'h	cc69;
59062	:douta	=	16'h	cc69;
59063	:douta	=	16'h	cc69;
59064	:douta	=	16'h	cc69;
59065	:douta	=	16'h	cc69;
59066	:douta	=	16'h	cc69;
59067	:douta	=	16'h	cc49;
59068	:douta	=	16'h	cc69;
59069	:douta	=	16'h	c468;
59070	:douta	=	16'h	c468;
59071	:douta	=	16'h	cc69;
59072	:douta	=	16'h	cc49;
59073	:douta	=	16'h	cc49;
59074	:douta	=	16'h	c449;
59075	:douta	=	16'h	c449;
59076	:douta	=	16'h	c449;
59077	:douta	=	16'h	c448;
59078	:douta	=	16'h	c449;
59079	:douta	=	16'h	c449;
59080	:douta	=	16'h	c429;
59081	:douta	=	16'h	c429;
59082	:douta	=	16'h	c429;
59083	:douta	=	16'h	c429;
59084	:douta	=	16'h	c429;
59085	:douta	=	16'h	c429;
59086	:douta	=	16'h	c429;
59087	:douta	=	16'h	bc29;
59088	:douta	=	16'h	c429;
59089	:douta	=	16'h	bc29;
59090	:douta	=	16'h	c429;
59091	:douta	=	16'h	c429;
59092	:douta	=	16'h	bc09;
59093	:douta	=	16'h	bc29;
59094	:douta	=	16'h	c429;
59095	:douta	=	16'h	bc09;
59096	:douta	=	16'h	bc29;
59097	:douta	=	16'h	bc09;
59098	:douta	=	16'h	bc09;
59099	:douta	=	16'h	bbe9;
59100	:douta	=	16'h	bc09;
59101	:douta	=	16'h	bc09;
59102	:douta	=	16'h	bbe9;
59103	:douta	=	16'h	bc09;
59104	:douta	=	16'h	bbe9;
59105	:douta	=	16'h	b3e9;
59106	:douta	=	16'h	b3e9;
59107	:douta	=	16'h	b3e9;
59108	:douta	=	16'h	b3c8;
59109	:douta	=	16'h	b3e9;
59110	:douta	=	16'h	b3c9;
59111	:douta	=	16'h	b3c9;
59112	:douta	=	16'h	b3c9;
59113	:douta	=	16'h	b3c9;
59114	:douta	=	16'h	b3c9;
59115	:douta	=	16'h	b3c9;
59116	:douta	=	16'h	b3c9;
59117	:douta	=	16'h	b3c8;
59118	:douta	=	16'h	aba9;
59119	:douta	=	16'h	b3c9;
59120	:douta	=	16'h	aba9;
59121	:douta	=	16'h	abc9;
59122	:douta	=	16'h	aba9;
59123	:douta	=	16'h	aba9;
59124	:douta	=	16'h	aba9;
59125	:douta	=	16'h	aba9;
59126	:douta	=	16'h	aba9;
59127	:douta	=	16'h	aba9;
59128	:douta	=	16'h	aba8;
59129	:douta	=	16'h	a389;
59130	:douta	=	16'h	ab89;
59131	:douta	=	16'h	ab89;
59132	:douta	=	16'h	ab89;
59133	:douta	=	16'h	a389;
59134	:douta	=	16'h	a388;
59135	:douta	=	16'h	a388;
59136	:douta	=	16'h	a515;
59137	:douta	=	16'h	8c95;
59138	:douta	=	16'h	94d6;
59139	:douta	=	16'h	94f7;
59140	:douta	=	16'h	8454;
59141	:douta	=	16'h	2924;
59142	:douta	=	16'h	2924;
59143	:douta	=	16'h	28e3;
59144	:douta	=	16'h	28e3;
59145	:douta	=	16'h	3124;
59146	:douta	=	16'h	28e3;
59147	:douta	=	16'h	28e3;
59148	:douta	=	16'h	28e3;
59149	:douta	=	16'h	28e3;
59150	:douta	=	16'h	28e3;
59151	:douta	=	16'h	28e3;
59152	:douta	=	16'h	20c3;
59153	:douta	=	16'h	20c3;
59154	:douta	=	16'h	20e3;
59155	:douta	=	16'h	20e3;
59156	:douta	=	16'h	2904;
59157	:douta	=	16'h	20a2;
59158	:douta	=	16'h	20a2;
59159	:douta	=	16'h	20c2;
59160	:douta	=	16'h	20c2;
59161	:douta	=	16'h	20c2;
59162	:douta	=	16'h	28c3;
59163	:douta	=	16'h	28e3;
59164	:douta	=	16'h	28e2;
59165	:douta	=	16'h	28e3;
59166	:douta	=	16'h	2903;
59167	:douta	=	16'h	28e3;
59168	:douta	=	16'h	3103;
59169	:douta	=	16'h	3103;
59170	:douta	=	16'h	3123;
59171	:douta	=	16'h	3123;
59172	:douta	=	16'h	4144;
59173	:douta	=	16'h	4124;
59174	:douta	=	16'h	4143;
59175	:douta	=	16'h	4963;
59176	:douta	=	16'h	4964;
59177	:douta	=	16'h	49c7;
59178	:douta	=	16'h	528a;
59179	:douta	=	16'h	0884;
59180	:douta	=	16'h	59c4;
59181	:douta	=	16'h	59c4;
59182	:douta	=	16'h	59c4;
59183	:douta	=	16'h	59c4;
59184	:douta	=	16'h	61e4;
59185	:douta	=	16'h	6204;
59186	:douta	=	16'h	61e4;
59187	:douta	=	16'h	6a24;
59188	:douta	=	16'h	6a04;
59189	:douta	=	16'h	7224;
59190	:douta	=	16'h	7266;
59191	:douta	=	16'h	9cd1;
59192	:douta	=	16'h	7244;
59193	:douta	=	16'h	7a64;
59194	:douta	=	16'h	7a85;
59195	:douta	=	16'h	7a85;
59196	:douta	=	16'h	7a85;
59197	:douta	=	16'h	82a5;
59198	:douta	=	16'h	82a5;
59199	:douta	=	16'h	82c6;
59200	:douta	=	16'h	8ae6;
59201	:douta	=	16'h	8ac6;
59202	:douta	=	16'h	8ac6;
59203	:douta	=	16'h	8ae6;
59204	:douta	=	16'h	8ae7;
59205	:douta	=	16'h	9307;
59206	:douta	=	16'h	9307;
59207	:douta	=	16'h	9306;
59208	:douta	=	16'h	9b27;
59209	:douta	=	16'h	9b27;
59210	:douta	=	16'h	9b28;
59211	:douta	=	16'h	8aa5;
59212	:douta	=	16'h	d6b7;
59213	:douta	=	16'h	2985;
59214	:douta	=	16'h	0000;
59215	:douta	=	16'h	0000;
59216	:douta	=	16'h	934a;
59217	:douta	=	16'h	ad52;
59218	:douta	=	16'h	59c4;
59219	:douta	=	16'h	b3c7;
59220	:douta	=	16'h	b3c7;
59221	:douta	=	16'h	aba7;
59222	:douta	=	16'h	b3e7;
59223	:douta	=	16'h	b3e7;
59224	:douta	=	16'h	b3e8;
59225	:douta	=	16'h	bbe7;
59226	:douta	=	16'h	bbe7;
59227	:douta	=	16'h	bc07;
59228	:douta	=	16'h	bc08;
59229	:douta	=	16'h	bc07;
59230	:douta	=	16'h	c407;
59231	:douta	=	16'h	c428;
59232	:douta	=	16'h	c428;
59233	:douta	=	16'h	c428;
59234	:douta	=	16'h	c428;
59235	:douta	=	16'h	c428;
59236	:douta	=	16'h	c428;
59237	:douta	=	16'h	c448;
59238	:douta	=	16'h	c448;
59239	:douta	=	16'h	c448;
59240	:douta	=	16'h	c448;
59241	:douta	=	16'h	cc68;
59242	:douta	=	16'h	cc49;
59243	:douta	=	16'h	cc49;
59244	:douta	=	16'h	cc49;
59245	:douta	=	16'h	cc49;
59246	:douta	=	16'h	c448;
59247	:douta	=	16'h	cc68;
59248	:douta	=	16'h	cc68;
59249	:douta	=	16'h	cc68;
59250	:douta	=	16'h	cc68;
59251	:douta	=	16'h	cc68;
59252	:douta	=	16'h	cc68;
59253	:douta	=	16'h	cc68;
59254	:douta	=	16'h	cc68;
59255	:douta	=	16'h	cc68;
59256	:douta	=	16'h	cc68;
59257	:douta	=	16'h	cc68;
59258	:douta	=	16'h	cc68;
59259	:douta	=	16'h	cc68;
59260	:douta	=	16'h	cc68;
59261	:douta	=	16'h	cc69;
59262	:douta	=	16'h	cc69;
59263	:douta	=	16'h	cc69;
59264	:douta	=	16'h	cc89;
59265	:douta	=	16'h	cc68;
59266	:douta	=	16'h	cc89;
59267	:douta	=	16'h	cc89;
59268	:douta	=	16'h	cc89;
59269	:douta	=	16'h	cc89;
59270	:douta	=	16'h	cc69;
59271	:douta	=	16'h	cc8a;
59272	:douta	=	16'h	cc69;
59273	:douta	=	16'h	cc89;
59274	:douta	=	16'h	cc69;
59275	:douta	=	16'h	cc89;
59276	:douta	=	16'h	cc89;
59277	:douta	=	16'h	cc89;
59278	:douta	=	16'h	cc69;
59279	:douta	=	16'h	cc89;
59280	:douta	=	16'h	cc89;
59281	:douta	=	16'h	cc89;
59282	:douta	=	16'h	cc89;
59283	:douta	=	16'h	cc8a;
59284	:douta	=	16'h	cc69;
59285	:douta	=	16'h	cc69;
59286	:douta	=	16'h	cc8a;
59287	:douta	=	16'h	cc89;
59288	:douta	=	16'h	cc89;
59289	:douta	=	16'h	cc89;
59290	:douta	=	16'h	cc69;
59291	:douta	=	16'h	cc89;
59292	:douta	=	16'h	cc69;
59293	:douta	=	16'h	cc89;
59294	:douta	=	16'h	cc89;
59295	:douta	=	16'h	cc89;
59296	:douta	=	16'h	cc89;
59297	:douta	=	16'h	cc89;
59298	:douta	=	16'h	d488;
59299	:douta	=	16'h	b594;
59300	:douta	=	16'h	e696;
59301	:douta	=	16'h	cc47;
59302	:douta	=	16'h	cc69;
59303	:douta	=	16'h	cc69;
59304	:douta	=	16'h	cc89;
59305	:douta	=	16'h	cc69;
59306	:douta	=	16'h	cc69;
59307	:douta	=	16'h	cc69;
59308	:douta	=	16'h	cc69;
59309	:douta	=	16'h	cc69;
59310	:douta	=	16'h	cc69;
59311	:douta	=	16'h	cc89;
59312	:douta	=	16'h	cc69;
59313	:douta	=	16'h	cc89;
59314	:douta	=	16'h	cc69;
59315	:douta	=	16'h	cc69;
59316	:douta	=	16'h	cc69;
59317	:douta	=	16'h	cc69;
59318	:douta	=	16'h	cc69;
59319	:douta	=	16'h	cc69;
59320	:douta	=	16'h	cc49;
59321	:douta	=	16'h	cc49;
59322	:douta	=	16'h	cc49;
59323	:douta	=	16'h	cc69;
59324	:douta	=	16'h	cc49;
59325	:douta	=	16'h	cc69;
59326	:douta	=	16'h	cc69;
59327	:douta	=	16'h	cc49;
59328	:douta	=	16'h	c449;
59329	:douta	=	16'h	c449;
59330	:douta	=	16'h	c449;
59331	:douta	=	16'h	c449;
59332	:douta	=	16'h	c449;
59333	:douta	=	16'h	c449;
59334	:douta	=	16'h	c429;
59335	:douta	=	16'h	c429;
59336	:douta	=	16'h	c429;
59337	:douta	=	16'h	c429;
59338	:douta	=	16'h	c449;
59339	:douta	=	16'h	c449;
59340	:douta	=	16'h	c449;
59341	:douta	=	16'h	c449;
59342	:douta	=	16'h	bc29;
59343	:douta	=	16'h	c429;
59344	:douta	=	16'h	bc09;
59345	:douta	=	16'h	c429;
59346	:douta	=	16'h	bc29;
59347	:douta	=	16'h	bc29;
59348	:douta	=	16'h	bc09;
59349	:douta	=	16'h	c429;
59350	:douta	=	16'h	bc09;
59351	:douta	=	16'h	bc09;
59352	:douta	=	16'h	bc09;
59353	:douta	=	16'h	bbe9;
59354	:douta	=	16'h	bc09;
59355	:douta	=	16'h	bc09;
59356	:douta	=	16'h	bbe9;
59357	:douta	=	16'h	bbe9;
59358	:douta	=	16'h	bc0a;
59359	:douta	=	16'h	b3e9;
59360	:douta	=	16'h	bbe9;
59361	:douta	=	16'h	b3e9;
59362	:douta	=	16'h	b3c9;
59363	:douta	=	16'h	bc09;
59364	:douta	=	16'h	b3e9;
59365	:douta	=	16'h	b3c9;
59366	:douta	=	16'h	b3c9;
59367	:douta	=	16'h	b3e9;
59368	:douta	=	16'h	b3c9;
59369	:douta	=	16'h	b3c9;
59370	:douta	=	16'h	b3c9;
59371	:douta	=	16'h	b3c9;
59372	:douta	=	16'h	b3c9;
59373	:douta	=	16'h	b3c9;
59374	:douta	=	16'h	abc9;
59375	:douta	=	16'h	aba9;
59376	:douta	=	16'h	abc9;
59377	:douta	=	16'h	aba9;
59378	:douta	=	16'h	abc9;
59379	:douta	=	16'h	aba9;
59380	:douta	=	16'h	aba9;
59381	:douta	=	16'h	aba9;
59382	:douta	=	16'h	ab89;
59383	:douta	=	16'h	aba8;
59384	:douta	=	16'h	aba8;
59385	:douta	=	16'h	aba9;
59386	:douta	=	16'h	ab89;
59387	:douta	=	16'h	aba9;
59388	:douta	=	16'h	a389;
59389	:douta	=	16'h	a389;
59390	:douta	=	16'h	ab89;
59391	:douta	=	16'h	a389;
59392	:douta	=	16'h	9cd5;
59393	:douta	=	16'h	8cb5;
59394	:douta	=	16'h	94d6;
59395	:douta	=	16'h	94b6;
59396	:douta	=	16'h	638f;
59397	:douta	=	16'h	2082;
59398	:douta	=	16'h	2903;
59399	:douta	=	16'h	2904;
59400	:douta	=	16'h	28e4;
59401	:douta	=	16'h	28e3;
59402	:douta	=	16'h	28e3;
59403	:douta	=	16'h	28e3;
59404	:douta	=	16'h	28e3;
59405	:douta	=	16'h	28e3;
59406	:douta	=	16'h	28e3;
59407	:douta	=	16'h	28e3;
59408	:douta	=	16'h	20e3;
59409	:douta	=	16'h	20e3;
59410	:douta	=	16'h	20e3;
59411	:douta	=	16'h	20e3;
59412	:douta	=	16'h	2904;
59413	:douta	=	16'h	20a2;
59414	:douta	=	16'h	20c2;
59415	:douta	=	16'h	20c2;
59416	:douta	=	16'h	20c2;
59417	:douta	=	16'h	20a2;
59418	:douta	=	16'h	28e3;
59419	:douta	=	16'h	28c3;
59420	:douta	=	16'h	28e3;
59421	:douta	=	16'h	28e3;
59422	:douta	=	16'h	28e3;
59423	:douta	=	16'h	3103;
59424	:douta	=	16'h	3103;
59425	:douta	=	16'h	3103;
59426	:douta	=	16'h	3923;
59427	:douta	=	16'h	3923;
59428	:douta	=	16'h	3943;
59429	:douta	=	16'h	4123;
59430	:douta	=	16'h	4143;
59431	:douta	=	16'h	4964;
59432	:douta	=	16'h	4964;
59433	:douta	=	16'h	5208;
59434	:douta	=	16'h	4a6a;
59435	:douta	=	16'h	0885;
59436	:douta	=	16'h	59c4;
59437	:douta	=	16'h	59c4;
59438	:douta	=	16'h	59c4;
59439	:douta	=	16'h	59e4;
59440	:douta	=	16'h	61e4;
59441	:douta	=	16'h	61e4;
59442	:douta	=	16'h	61e4;
59443	:douta	=	16'h	6a24;
59444	:douta	=	16'h	6a25;
59445	:douta	=	16'h	7224;
59446	:douta	=	16'h	72a8;
59447	:douta	=	16'h	a513;
59448	:douta	=	16'h	7204;
59449	:douta	=	16'h	7a84;
59450	:douta	=	16'h	7a85;
59451	:douta	=	16'h	82a5;
59452	:douta	=	16'h	7a85;
59453	:douta	=	16'h	82c6;
59454	:douta	=	16'h	82c6;
59455	:douta	=	16'h	82c6;
59456	:douta	=	16'h	8ac6;
59457	:douta	=	16'h	8ae6;
59458	:douta	=	16'h	8ac6;
59459	:douta	=	16'h	8ac6;
59460	:douta	=	16'h	8b06;
59461	:douta	=	16'h	92e6;
59462	:douta	=	16'h	9307;
59463	:douta	=	16'h	9326;
59464	:douta	=	16'h	9b27;
59465	:douta	=	16'h	9b47;
59466	:douta	=	16'h	9b27;
59467	:douta	=	16'h	92c4;
59468	:douta	=	16'h	f71a;
59469	:douta	=	16'h	73cc;
59470	:douta	=	16'h	4a28;
59471	:douta	=	16'h	0000;
59472	:douta	=	16'h	8b4a;
59473	:douta	=	16'h	94d0;
59474	:douta	=	16'h	59c3;
59475	:douta	=	16'h	b3a8;
59476	:douta	=	16'h	b3c7;
59477	:douta	=	16'h	b3c7;
59478	:douta	=	16'h	b3e7;
59479	:douta	=	16'h	b3c7;
59480	:douta	=	16'h	bbe8;
59481	:douta	=	16'h	bbe7;
59482	:douta	=	16'h	bc07;
59483	:douta	=	16'h	bc07;
59484	:douta	=	16'h	bc07;
59485	:douta	=	16'h	bc07;
59486	:douta	=	16'h	bc07;
59487	:douta	=	16'h	c428;
59488	:douta	=	16'h	c428;
59489	:douta	=	16'h	c428;
59490	:douta	=	16'h	c428;
59491	:douta	=	16'h	c428;
59492	:douta	=	16'h	c448;
59493	:douta	=	16'h	c448;
59494	:douta	=	16'h	c448;
59495	:douta	=	16'h	c448;
59496	:douta	=	16'h	c448;
59497	:douta	=	16'h	c448;
59498	:douta	=	16'h	cc49;
59499	:douta	=	16'h	cc49;
59500	:douta	=	16'h	cc49;
59501	:douta	=	16'h	c449;
59502	:douta	=	16'h	cc68;
59503	:douta	=	16'h	c448;
59504	:douta	=	16'h	cc68;
59505	:douta	=	16'h	cc68;
59506	:douta	=	16'h	cc68;
59507	:douta	=	16'h	cc67;
59508	:douta	=	16'h	cc68;
59509	:douta	=	16'h	cc68;
59510	:douta	=	16'h	cc68;
59511	:douta	=	16'h	cc48;
59512	:douta	=	16'h	cc69;
59513	:douta	=	16'h	cc68;
59514	:douta	=	16'h	cc68;
59515	:douta	=	16'h	cc68;
59516	:douta	=	16'h	cc68;
59517	:douta	=	16'h	cc69;
59518	:douta	=	16'h	cc69;
59519	:douta	=	16'h	cc69;
59520	:douta	=	16'h	cc69;
59521	:douta	=	16'h	cc68;
59522	:douta	=	16'h	cc69;
59523	:douta	=	16'h	cc69;
59524	:douta	=	16'h	cc69;
59525	:douta	=	16'h	cc89;
59526	:douta	=	16'h	cc89;
59527	:douta	=	16'h	cc69;
59528	:douta	=	16'h	cc89;
59529	:douta	=	16'h	cc89;
59530	:douta	=	16'h	cc89;
59531	:douta	=	16'h	cc8a;
59532	:douta	=	16'h	cc69;
59533	:douta	=	16'h	cc89;
59534	:douta	=	16'h	cc69;
59535	:douta	=	16'h	cc89;
59536	:douta	=	16'h	cc89;
59537	:douta	=	16'h	cc89;
59538	:douta	=	16'h	cc89;
59539	:douta	=	16'h	cc89;
59540	:douta	=	16'h	cc89;
59541	:douta	=	16'h	cc8a;
59542	:douta	=	16'h	cc89;
59543	:douta	=	16'h	cc8a;
59544	:douta	=	16'h	cc89;
59545	:douta	=	16'h	cc89;
59546	:douta	=	16'h	cc89;
59547	:douta	=	16'h	cc89;
59548	:douta	=	16'h	cc69;
59549	:douta	=	16'h	cc89;
59550	:douta	=	16'h	cc69;
59551	:douta	=	16'h	cc89;
59552	:douta	=	16'h	cc89;
59553	:douta	=	16'h	cc69;
59554	:douta	=	16'h	d488;
59555	:douta	=	16'h	ad74;
59556	:douta	=	16'h	e696;
59557	:douta	=	16'h	cc47;
59558	:douta	=	16'h	cc69;
59559	:douta	=	16'h	cc69;
59560	:douta	=	16'h	cc89;
59561	:douta	=	16'h	cc69;
59562	:douta	=	16'h	cc69;
59563	:douta	=	16'h	cc69;
59564	:douta	=	16'h	cc69;
59565	:douta	=	16'h	cc69;
59566	:douta	=	16'h	cc49;
59567	:douta	=	16'h	cc69;
59568	:douta	=	16'h	cc69;
59569	:douta	=	16'h	cc69;
59570	:douta	=	16'h	cc69;
59571	:douta	=	16'h	cc69;
59572	:douta	=	16'h	cc69;
59573	:douta	=	16'h	cc69;
59574	:douta	=	16'h	cc69;
59575	:douta	=	16'h	cc69;
59576	:douta	=	16'h	cc69;
59577	:douta	=	16'h	cc69;
59578	:douta	=	16'h	cc49;
59579	:douta	=	16'h	cc49;
59580	:douta	=	16'h	cc49;
59581	:douta	=	16'h	c449;
59582	:douta	=	16'h	cc49;
59583	:douta	=	16'h	cc69;
59584	:douta	=	16'h	c449;
59585	:douta	=	16'h	c449;
59586	:douta	=	16'h	c449;
59587	:douta	=	16'h	c449;
59588	:douta	=	16'h	c449;
59589	:douta	=	16'h	c449;
59590	:douta	=	16'h	c449;
59591	:douta	=	16'h	c449;
59592	:douta	=	16'h	c429;
59593	:douta	=	16'h	c429;
59594	:douta	=	16'h	c429;
59595	:douta	=	16'h	c449;
59596	:douta	=	16'h	c429;
59597	:douta	=	16'h	c429;
59598	:douta	=	16'h	c449;
59599	:douta	=	16'h	c429;
59600	:douta	=	16'h	bc29;
59601	:douta	=	16'h	c429;
59602	:douta	=	16'h	c429;
59603	:douta	=	16'h	bc29;
59604	:douta	=	16'h	bc29;
59605	:douta	=	16'h	bc09;
59606	:douta	=	16'h	bc09;
59607	:douta	=	16'h	bc09;
59608	:douta	=	16'h	bc29;
59609	:douta	=	16'h	bbe9;
59610	:douta	=	16'h	bc09;
59611	:douta	=	16'h	bbe9;
59612	:douta	=	16'h	bc09;
59613	:douta	=	16'h	bc09;
59614	:douta	=	16'h	bc09;
59615	:douta	=	16'h	bbe9;
59616	:douta	=	16'h	bc09;
59617	:douta	=	16'h	bbe9;
59618	:douta	=	16'h	b3e9;
59619	:douta	=	16'h	b3e9;
59620	:douta	=	16'h	b3c9;
59621	:douta	=	16'h	b3c9;
59622	:douta	=	16'h	b3c9;
59623	:douta	=	16'h	b3e9;
59624	:douta	=	16'h	b3e9;
59625	:douta	=	16'h	b3c9;
59626	:douta	=	16'h	b3e9;
59627	:douta	=	16'h	b3c9;
59628	:douta	=	16'h	b3c9;
59629	:douta	=	16'h	b3ca;
59630	:douta	=	16'h	b3a9;
59631	:douta	=	16'h	abc9;
59632	:douta	=	16'h	aba9;
59633	:douta	=	16'h	aba9;
59634	:douta	=	16'h	b3c9;
59635	:douta	=	16'h	aba9;
59636	:douta	=	16'h	aba9;
59637	:douta	=	16'h	ab89;
59638	:douta	=	16'h	aba9;
59639	:douta	=	16'h	aba9;
59640	:douta	=	16'h	abc9;
59641	:douta	=	16'h	aba9;
59642	:douta	=	16'h	ab89;
59643	:douta	=	16'h	aba9;
59644	:douta	=	16'h	a389;
59645	:douta	=	16'h	ab89;
59646	:douta	=	16'h	a389;
59647	:douta	=	16'h	a388;
59648	:douta	=	16'h	8c54;
59649	:douta	=	16'h	94b6;
59650	:douta	=	16'h	94d6;
59651	:douta	=	16'h	8496;
59652	:douta	=	16'h	39c7;
59653	:douta	=	16'h	2082;
59654	:douta	=	16'h	2904;
59655	:douta	=	16'h	28e3;
59656	:douta	=	16'h	28e3;
59657	:douta	=	16'h	28e3;
59658	:douta	=	16'h	28e3;
59659	:douta	=	16'h	28e3;
59660	:douta	=	16'h	28e3;
59661	:douta	=	16'h	28e3;
59662	:douta	=	16'h	20c3;
59663	:douta	=	16'h	20e3;
59664	:douta	=	16'h	20e3;
59665	:douta	=	16'h	20e3;
59666	:douta	=	16'h	20c3;
59667	:douta	=	16'h	20e3;
59668	:douta	=	16'h	20e3;
59669	:douta	=	16'h	20a2;
59670	:douta	=	16'h	20a2;
59671	:douta	=	16'h	20c2;
59672	:douta	=	16'h	20c2;
59673	:douta	=	16'h	28c3;
59674	:douta	=	16'h	28e3;
59675	:douta	=	16'h	28e3;
59676	:douta	=	16'h	28e3;
59677	:douta	=	16'h	3103;
59678	:douta	=	16'h	3103;
59679	:douta	=	16'h	30e3;
59680	:douta	=	16'h	3103;
59681	:douta	=	16'h	3103;
59682	:douta	=	16'h	3923;
59683	:douta	=	16'h	3923;
59684	:douta	=	16'h	4124;
59685	:douta	=	16'h	4143;
59686	:douta	=	16'h	4143;
59687	:douta	=	16'h	4964;
59688	:douta	=	16'h	4964;
59689	:douta	=	16'h	524a;
59690	:douta	=	16'h	4a49;
59691	:douta	=	16'h	1084;
59692	:douta	=	16'h	59c4;
59693	:douta	=	16'h	61c4;
59694	:douta	=	16'h	59c4;
59695	:douta	=	16'h	59c4;
59696	:douta	=	16'h	61e4;
59697	:douta	=	16'h	6204;
59698	:douta	=	16'h	6a04;
59699	:douta	=	16'h	6a24;
59700	:douta	=	16'h	6a24;
59701	:douta	=	16'h	7224;
59702	:douta	=	16'h	7b6c;
59703	:douta	=	16'h	b593;
59704	:douta	=	16'h	7203;
59705	:douta	=	16'h	7a64;
59706	:douta	=	16'h	7a85;
59707	:douta	=	16'h	7a85;
59708	:douta	=	16'h	82a5;
59709	:douta	=	16'h	82a5;
59710	:douta	=	16'h	82a6;
59711	:douta	=	16'h	82c6;
59712	:douta	=	16'h	8ac6;
59713	:douta	=	16'h	8ae7;
59714	:douta	=	16'h	8ac6;
59715	:douta	=	16'h	8ae7;
59716	:douta	=	16'h	8ae6;
59717	:douta	=	16'h	9307;
59718	:douta	=	16'h	9307;
59719	:douta	=	16'h	9326;
59720	:douta	=	16'h	9b27;
59721	:douta	=	16'h	9b47;
59722	:douta	=	16'h	9b27;
59723	:douta	=	16'h	9b46;
59724	:douta	=	16'h	eef9;
59725	:douta	=	16'h	8caf;
59726	:douta	=	16'h	0000;
59727	:douta	=	16'h	7b8a;
59728	:douta	=	16'h	e696;
59729	:douta	=	16'h	7bad;
59730	:douta	=	16'h	71c3;
59731	:douta	=	16'h	b3c7;
59732	:douta	=	16'h	b3c7;
59733	:douta	=	16'h	b3c8;
59734	:douta	=	16'h	b3c7;
59735	:douta	=	16'h	bc08;
59736	:douta	=	16'h	b3e8;
59737	:douta	=	16'h	bc07;
59738	:douta	=	16'h	bbe7;
59739	:douta	=	16'h	bc07;
59740	:douta	=	16'h	bc08;
59741	:douta	=	16'h	bc07;
59742	:douta	=	16'h	bc07;
59743	:douta	=	16'h	c428;
59744	:douta	=	16'h	c428;
59745	:douta	=	16'h	c428;
59746	:douta	=	16'h	c428;
59747	:douta	=	16'h	c428;
59748	:douta	=	16'h	c428;
59749	:douta	=	16'h	c448;
59750	:douta	=	16'h	c448;
59751	:douta	=	16'h	c428;
59752	:douta	=	16'h	c448;
59753	:douta	=	16'h	c448;
59754	:douta	=	16'h	c448;
59755	:douta	=	16'h	c448;
59756	:douta	=	16'h	c449;
59757	:douta	=	16'h	cc68;
59758	:douta	=	16'h	cc68;
59759	:douta	=	16'h	c448;
59760	:douta	=	16'h	c448;
59761	:douta	=	16'h	cc68;
59762	:douta	=	16'h	c448;
59763	:douta	=	16'h	cc68;
59764	:douta	=	16'h	cc68;
59765	:douta	=	16'h	cc68;
59766	:douta	=	16'h	cc68;
59767	:douta	=	16'h	cc69;
59768	:douta	=	16'h	cc68;
59769	:douta	=	16'h	cc68;
59770	:douta	=	16'h	cc69;
59771	:douta	=	16'h	cc89;
59772	:douta	=	16'h	cc68;
59773	:douta	=	16'h	cc69;
59774	:douta	=	16'h	cc69;
59775	:douta	=	16'h	cc69;
59776	:douta	=	16'h	cc69;
59777	:douta	=	16'h	cc69;
59778	:douta	=	16'h	d489;
59779	:douta	=	16'h	cc69;
59780	:douta	=	16'h	cc69;
59781	:douta	=	16'h	cc69;
59782	:douta	=	16'h	cc69;
59783	:douta	=	16'h	cc89;
59784	:douta	=	16'h	cc69;
59785	:douta	=	16'h	cc89;
59786	:douta	=	16'h	cc69;
59787	:douta	=	16'h	cc89;
59788	:douta	=	16'h	cc8a;
59789	:douta	=	16'h	cc89;
59790	:douta	=	16'h	cc89;
59791	:douta	=	16'h	cc89;
59792	:douta	=	16'h	cc89;
59793	:douta	=	16'h	cc89;
59794	:douta	=	16'h	cc89;
59795	:douta	=	16'h	cc89;
59796	:douta	=	16'h	cc89;
59797	:douta	=	16'h	cc89;
59798	:douta	=	16'h	cc89;
59799	:douta	=	16'h	cc89;
59800	:douta	=	16'h	cc89;
59801	:douta	=	16'h	cc89;
59802	:douta	=	16'h	cc89;
59803	:douta	=	16'h	cc89;
59804	:douta	=	16'h	d489;
59805	:douta	=	16'h	cc69;
59806	:douta	=	16'h	cc69;
59807	:douta	=	16'h	cc69;
59808	:douta	=	16'h	cc69;
59809	:douta	=	16'h	cc69;
59810	:douta	=	16'h	d467;
59811	:douta	=	16'h	b594;
59812	:douta	=	16'h	e696;
59813	:douta	=	16'h	cc48;
59814	:douta	=	16'h	cc69;
59815	:douta	=	16'h	cc69;
59816	:douta	=	16'h	cc8a;
59817	:douta	=	16'h	cc69;
59818	:douta	=	16'h	cc69;
59819	:douta	=	16'h	cc69;
59820	:douta	=	16'h	cc69;
59821	:douta	=	16'h	cc69;
59822	:douta	=	16'h	cc89;
59823	:douta	=	16'h	cc69;
59824	:douta	=	16'h	cc69;
59825	:douta	=	16'h	cc69;
59826	:douta	=	16'h	cc69;
59827	:douta	=	16'h	cc69;
59828	:douta	=	16'h	cc69;
59829	:douta	=	16'h	cc49;
59830	:douta	=	16'h	cc69;
59831	:douta	=	16'h	cc69;
59832	:douta	=	16'h	cc69;
59833	:douta	=	16'h	cc49;
59834	:douta	=	16'h	cc69;
59835	:douta	=	16'h	cc49;
59836	:douta	=	16'h	cc49;
59837	:douta	=	16'h	cc49;
59838	:douta	=	16'h	cc49;
59839	:douta	=	16'h	cc69;
59840	:douta	=	16'h	cc49;
59841	:douta	=	16'h	cc69;
59842	:douta	=	16'h	cc49;
59843	:douta	=	16'h	c449;
59844	:douta	=	16'h	c449;
59845	:douta	=	16'h	c449;
59846	:douta	=	16'h	c429;
59847	:douta	=	16'h	c429;
59848	:douta	=	16'h	c449;
59849	:douta	=	16'h	c429;
59850	:douta	=	16'h	c429;
59851	:douta	=	16'h	c429;
59852	:douta	=	16'h	c449;
59853	:douta	=	16'h	bc29;
59854	:douta	=	16'h	c429;
59855	:douta	=	16'h	c429;
59856	:douta	=	16'h	bc29;
59857	:douta	=	16'h	c429;
59858	:douta	=	16'h	bc29;
59859	:douta	=	16'h	bc29;
59860	:douta	=	16'h	bc09;
59861	:douta	=	16'h	bc09;
59862	:douta	=	16'h	bc09;
59863	:douta	=	16'h	bc29;
59864	:douta	=	16'h	bc09;
59865	:douta	=	16'h	bc09;
59866	:douta	=	16'h	bc09;
59867	:douta	=	16'h	bc09;
59868	:douta	=	16'h	bc09;
59869	:douta	=	16'h	bc09;
59870	:douta	=	16'h	bc09;
59871	:douta	=	16'h	bbe9;
59872	:douta	=	16'h	bbe9;
59873	:douta	=	16'h	bbe9;
59874	:douta	=	16'h	bc09;
59875	:douta	=	16'h	b3e9;
59876	:douta	=	16'h	b3e9;
59877	:douta	=	16'h	b3c9;
59878	:douta	=	16'h	b3c9;
59879	:douta	=	16'h	b3c9;
59880	:douta	=	16'h	b3c9;
59881	:douta	=	16'h	b3e9;
59882	:douta	=	16'h	b3c9;
59883	:douta	=	16'h	b3c9;
59884	:douta	=	16'h	b3c8;
59885	:douta	=	16'h	b3c9;
59886	:douta	=	16'h	b3ca;
59887	:douta	=	16'h	b3c9;
59888	:douta	=	16'h	b3c9;
59889	:douta	=	16'h	aba9;
59890	:douta	=	16'h	aba9;
59891	:douta	=	16'h	aba9;
59892	:douta	=	16'h	abc9;
59893	:douta	=	16'h	aba9;
59894	:douta	=	16'h	aba9;
59895	:douta	=	16'h	aba9;
59896	:douta	=	16'h	aba8;
59897	:douta	=	16'h	aba9;
59898	:douta	=	16'h	a388;
59899	:douta	=	16'h	a389;
59900	:douta	=	16'h	a389;
59901	:douta	=	16'h	a389;
59902	:douta	=	16'h	a388;
59903	:douta	=	16'h	a389;
59904	:douta	=	16'h	8c54;
59905	:douta	=	16'h	8c95;
59906	:douta	=	16'h	94b6;
59907	:douta	=	16'h	8cf7;
59908	:douta	=	16'h	20e3;
59909	:douta	=	16'h	28e3;
59910	:douta	=	16'h	2904;
59911	:douta	=	16'h	28e3;
59912	:douta	=	16'h	28e3;
59913	:douta	=	16'h	20e3;
59914	:douta	=	16'h	28e3;
59915	:douta	=	16'h	28e3;
59916	:douta	=	16'h	28e3;
59917	:douta	=	16'h	28e3;
59918	:douta	=	16'h	20e3;
59919	:douta	=	16'h	20e3;
59920	:douta	=	16'h	20e3;
59921	:douta	=	16'h	20e3;
59922	:douta	=	16'h	20e3;
59923	:douta	=	16'h	20e3;
59924	:douta	=	16'h	20e3;
59925	:douta	=	16'h	20a2;
59926	:douta	=	16'h	20a2;
59927	:douta	=	16'h	20c2;
59928	:douta	=	16'h	20c3;
59929	:douta	=	16'h	20c2;
59930	:douta	=	16'h	28c3;
59931	:douta	=	16'h	28e3;
59932	:douta	=	16'h	28e3;
59933	:douta	=	16'h	30e3;
59934	:douta	=	16'h	30e3;
59935	:douta	=	16'h	3103;
59936	:douta	=	16'h	3103;
59937	:douta	=	16'h	3103;
59938	:douta	=	16'h	3923;
59939	:douta	=	16'h	3923;
59940	:douta	=	16'h	4124;
59941	:douta	=	16'h	4164;
59942	:douta	=	16'h	4143;
59943	:douta	=	16'h	4964;
59944	:douta	=	16'h	4964;
59945	:douta	=	16'h	5a8b;
59946	:douta	=	16'h	39c8;
59947	:douta	=	16'h	18a4;
59948	:douta	=	16'h	59c4;
59949	:douta	=	16'h	59c4;
59950	:douta	=	16'h	59e4;
59951	:douta	=	16'h	59c4;
59952	:douta	=	16'h	61e4;
59953	:douta	=	16'h	6204;
59954	:douta	=	16'h	6a04;
59955	:douta	=	16'h	6a24;
59956	:douta	=	16'h	6a24;
59957	:douta	=	16'h	7244;
59958	:douta	=	16'h	83ee;
59959	:douta	=	16'h	b573;
59960	:douta	=	16'h	7203;
59961	:douta	=	16'h	7a85;
59962	:douta	=	16'h	7a85;
59963	:douta	=	16'h	7a85;
59964	:douta	=	16'h	7a85;
59965	:douta	=	16'h	82a6;
59966	:douta	=	16'h	82c6;
59967	:douta	=	16'h	82c6;
59968	:douta	=	16'h	8ac6;
59969	:douta	=	16'h	8ac6;
59970	:douta	=	16'h	8ae6;
59971	:douta	=	16'h	8ae6;
59972	:douta	=	16'h	8ae7;
59973	:douta	=	16'h	9307;
59974	:douta	=	16'h	9307;
59975	:douta	=	16'h	9b27;
59976	:douta	=	16'h	9b47;
59977	:douta	=	16'h	9b47;
59978	:douta	=	16'h	9306;
59979	:douta	=	16'h	a387;
59980	:douta	=	16'h	de37;
59981	:douta	=	16'h	d675;
59982	:douta	=	16'h	5269;
59983	:douta	=	16'h	de96;
59984	:douta	=	16'h	de55;
59985	:douta	=	16'h	732a;
59986	:douta	=	16'h	79e2;
59987	:douta	=	16'h	b3c8;
59988	:douta	=	16'h	aba7;
59989	:douta	=	16'h	b3c7;
59990	:douta	=	16'h	b3e8;
59991	:douta	=	16'h	b3e7;
59992	:douta	=	16'h	bbe8;
59993	:douta	=	16'h	bbe7;
59994	:douta	=	16'h	bc07;
59995	:douta	=	16'h	bc07;
59996	:douta	=	16'h	bc08;
59997	:douta	=	16'h	bc07;
59998	:douta	=	16'h	c407;
59999	:douta	=	16'h	c407;
60000	:douta	=	16'h	bc07;
60001	:douta	=	16'h	c428;
60002	:douta	=	16'h	c448;
60003	:douta	=	16'h	c428;
60004	:douta	=	16'h	c448;
60005	:douta	=	16'h	c448;
60006	:douta	=	16'h	c448;
60007	:douta	=	16'h	c448;
60008	:douta	=	16'h	c448;
60009	:douta	=	16'h	c448;
60010	:douta	=	16'h	c448;
60011	:douta	=	16'h	c449;
60012	:douta	=	16'h	cc49;
60013	:douta	=	16'h	cc49;
60014	:douta	=	16'h	c448;
60015	:douta	=	16'h	c448;
60016	:douta	=	16'h	cc68;
60017	:douta	=	16'h	cc68;
60018	:douta	=	16'h	cc68;
60019	:douta	=	16'h	cc68;
60020	:douta	=	16'h	cc68;
60021	:douta	=	16'h	cc69;
60022	:douta	=	16'h	cc69;
60023	:douta	=	16'h	cc68;
60024	:douta	=	16'h	cc69;
60025	:douta	=	16'h	cc68;
60026	:douta	=	16'h	cc68;
60027	:douta	=	16'h	cc69;
60028	:douta	=	16'h	cc69;
60029	:douta	=	16'h	cc69;
60030	:douta	=	16'h	cc69;
60031	:douta	=	16'h	cc68;
60032	:douta	=	16'h	cc69;
60033	:douta	=	16'h	cc69;
60034	:douta	=	16'h	cc69;
60035	:douta	=	16'h	cc69;
60036	:douta	=	16'h	cc69;
60037	:douta	=	16'h	cc69;
60038	:douta	=	16'h	cc89;
60039	:douta	=	16'h	cc69;
60040	:douta	=	16'h	cc89;
60041	:douta	=	16'h	cc69;
60042	:douta	=	16'h	cc89;
60043	:douta	=	16'h	cc89;
60044	:douta	=	16'h	cc89;
60045	:douta	=	16'h	cc89;
60046	:douta	=	16'h	cc69;
60047	:douta	=	16'h	cc89;
60048	:douta	=	16'h	cc89;
60049	:douta	=	16'h	cc89;
60050	:douta	=	16'h	cc89;
60051	:douta	=	16'h	cc89;
60052	:douta	=	16'h	cc8a;
60053	:douta	=	16'h	cc89;
60054	:douta	=	16'h	cc89;
60055	:douta	=	16'h	cc89;
60056	:douta	=	16'h	cc89;
60057	:douta	=	16'h	cc89;
60058	:douta	=	16'h	cc69;
60059	:douta	=	16'h	cc69;
60060	:douta	=	16'h	cc89;
60061	:douta	=	16'h	cc69;
60062	:douta	=	16'h	cc69;
60063	:douta	=	16'h	cc69;
60064	:douta	=	16'h	cc69;
60065	:douta	=	16'h	cc69;
60066	:douta	=	16'h	d488;
60067	:douta	=	16'h	b594;
60068	:douta	=	16'h	de76;
60069	:douta	=	16'h	cc48;
60070	:douta	=	16'h	cc69;
60071	:douta	=	16'h	cc69;
60072	:douta	=	16'h	cc69;
60073	:douta	=	16'h	cc69;
60074	:douta	=	16'h	cc69;
60075	:douta	=	16'h	cc69;
60076	:douta	=	16'h	cc69;
60077	:douta	=	16'h	cc69;
60078	:douta	=	16'h	cc69;
60079	:douta	=	16'h	cc69;
60080	:douta	=	16'h	cc69;
60081	:douta	=	16'h	cc69;
60082	:douta	=	16'h	cc69;
60083	:douta	=	16'h	cc69;
60084	:douta	=	16'h	cc69;
60085	:douta	=	16'h	cc69;
60086	:douta	=	16'h	cc6a;
60087	:douta	=	16'h	cc69;
60088	:douta	=	16'h	cc69;
60089	:douta	=	16'h	cc49;
60090	:douta	=	16'h	cc69;
60091	:douta	=	16'h	c449;
60092	:douta	=	16'h	c449;
60093	:douta	=	16'h	cc49;
60094	:douta	=	16'h	c449;
60095	:douta	=	16'h	c448;
60096	:douta	=	16'h	c449;
60097	:douta	=	16'h	cc49;
60098	:douta	=	16'h	cc49;
60099	:douta	=	16'h	c449;
60100	:douta	=	16'h	c449;
60101	:douta	=	16'h	c449;
60102	:douta	=	16'h	c429;
60103	:douta	=	16'h	c429;
60104	:douta	=	16'h	c429;
60105	:douta	=	16'h	c449;
60106	:douta	=	16'h	c429;
60107	:douta	=	16'h	c429;
60108	:douta	=	16'h	c449;
60109	:douta	=	16'h	c429;
60110	:douta	=	16'h	c429;
60111	:douta	=	16'h	c429;
60112	:douta	=	16'h	c429;
60113	:douta	=	16'h	bc29;
60114	:douta	=	16'h	bc09;
60115	:douta	=	16'h	bc09;
60116	:douta	=	16'h	bc09;
60117	:douta	=	16'h	c429;
60118	:douta	=	16'h	c429;
60119	:douta	=	16'h	bc09;
60120	:douta	=	16'h	bc09;
60121	:douta	=	16'h	bc09;
60122	:douta	=	16'h	bc09;
60123	:douta	=	16'h	bc09;
60124	:douta	=	16'h	bc09;
60125	:douta	=	16'h	bc09;
60126	:douta	=	16'h	bc09;
60127	:douta	=	16'h	bbe9;
60128	:douta	=	16'h	bbe9;
60129	:douta	=	16'h	b3e9;
60130	:douta	=	16'h	b3e9;
60131	:douta	=	16'h	bbe9;
60132	:douta	=	16'h	b3e9;
60133	:douta	=	16'h	b3e9;
60134	:douta	=	16'h	b3e9;
60135	:douta	=	16'h	b3c9;
60136	:douta	=	16'h	bbe9;
60137	:douta	=	16'h	b3c9;
60138	:douta	=	16'h	b3e9;
60139	:douta	=	16'h	b3c9;
60140	:douta	=	16'h	b3c8;
60141	:douta	=	16'h	b3c9;
60142	:douta	=	16'h	b3a9;
60143	:douta	=	16'h	b3ca;
60144	:douta	=	16'h	aba9;
60145	:douta	=	16'h	aba9;
60146	:douta	=	16'h	aba9;
60147	:douta	=	16'h	aba9;
60148	:douta	=	16'h	b3c9;
60149	:douta	=	16'h	aba9;
60150	:douta	=	16'h	aba9;
60151	:douta	=	16'h	aba9;
60152	:douta	=	16'h	aba9;
60153	:douta	=	16'h	aba8;
60154	:douta	=	16'h	a388;
60155	:douta	=	16'h	a389;
60156	:douta	=	16'h	a389;
60157	:douta	=	16'h	ab89;
60158	:douta	=	16'h	a389;
60159	:douta	=	16'h	a389;
60160	:douta	=	16'h	8c95;
60161	:douta	=	16'h	94b5;
60162	:douta	=	16'h	94b6;
60163	:douta	=	16'h	9518;
60164	:douta	=	16'h	2061;
60165	:douta	=	16'h	2903;
60166	:douta	=	16'h	3104;
60167	:douta	=	16'h	28e3;
60168	:douta	=	16'h	28e3;
60169	:douta	=	16'h	28e3;
60170	:douta	=	16'h	20e3;
60171	:douta	=	16'h	28e3;
60172	:douta	=	16'h	28e3;
60173	:douta	=	16'h	20e3;
60174	:douta	=	16'h	20e3;
60175	:douta	=	16'h	20e3;
60176	:douta	=	16'h	28e3;
60177	:douta	=	16'h	20e3;
60178	:douta	=	16'h	20c3;
60179	:douta	=	16'h	28e3;
60180	:douta	=	16'h	18a2;
60181	:douta	=	16'h	20c3;
60182	:douta	=	16'h	20a2;
60183	:douta	=	16'h	20c3;
60184	:douta	=	16'h	20c2;
60185	:douta	=	16'h	28c3;
60186	:douta	=	16'h	28c3;
60187	:douta	=	16'h	28e3;
60188	:douta	=	16'h	28e3;
60189	:douta	=	16'h	3103;
60190	:douta	=	16'h	3103;
60191	:douta	=	16'h	3103;
60192	:douta	=	16'h	3123;
60193	:douta	=	16'h	3103;
60194	:douta	=	16'h	3943;
60195	:douta	=	16'h	3923;
60196	:douta	=	16'h	4144;
60197	:douta	=	16'h	4143;
60198	:douta	=	16'h	4163;
60199	:douta	=	16'h	4964;
60200	:douta	=	16'h	4964;
60201	:douta	=	16'h	528b;
60202	:douta	=	16'h	2967;
60203	:douta	=	16'h	3104;
60204	:douta	=	16'h	59c4;
60205	:douta	=	16'h	59c4;
60206	:douta	=	16'h	59e4;
60207	:douta	=	16'h	61e4;
60208	:douta	=	16'h	61e4;
60209	:douta	=	16'h	6a24;
60210	:douta	=	16'h	6a24;
60211	:douta	=	16'h	7245;
60212	:douta	=	16'h	7224;
60213	:douta	=	16'h	7223;
60214	:douta	=	16'h	9cf2;
60215	:douta	=	16'h	acf0;
60216	:douta	=	16'h	7a64;
60217	:douta	=	16'h	7a85;
60218	:douta	=	16'h	7a85;
60219	:douta	=	16'h	7a85;
60220	:douta	=	16'h	82a5;
60221	:douta	=	16'h	82a6;
60222	:douta	=	16'h	82c6;
60223	:douta	=	16'h	82c6;
60224	:douta	=	16'h	8ac6;
60225	:douta	=	16'h	8ac6;
60226	:douta	=	16'h	8ac6;
60227	:douta	=	16'h	8ae6;
60228	:douta	=	16'h	92e6;
60229	:douta	=	16'h	9307;
60230	:douta	=	16'h	9307;
60231	:douta	=	16'h	9b27;
60232	:douta	=	16'h	9b47;
60233	:douta	=	16'h	9b47;
60234	:douta	=	16'h	92c6;
60235	:douta	=	16'h	ac4b;
60236	:douta	=	16'h	e6d7;
60237	:douta	=	16'h	acb0;
60238	:douta	=	16'h	29e7;
60239	:douta	=	16'h	b44e;
60240	:douta	=	16'h	eef8;
60241	:douta	=	16'h	5a47;
60242	:douta	=	16'h	9ae4;
60243	:douta	=	16'h	aba7;
60244	:douta	=	16'h	aba7;
60245	:douta	=	16'h	b3c7;
60246	:douta	=	16'h	b3e7;
60247	:douta	=	16'h	bbe8;
60248	:douta	=	16'h	b3e7;
60249	:douta	=	16'h	bbe7;
60250	:douta	=	16'h	bc07;
60251	:douta	=	16'h	bc08;
60252	:douta	=	16'h	bc08;
60253	:douta	=	16'h	c407;
60254	:douta	=	16'h	c407;
60255	:douta	=	16'h	c407;
60256	:douta	=	16'h	c428;
60257	:douta	=	16'h	c448;
60258	:douta	=	16'h	c428;
60259	:douta	=	16'h	c448;
60260	:douta	=	16'h	c428;
60261	:douta	=	16'h	c448;
60262	:douta	=	16'h	c448;
60263	:douta	=	16'h	cc49;
60264	:douta	=	16'h	c448;
60265	:douta	=	16'h	c428;
60266	:douta	=	16'h	c448;
60267	:douta	=	16'h	c449;
60268	:douta	=	16'h	c448;
60269	:douta	=	16'h	cc49;
60270	:douta	=	16'h	c448;
60271	:douta	=	16'h	c448;
60272	:douta	=	16'h	c448;
60273	:douta	=	16'h	cc68;
60274	:douta	=	16'h	cc68;
60275	:douta	=	16'h	cc68;
60276	:douta	=	16'h	cc68;
60277	:douta	=	16'h	cc68;
60278	:douta	=	16'h	cc68;
60279	:douta	=	16'h	cc68;
60280	:douta	=	16'h	cc68;
60281	:douta	=	16'h	cc68;
60282	:douta	=	16'h	cc69;
60283	:douta	=	16'h	cc69;
60284	:douta	=	16'h	cc69;
60285	:douta	=	16'h	cc69;
60286	:douta	=	16'h	cc69;
60287	:douta	=	16'h	cc69;
60288	:douta	=	16'h	cc69;
60289	:douta	=	16'h	cc69;
60290	:douta	=	16'h	cc69;
60291	:douta	=	16'h	cc69;
60292	:douta	=	16'h	cc69;
60293	:douta	=	16'h	cc89;
60294	:douta	=	16'h	cc69;
60295	:douta	=	16'h	cc89;
60296	:douta	=	16'h	cc69;
60297	:douta	=	16'h	cc89;
60298	:douta	=	16'h	cc89;
60299	:douta	=	16'h	cc89;
60300	:douta	=	16'h	cc89;
60301	:douta	=	16'h	cc89;
60302	:douta	=	16'h	cc89;
60303	:douta	=	16'h	cc89;
60304	:douta	=	16'h	cc89;
60305	:douta	=	16'h	cc89;
60306	:douta	=	16'h	cc89;
60307	:douta	=	16'h	cc69;
60308	:douta	=	16'h	cc89;
60309	:douta	=	16'h	cc89;
60310	:douta	=	16'h	cc89;
60311	:douta	=	16'h	cc89;
60312	:douta	=	16'h	cc69;
60313	:douta	=	16'h	cc89;
60314	:douta	=	16'h	cc89;
60315	:douta	=	16'h	cc69;
60316	:douta	=	16'h	cc89;
60317	:douta	=	16'h	cc89;
60318	:douta	=	16'h	cc69;
60319	:douta	=	16'h	cc69;
60320	:douta	=	16'h	cc69;
60321	:douta	=	16'h	cc69;
60322	:douta	=	16'h	cc68;
60323	:douta	=	16'h	b594;
60324	:douta	=	16'h	e696;
60325	:douta	=	16'h	cc48;
60326	:douta	=	16'h	cc89;
60327	:douta	=	16'h	cc69;
60328	:douta	=	16'h	cc69;
60329	:douta	=	16'h	cc69;
60330	:douta	=	16'h	cc69;
60331	:douta	=	16'h	cc69;
60332	:douta	=	16'h	cc69;
60333	:douta	=	16'h	cc69;
60334	:douta	=	16'h	cc69;
60335	:douta	=	16'h	cc69;
60336	:douta	=	16'h	cc69;
60337	:douta	=	16'h	cc69;
60338	:douta	=	16'h	cc69;
60339	:douta	=	16'h	cc69;
60340	:douta	=	16'h	cc69;
60341	:douta	=	16'h	cc8a;
60342	:douta	=	16'h	cc69;
60343	:douta	=	16'h	cc69;
60344	:douta	=	16'h	cc69;
60345	:douta	=	16'h	c449;
60346	:douta	=	16'h	cc69;
60347	:douta	=	16'h	cc69;
60348	:douta	=	16'h	cc49;
60349	:douta	=	16'h	c449;
60350	:douta	=	16'h	cc69;
60351	:douta	=	16'h	c449;
60352	:douta	=	16'h	cc69;
60353	:douta	=	16'h	c449;
60354	:douta	=	16'h	c449;
60355	:douta	=	16'h	c449;
60356	:douta	=	16'h	c449;
60357	:douta	=	16'h	c429;
60358	:douta	=	16'h	c429;
60359	:douta	=	16'h	c429;
60360	:douta	=	16'h	c449;
60361	:douta	=	16'h	c429;
60362	:douta	=	16'h	c429;
60363	:douta	=	16'h	c429;
60364	:douta	=	16'h	c429;
60365	:douta	=	16'h	c429;
60366	:douta	=	16'h	c429;
60367	:douta	=	16'h	c429;
60368	:douta	=	16'h	c429;
60369	:douta	=	16'h	c429;
60370	:douta	=	16'h	bc09;
60371	:douta	=	16'h	bc29;
60372	:douta	=	16'h	bc29;
60373	:douta	=	16'h	bc29;
60374	:douta	=	16'h	bc09;
60375	:douta	=	16'h	bc09;
60376	:douta	=	16'h	bc09;
60377	:douta	=	16'h	bc2a;
60378	:douta	=	16'h	bc09;
60379	:douta	=	16'h	bc09;
60380	:douta	=	16'h	bc09;
60381	:douta	=	16'h	bc09;
60382	:douta	=	16'h	bbe9;
60383	:douta	=	16'h	bc09;
60384	:douta	=	16'h	bc09;
60385	:douta	=	16'h	bc09;
60386	:douta	=	16'h	bbe9;
60387	:douta	=	16'h	bbe9;
60388	:douta	=	16'h	bbe9;
60389	:douta	=	16'h	b3e9;
60390	:douta	=	16'h	b3e9;
60391	:douta	=	16'h	b3e9;
60392	:douta	=	16'h	b3e9;
60393	:douta	=	16'h	b3e9;
60394	:douta	=	16'h	b3c9;
60395	:douta	=	16'h	b3c9;
60396	:douta	=	16'h	b3c9;
60397	:douta	=	16'h	abc9;
60398	:douta	=	16'h	aba9;
60399	:douta	=	16'h	aba9;
60400	:douta	=	16'h	abc9;
60401	:douta	=	16'h	abc9;
60402	:douta	=	16'h	aba9;
60403	:douta	=	16'h	aba9;
60404	:douta	=	16'h	aba9;
60405	:douta	=	16'h	aba9;
60406	:douta	=	16'h	abc9;
60407	:douta	=	16'h	aba9;
60408	:douta	=	16'h	aba9;
60409	:douta	=	16'h	aba9;
60410	:douta	=	16'h	aba9;
60411	:douta	=	16'h	aba9;
60412	:douta	=	16'h	a389;
60413	:douta	=	16'h	a389;
60414	:douta	=	16'h	a389;
60415	:douta	=	16'h	a389;
60416	:douta	=	16'h	8c95;
60417	:douta	=	16'h	94d6;
60418	:douta	=	16'h	8c96;
60419	:douta	=	16'h	8495;
60420	:douta	=	16'h	20a2;
60421	:douta	=	16'h	2904;
60422	:douta	=	16'h	2904;
60423	:douta	=	16'h	20e3;
60424	:douta	=	16'h	2904;
60425	:douta	=	16'h	28e3;
60426	:douta	=	16'h	28e3;
60427	:douta	=	16'h	28e3;
60428	:douta	=	16'h	28e3;
60429	:douta	=	16'h	2904;
60430	:douta	=	16'h	20e3;
60431	:douta	=	16'h	20e3;
60432	:douta	=	16'h	20e3;
60433	:douta	=	16'h	20e3;
60434	:douta	=	16'h	20c3;
60435	:douta	=	16'h	28e3;
60436	:douta	=	16'h	18a2;
60437	:douta	=	16'h	20a3;
60438	:douta	=	16'h	20a2;
60439	:douta	=	16'h	20c2;
60440	:douta	=	16'h	28c3;
60441	:douta	=	16'h	28e3;
60442	:douta	=	16'h	28e3;
60443	:douta	=	16'h	28e3;
60444	:douta	=	16'h	28e3;
60445	:douta	=	16'h	3103;
60446	:douta	=	16'h	30e3;
60447	:douta	=	16'h	3103;
60448	:douta	=	16'h	3103;
60449	:douta	=	16'h	3903;
60450	:douta	=	16'h	3923;
60451	:douta	=	16'h	3943;
60452	:douta	=	16'h	4164;
60453	:douta	=	16'h	4164;
60454	:douta	=	16'h	4163;
60455	:douta	=	16'h	4964;
60456	:douta	=	16'h	4144;
60457	:douta	=	16'h	528a;
60458	:douta	=	16'h	2967;
60459	:douta	=	16'h	3924;
60460	:douta	=	16'h	59c4;
60461	:douta	=	16'h	59c4;
60462	:douta	=	16'h	59e4;
60463	:douta	=	16'h	61e4;
60464	:douta	=	16'h	61e4;
60465	:douta	=	16'h	6a24;
60466	:douta	=	16'h	6a24;
60467	:douta	=	16'h	6a25;
60468	:douta	=	16'h	7245;
60469	:douta	=	16'h	7204;
60470	:douta	=	16'h	a553;
60471	:douta	=	16'h	a4af;
60472	:douta	=	16'h	7a64;
60473	:douta	=	16'h	7a85;
60474	:douta	=	16'h	7a85;
60475	:douta	=	16'h	82a5;
60476	:douta	=	16'h	82a5;
60477	:douta	=	16'h	82a6;
60478	:douta	=	16'h	82c6;
60479	:douta	=	16'h	82c6;
60480	:douta	=	16'h	8ac6;
60481	:douta	=	16'h	8ae7;
60482	:douta	=	16'h	8ae7;
60483	:douta	=	16'h	8ae7;
60484	:douta	=	16'h	9307;
60485	:douta	=	16'h	92e7;
60486	:douta	=	16'h	9307;
60487	:douta	=	16'h	9326;
60488	:douta	=	16'h	9b27;
60489	:douta	=	16'h	9b27;
60490	:douta	=	16'h	92c5;
60491	:douta	=	16'h	bc8e;
60492	:douta	=	16'h	c5d4;
60493	:douta	=	16'h	18c3;
60494	:douta	=	16'h	41e6;
60495	:douta	=	16'h	8aea;
60496	:douta	=	16'h	f739;
60497	:douta	=	16'h	59e5;
60498	:douta	=	16'h	a325;
60499	:douta	=	16'h	b3c8;
60500	:douta	=	16'h	b3c7;
60501	:douta	=	16'h	b3c7;
60502	:douta	=	16'h	bc08;
60503	:douta	=	16'h	bc08;
60504	:douta	=	16'h	bc08;
60505	:douta	=	16'h	bc07;
60506	:douta	=	16'h	bc07;
60507	:douta	=	16'h	bc07;
60508	:douta	=	16'h	bc08;
60509	:douta	=	16'h	bc08;
60510	:douta	=	16'h	c428;
60511	:douta	=	16'h	c428;
60512	:douta	=	16'h	c428;
60513	:douta	=	16'h	c428;
60514	:douta	=	16'h	c428;
60515	:douta	=	16'h	c448;
60516	:douta	=	16'h	c448;
60517	:douta	=	16'h	c448;
60518	:douta	=	16'h	c448;
60519	:douta	=	16'h	c448;
60520	:douta	=	16'h	c428;
60521	:douta	=	16'h	c448;
60522	:douta	=	16'h	c448;
60523	:douta	=	16'h	c448;
60524	:douta	=	16'h	c448;
60525	:douta	=	16'h	cc49;
60526	:douta	=	16'h	cc68;
60527	:douta	=	16'h	cc68;
60528	:douta	=	16'h	c448;
60529	:douta	=	16'h	cc68;
60530	:douta	=	16'h	cc68;
60531	:douta	=	16'h	cc68;
60532	:douta	=	16'h	cc68;
60533	:douta	=	16'h	cc68;
60534	:douta	=	16'h	cc68;
60535	:douta	=	16'h	cc68;
60536	:douta	=	16'h	cc69;
60537	:douta	=	16'h	cc68;
60538	:douta	=	16'h	cc69;
60539	:douta	=	16'h	cc69;
60540	:douta	=	16'h	cc68;
60541	:douta	=	16'h	cc69;
60542	:douta	=	16'h	cc69;
60543	:douta	=	16'h	cc69;
60544	:douta	=	16'h	cc69;
60545	:douta	=	16'h	cc69;
60546	:douta	=	16'h	cc69;
60547	:douta	=	16'h	cc69;
60548	:douta	=	16'h	cc69;
60549	:douta	=	16'h	cc89;
60550	:douta	=	16'h	cc89;
60551	:douta	=	16'h	cc69;
60552	:douta	=	16'h	cc89;
60553	:douta	=	16'h	cc89;
60554	:douta	=	16'h	cc89;
60555	:douta	=	16'h	cc89;
60556	:douta	=	16'h	cc89;
60557	:douta	=	16'h	cc89;
60558	:douta	=	16'h	cc89;
60559	:douta	=	16'h	cc89;
60560	:douta	=	16'h	cc89;
60561	:douta	=	16'h	cc89;
60562	:douta	=	16'h	cc89;
60563	:douta	=	16'h	cc89;
60564	:douta	=	16'h	cc89;
60565	:douta	=	16'h	cc89;
60566	:douta	=	16'h	cc89;
60567	:douta	=	16'h	cc89;
60568	:douta	=	16'h	cc89;
60569	:douta	=	16'h	cc69;
60570	:douta	=	16'h	cc89;
60571	:douta	=	16'h	cc69;
60572	:douta	=	16'h	cc69;
60573	:douta	=	16'h	cc89;
60574	:douta	=	16'h	cc89;
60575	:douta	=	16'h	cc89;
60576	:douta	=	16'h	cc69;
60577	:douta	=	16'h	cc89;
60578	:douta	=	16'h	cc88;
60579	:douta	=	16'h	b594;
60580	:douta	=	16'h	e696;
60581	:douta	=	16'h	cc48;
60582	:douta	=	16'h	cc69;
60583	:douta	=	16'h	cc89;
60584	:douta	=	16'h	cc68;
60585	:douta	=	16'h	cc69;
60586	:douta	=	16'h	cc89;
60587	:douta	=	16'h	cc69;
60588	:douta	=	16'h	cc69;
60589	:douta	=	16'h	cc69;
60590	:douta	=	16'h	cc69;
60591	:douta	=	16'h	cc69;
60592	:douta	=	16'h	cc69;
60593	:douta	=	16'h	cc69;
60594	:douta	=	16'h	cc6a;
60595	:douta	=	16'h	cc69;
60596	:douta	=	16'h	cc69;
60597	:douta	=	16'h	cc69;
60598	:douta	=	16'h	cc69;
60599	:douta	=	16'h	cc69;
60600	:douta	=	16'h	cc69;
60601	:douta	=	16'h	cc49;
60602	:douta	=	16'h	cc69;
60603	:douta	=	16'h	c449;
60604	:douta	=	16'h	cc49;
60605	:douta	=	16'h	cc69;
60606	:douta	=	16'h	cc6a;
60607	:douta	=	16'h	c449;
60608	:douta	=	16'h	c449;
60609	:douta	=	16'h	c449;
60610	:douta	=	16'h	c449;
60611	:douta	=	16'h	c449;
60612	:douta	=	16'h	c449;
60613	:douta	=	16'h	c449;
60614	:douta	=	16'h	c429;
60615	:douta	=	16'h	c449;
60616	:douta	=	16'h	c449;
60617	:douta	=	16'h	c429;
60618	:douta	=	16'h	c429;
60619	:douta	=	16'h	c429;
60620	:douta	=	16'h	c429;
60621	:douta	=	16'h	c429;
60622	:douta	=	16'h	c44a;
60623	:douta	=	16'h	c429;
60624	:douta	=	16'h	c429;
60625	:douta	=	16'h	c429;
60626	:douta	=	16'h	c429;
60627	:douta	=	16'h	c429;
60628	:douta	=	16'h	c429;
60629	:douta	=	16'h	bc09;
60630	:douta	=	16'h	bc09;
60631	:douta	=	16'h	bc09;
60632	:douta	=	16'h	bc09;
60633	:douta	=	16'h	bc09;
60634	:douta	=	16'h	bc09;
60635	:douta	=	16'h	bbe9;
60636	:douta	=	16'h	bc09;
60637	:douta	=	16'h	bc09;
60638	:douta	=	16'h	bc09;
60639	:douta	=	16'h	b3e9;
60640	:douta	=	16'h	b3e9;
60641	:douta	=	16'h	bbe9;
60642	:douta	=	16'h	bc09;
60643	:douta	=	16'h	b3e9;
60644	:douta	=	16'h	bbe9;
60645	:douta	=	16'h	bbe9;
60646	:douta	=	16'h	bbe9;
60647	:douta	=	16'h	b3e9;
60648	:douta	=	16'h	b3e9;
60649	:douta	=	16'h	b3e9;
60650	:douta	=	16'h	b3c9;
60651	:douta	=	16'h	b3c9;
60652	:douta	=	16'h	b3c9;
60653	:douta	=	16'h	aba9;
60654	:douta	=	16'h	b3ea;
60655	:douta	=	16'h	b3ca;
60656	:douta	=	16'h	b3ca;
60657	:douta	=	16'h	abc9;
60658	:douta	=	16'h	aba9;
60659	:douta	=	16'h	aba9;
60660	:douta	=	16'h	aba9;
60661	:douta	=	16'h	aba9;
60662	:douta	=	16'h	aba9;
60663	:douta	=	16'h	abc9;
60664	:douta	=	16'h	aba9;
60665	:douta	=	16'h	aba9;
60666	:douta	=	16'h	a388;
60667	:douta	=	16'h	aba8;
60668	:douta	=	16'h	a389;
60669	:douta	=	16'h	a389;
60670	:douta	=	16'h	a389;
60671	:douta	=	16'h	a389;
60672	:douta	=	16'h	9495;
60673	:douta	=	16'h	8cb6;
60674	:douta	=	16'h	8496;
60675	:douta	=	16'h	528c;
60676	:douta	=	16'h	2924;
60677	:douta	=	16'h	2904;
60678	:douta	=	16'h	2904;
60679	:douta	=	16'h	2904;
60680	:douta	=	16'h	20e3;
60681	:douta	=	16'h	20e3;
60682	:douta	=	16'h	28e3;
60683	:douta	=	16'h	2904;
60684	:douta	=	16'h	2904;
60685	:douta	=	16'h	28e3;
60686	:douta	=	16'h	2904;
60687	:douta	=	16'h	2904;
60688	:douta	=	16'h	20e3;
60689	:douta	=	16'h	20e3;
60690	:douta	=	16'h	20e3;
60691	:douta	=	16'h	20e3;
60692	:douta	=	16'h	1882;
60693	:douta	=	16'h	20a3;
60694	:douta	=	16'h	20c3;
60695	:douta	=	16'h	28e3;
60696	:douta	=	16'h	28e3;
60697	:douta	=	16'h	28e3;
60698	:douta	=	16'h	28c3;
60699	:douta	=	16'h	28e3;
60700	:douta	=	16'h	28e3;
60701	:douta	=	16'h	30e3;
60702	:douta	=	16'h	30e3;
60703	:douta	=	16'h	3103;
60704	:douta	=	16'h	3103;
60705	:douta	=	16'h	3123;
60706	:douta	=	16'h	3943;
60707	:douta	=	16'h	3943;
60708	:douta	=	16'h	4164;
60709	:douta	=	16'h	4144;
60710	:douta	=	16'h	4163;
60711	:douta	=	16'h	4964;
60712	:douta	=	16'h	49a5;
60713	:douta	=	16'h	4249;
60714	:douta	=	16'h	18e5;
60715	:douta	=	16'h	4984;
60716	:douta	=	16'h	59c4;
60717	:douta	=	16'h	59c4;
60718	:douta	=	16'h	61e4;
60719	:douta	=	16'h	61e4;
60720	:douta	=	16'h	6204;
60721	:douta	=	16'h	6a24;
60722	:douta	=	16'h	6a24;
60723	:douta	=	16'h	7245;
60724	:douta	=	16'h	7224;
60725	:douta	=	16'h	7224;
60726	:douta	=	16'h	b594;
60727	:douta	=	16'h	93eb;
60728	:douta	=	16'h	7a84;
60729	:douta	=	16'h	7a85;
60730	:douta	=	16'h	8285;
60731	:douta	=	16'h	8285;
60732	:douta	=	16'h	82c6;
60733	:douta	=	16'h	82c6;
60734	:douta	=	16'h	82c6;
60735	:douta	=	16'h	82c6;
60736	:douta	=	16'h	8ae7;
60737	:douta	=	16'h	8ae7;
60738	:douta	=	16'h	8b07;
60739	:douta	=	16'h	8ae7;
60740	:douta	=	16'h	9307;
60741	:douta	=	16'h	9307;
60742	:douta	=	16'h	9307;
60743	:douta	=	16'h	9b27;
60744	:douta	=	16'h	9b27;
60745	:douta	=	16'h	9b27;
60746	:douta	=	16'h	92e5;
60747	:douta	=	16'h	cd52;
60748	:douta	=	16'h	7c0c;
60749	:douta	=	16'h	0000;
60750	:douta	=	16'h	20a3;
60751	:douta	=	16'h	cdb3;
60752	:douta	=	16'h	f75a;
60753	:douta	=	16'h	59a4;
60754	:douta	=	16'h	b3c7;
60755	:douta	=	16'h	aba7;
60756	:douta	=	16'h	b3c7;
60757	:douta	=	16'h	b3c7;
60758	:douta	=	16'h	b3e8;
60759	:douta	=	16'h	b3c7;
60760	:douta	=	16'h	bc08;
60761	:douta	=	16'h	bc08;
60762	:douta	=	16'h	bc07;
60763	:douta	=	16'h	bc08;
60764	:douta	=	16'h	bc08;
60765	:douta	=	16'h	bc08;
60766	:douta	=	16'h	bc07;
60767	:douta	=	16'h	c428;
60768	:douta	=	16'h	c428;
60769	:douta	=	16'h	c428;
60770	:douta	=	16'h	c448;
60771	:douta	=	16'h	c448;
60772	:douta	=	16'h	c449;
60773	:douta	=	16'h	cc49;
60774	:douta	=	16'h	cc49;
60775	:douta	=	16'h	c428;
60776	:douta	=	16'h	c448;
60777	:douta	=	16'h	c448;
60778	:douta	=	16'h	c449;
60779	:douta	=	16'h	c449;
60780	:douta	=	16'h	c448;
60781	:douta	=	16'h	c448;
60782	:douta	=	16'h	c448;
60783	:douta	=	16'h	c448;
60784	:douta	=	16'h	cc68;
60785	:douta	=	16'h	cc69;
60786	:douta	=	16'h	cc69;
60787	:douta	=	16'h	cc49;
60788	:douta	=	16'h	cc68;
60789	:douta	=	16'h	cc68;
60790	:douta	=	16'h	cc68;
60791	:douta	=	16'h	cc69;
60792	:douta	=	16'h	cc68;
60793	:douta	=	16'h	cc69;
60794	:douta	=	16'h	cc69;
60795	:douta	=	16'h	cc69;
60796	:douta	=	16'h	cc89;
60797	:douta	=	16'h	cc69;
60798	:douta	=	16'h	cc89;
60799	:douta	=	16'h	cc89;
60800	:douta	=	16'h	cc89;
60801	:douta	=	16'h	cc89;
60802	:douta	=	16'h	cc69;
60803	:douta	=	16'h	cc69;
60804	:douta	=	16'h	cc69;
60805	:douta	=	16'h	cc89;
60806	:douta	=	16'h	cc69;
60807	:douta	=	16'h	cc89;
60808	:douta	=	16'h	cc89;
60809	:douta	=	16'h	cc89;
60810	:douta	=	16'h	cc89;
60811	:douta	=	16'h	cc89;
60812	:douta	=	16'h	cc89;
60813	:douta	=	16'h	cc89;
60814	:douta	=	16'h	cc89;
60815	:douta	=	16'h	cc69;
60816	:douta	=	16'h	cc89;
60817	:douta	=	16'h	cc89;
60818	:douta	=	16'h	cc89;
60819	:douta	=	16'h	cc89;
60820	:douta	=	16'h	cc89;
60821	:douta	=	16'h	cc89;
60822	:douta	=	16'h	cc69;
60823	:douta	=	16'h	cc89;
60824	:douta	=	16'h	cc69;
60825	:douta	=	16'h	cc89;
60826	:douta	=	16'h	cc69;
60827	:douta	=	16'h	cc69;
60828	:douta	=	16'h	cc69;
60829	:douta	=	16'h	cc69;
60830	:douta	=	16'h	cc69;
60831	:douta	=	16'h	cc89;
60832	:douta	=	16'h	cc89;
60833	:douta	=	16'h	cc69;
60834	:douta	=	16'h	cc69;
60835	:douta	=	16'h	b5b5;
60836	:douta	=	16'h	e696;
60837	:douta	=	16'h	cc48;
60838	:douta	=	16'h	cc69;
60839	:douta	=	16'h	cc69;
60840	:douta	=	16'h	cc69;
60841	:douta	=	16'h	cc6a;
60842	:douta	=	16'h	cc69;
60843	:douta	=	16'h	cc69;
60844	:douta	=	16'h	cc69;
60845	:douta	=	16'h	cc69;
60846	:douta	=	16'h	cc69;
60847	:douta	=	16'h	cc69;
60848	:douta	=	16'h	cc6a;
60849	:douta	=	16'h	cc6a;
60850	:douta	=	16'h	cc69;
60851	:douta	=	16'h	cc69;
60852	:douta	=	16'h	cc69;
60853	:douta	=	16'h	cc69;
60854	:douta	=	16'h	cc69;
60855	:douta	=	16'h	cc49;
60856	:douta	=	16'h	cc49;
60857	:douta	=	16'h	c449;
60858	:douta	=	16'h	cc49;
60859	:douta	=	16'h	cc49;
60860	:douta	=	16'h	cc49;
60861	:douta	=	16'h	cc49;
60862	:douta	=	16'h	c449;
60863	:douta	=	16'h	c449;
60864	:douta	=	16'h	cc6a;
60865	:douta	=	16'h	c429;
60866	:douta	=	16'h	c44a;
60867	:douta	=	16'h	c449;
60868	:douta	=	16'h	c44a;
60869	:douta	=	16'h	c429;
60870	:douta	=	16'h	c44a;
60871	:douta	=	16'h	c429;
60872	:douta	=	16'h	c429;
60873	:douta	=	16'h	c429;
60874	:douta	=	16'h	c449;
60875	:douta	=	16'h	bc29;
60876	:douta	=	16'h	c429;
60877	:douta	=	16'h	c429;
60878	:douta	=	16'h	c429;
60879	:douta	=	16'h	c429;
60880	:douta	=	16'h	c429;
60881	:douta	=	16'h	c429;
60882	:douta	=	16'h	bc09;
60883	:douta	=	16'h	bc29;
60884	:douta	=	16'h	bc09;
60885	:douta	=	16'h	bc09;
60886	:douta	=	16'h	c40a;
60887	:douta	=	16'h	bc2a;
60888	:douta	=	16'h	bc2a;
60889	:douta	=	16'h	bc09;
60890	:douta	=	16'h	bc09;
60891	:douta	=	16'h	bc09;
60892	:douta	=	16'h	bc09;
60893	:douta	=	16'h	bc09;
60894	:douta	=	16'h	bbe9;
60895	:douta	=	16'h	bc09;
60896	:douta	=	16'h	bc09;
60897	:douta	=	16'h	bbe9;
60898	:douta	=	16'h	b3e9;
60899	:douta	=	16'h	bc09;
60900	:douta	=	16'h	bbe9;
60901	:douta	=	16'h	b3c9;
60902	:douta	=	16'h	bbe9;
60903	:douta	=	16'h	bbe9;
60904	:douta	=	16'h	b3e9;
60905	:douta	=	16'h	b3e9;
60906	:douta	=	16'h	b3e9;
60907	:douta	=	16'h	b3e9;
60908	:douta	=	16'h	b3c9;
60909	:douta	=	16'h	abc9;
60910	:douta	=	16'h	b3ca;
60911	:douta	=	16'h	b3c9;
60912	:douta	=	16'h	aba9;
60913	:douta	=	16'h	aba9;
60914	:douta	=	16'h	b3c9;
60915	:douta	=	16'h	abc9;
60916	:douta	=	16'h	aba9;
60917	:douta	=	16'h	aba9;
60918	:douta	=	16'h	abc9;
60919	:douta	=	16'h	aba8;
60920	:douta	=	16'h	aba9;
60921	:douta	=	16'h	ab89;
60922	:douta	=	16'h	aba9;
60923	:douta	=	16'h	a388;
60924	:douta	=	16'h	ab89;
60925	:douta	=	16'h	a389;
60926	:douta	=	16'h	a389;
60927	:douta	=	16'h	a389;
60928	:douta	=	16'h	9495;
60929	:douta	=	16'h	8495;
60930	:douta	=	16'h	84b7;
60931	:douta	=	16'h	3166;
60932	:douta	=	16'h	2904;
60933	:douta	=	16'h	2904;
60934	:douta	=	16'h	2904;
60935	:douta	=	16'h	28e3;
60936	:douta	=	16'h	28e3;
60937	:douta	=	16'h	20e3;
60938	:douta	=	16'h	28e3;
60939	:douta	=	16'h	2904;
60940	:douta	=	16'h	2904;
60941	:douta	=	16'h	20e3;
60942	:douta	=	16'h	20e4;
60943	:douta	=	16'h	20e3;
60944	:douta	=	16'h	2904;
60945	:douta	=	16'h	20e3;
60946	:douta	=	16'h	20e3;
60947	:douta	=	16'h	20a2;
60948	:douta	=	16'h	20a2;
60949	:douta	=	16'h	20c3;
60950	:douta	=	16'h	20c3;
60951	:douta	=	16'h	20c2;
60952	:douta	=	16'h	28e2;
60953	:douta	=	16'h	28e3;
60954	:douta	=	16'h	28e3;
60955	:douta	=	16'h	28e3;
60956	:douta	=	16'h	28e3;
60957	:douta	=	16'h	3103;
60958	:douta	=	16'h	3103;
60959	:douta	=	16'h	3103;
60960	:douta	=	16'h	3103;
60961	:douta	=	16'h	3923;
60962	:douta	=	16'h	3944;
60963	:douta	=	16'h	3923;
60964	:douta	=	16'h	4144;
60965	:douta	=	16'h	4164;
60966	:douta	=	16'h	4163;
60967	:douta	=	16'h	4943;
60968	:douta	=	16'h	49c6;
60969	:douta	=	16'h	3a09;
60970	:douta	=	16'h	10c4;
60971	:douta	=	16'h	51a5;
60972	:douta	=	16'h	59c4;
60973	:douta	=	16'h	59c4;
60974	:douta	=	16'h	6205;
60975	:douta	=	16'h	6204;
60976	:douta	=	16'h	6205;
60977	:douta	=	16'h	6a24;
60978	:douta	=	16'h	6a44;
60979	:douta	=	16'h	7245;
60980	:douta	=	16'h	7244;
60981	:douta	=	16'h	7246;
60982	:douta	=	16'h	b572;
60983	:douta	=	16'h	8b49;
60984	:douta	=	16'h	7a85;
60985	:douta	=	16'h	82a5;
60986	:douta	=	16'h	7a85;
60987	:douta	=	16'h	82a5;
60988	:douta	=	16'h	82c6;
60989	:douta	=	16'h	82c6;
60990	:douta	=	16'h	82c6;
60991	:douta	=	16'h	8ac6;
60992	:douta	=	16'h	8ae7;
60993	:douta	=	16'h	8b07;
60994	:douta	=	16'h	8b07;
60995	:douta	=	16'h	9307;
60996	:douta	=	16'h	9307;
60997	:douta	=	16'h	8b07;
60998	:douta	=	16'h	9307;
60999	:douta	=	16'h	9b27;
61000	:douta	=	16'h	9b47;
61001	:douta	=	16'h	9b47;
61002	:douta	=	16'h	9b26;
61003	:douta	=	16'h	d5b3;
61004	:douta	=	16'h	bdd3;
61005	:douta	=	16'h	10e2;
61006	:douta	=	16'h	1861;
61007	:douta	=	16'h	e6d8;
61008	:douta	=	16'h	eed8;
61009	:douta	=	16'h	61c3;
61010	:douta	=	16'h	bbe8;
61011	:douta	=	16'h	abc7;
61012	:douta	=	16'h	b3c7;
61013	:douta	=	16'h	b3e8;
61014	:douta	=	16'h	b3c8;
61015	:douta	=	16'h	b3e7;
61016	:douta	=	16'h	bbe8;
61017	:douta	=	16'h	bc08;
61018	:douta	=	16'h	bbe8;
61019	:douta	=	16'h	bc08;
61020	:douta	=	16'h	bc08;
61021	:douta	=	16'h	bc08;
61022	:douta	=	16'h	c428;
61023	:douta	=	16'h	c408;
61024	:douta	=	16'h	c428;
61025	:douta	=	16'h	c428;
61026	:douta	=	16'h	c448;
61027	:douta	=	16'h	c428;
61028	:douta	=	16'h	c449;
61029	:douta	=	16'h	c448;
61030	:douta	=	16'h	c448;
61031	:douta	=	16'h	c448;
61032	:douta	=	16'h	c448;
61033	:douta	=	16'h	c449;
61034	:douta	=	16'h	c449;
61035	:douta	=	16'h	c448;
61036	:douta	=	16'h	cc49;
61037	:douta	=	16'h	cc49;
61038	:douta	=	16'h	c449;
61039	:douta	=	16'h	cc69;
61040	:douta	=	16'h	cc69;
61041	:douta	=	16'h	c449;
61042	:douta	=	16'h	cc69;
61043	:douta	=	16'h	cc69;
61044	:douta	=	16'h	cc68;
61045	:douta	=	16'h	cc68;
61046	:douta	=	16'h	cc69;
61047	:douta	=	16'h	cc68;
61048	:douta	=	16'h	cc68;
61049	:douta	=	16'h	cc69;
61050	:douta	=	16'h	cc69;
61051	:douta	=	16'h	cc69;
61052	:douta	=	16'h	cc69;
61053	:douta	=	16'h	cc69;
61054	:douta	=	16'h	cc69;
61055	:douta	=	16'h	cc89;
61056	:douta	=	16'h	cc69;
61057	:douta	=	16'h	cc89;
61058	:douta	=	16'h	cc69;
61059	:douta	=	16'h	cc89;
61060	:douta	=	16'h	cc69;
61061	:douta	=	16'h	cc69;
61062	:douta	=	16'h	cc89;
61063	:douta	=	16'h	cc89;
61064	:douta	=	16'h	cc89;
61065	:douta	=	16'h	cc89;
61066	:douta	=	16'h	cc89;
61067	:douta	=	16'h	cc89;
61068	:douta	=	16'h	cc89;
61069	:douta	=	16'h	cc89;
61070	:douta	=	16'h	cc89;
61071	:douta	=	16'h	cc89;
61072	:douta	=	16'h	cc8a;
61073	:douta	=	16'h	cc89;
61074	:douta	=	16'h	cc89;
61075	:douta	=	16'h	cc69;
61076	:douta	=	16'h	cc69;
61077	:douta	=	16'h	cc69;
61078	:douta	=	16'h	cc69;
61079	:douta	=	16'h	cc89;
61080	:douta	=	16'h	cc89;
61081	:douta	=	16'h	cc69;
61082	:douta	=	16'h	cc69;
61083	:douta	=	16'h	cc69;
61084	:douta	=	16'h	cc89;
61085	:douta	=	16'h	cc89;
61086	:douta	=	16'h	cc69;
61087	:douta	=	16'h	cc89;
61088	:douta	=	16'h	cc69;
61089	:douta	=	16'h	cc89;
61090	:douta	=	16'h	cc69;
61091	:douta	=	16'h	b5b5;
61092	:douta	=	16'h	e696;
61093	:douta	=	16'h	cc49;
61094	:douta	=	16'h	cc6a;
61095	:douta	=	16'h	cc69;
61096	:douta	=	16'h	cc49;
61097	:douta	=	16'h	cc69;
61098	:douta	=	16'h	cc89;
61099	:douta	=	16'h	cc69;
61100	:douta	=	16'h	cc69;
61101	:douta	=	16'h	cc69;
61102	:douta	=	16'h	cc69;
61103	:douta	=	16'h	cc69;
61104	:douta	=	16'h	cc69;
61105	:douta	=	16'h	cc6a;
61106	:douta	=	16'h	cc69;
61107	:douta	=	16'h	cc69;
61108	:douta	=	16'h	cc49;
61109	:douta	=	16'h	cc49;
61110	:douta	=	16'h	cc69;
61111	:douta	=	16'h	cc49;
61112	:douta	=	16'h	cc69;
61113	:douta	=	16'h	cc69;
61114	:douta	=	16'h	cc69;
61115	:douta	=	16'h	c449;
61116	:douta	=	16'h	c449;
61117	:douta	=	16'h	c449;
61118	:douta	=	16'h	c449;
61119	:douta	=	16'h	cc49;
61120	:douta	=	16'h	c449;
61121	:douta	=	16'h	c449;
61122	:douta	=	16'h	c449;
61123	:douta	=	16'h	c429;
61124	:douta	=	16'h	c449;
61125	:douta	=	16'h	c44a;
61126	:douta	=	16'h	c449;
61127	:douta	=	16'h	c429;
61128	:douta	=	16'h	c429;
61129	:douta	=	16'h	c429;
61130	:douta	=	16'h	c429;
61131	:douta	=	16'h	c429;
61132	:douta	=	16'h	c429;
61133	:douta	=	16'h	c429;
61134	:douta	=	16'h	c429;
61135	:douta	=	16'h	c44a;
61136	:douta	=	16'h	bc09;
61137	:douta	=	16'h	c429;
61138	:douta	=	16'h	bc09;
61139	:douta	=	16'h	c429;
61140	:douta	=	16'h	c40a;
61141	:douta	=	16'h	bc2a;
61142	:douta	=	16'h	bc09;
61143	:douta	=	16'h	bc09;
61144	:douta	=	16'h	bc09;
61145	:douta	=	16'h	bc09;
61146	:douta	=	16'h	bc09;
61147	:douta	=	16'h	bc09;
61148	:douta	=	16'h	bc09;
61149	:douta	=	16'h	bc09;
61150	:douta	=	16'h	bc09;
61151	:douta	=	16'h	bc09;
61152	:douta	=	16'h	bbe9;
61153	:douta	=	16'h	b3e9;
61154	:douta	=	16'h	bbe9;
61155	:douta	=	16'h	bbe9;
61156	:douta	=	16'h	bc09;
61157	:douta	=	16'h	bbe9;
61158	:douta	=	16'h	bbe9;
61159	:douta	=	16'h	bbe9;
61160	:douta	=	16'h	b3e9;
61161	:douta	=	16'h	b3c9;
61162	:douta	=	16'h	b3e9;
61163	:douta	=	16'h	b3ca;
61164	:douta	=	16'h	b3ca;
61165	:douta	=	16'h	b3ca;
61166	:douta	=	16'h	b3c9;
61167	:douta	=	16'h	b3c9;
61168	:douta	=	16'h	abc9;
61169	:douta	=	16'h	abc9;
61170	:douta	=	16'h	abc9;
61171	:douta	=	16'h	aba9;
61172	:douta	=	16'h	aba9;
61173	:douta	=	16'h	abc9;
61174	:douta	=	16'h	abc9;
61175	:douta	=	16'h	aba9;
61176	:douta	=	16'h	aba8;
61177	:douta	=	16'h	aba9;
61178	:douta	=	16'h	aba9;
61179	:douta	=	16'h	a389;
61180	:douta	=	16'h	a389;
61181	:douta	=	16'h	aba9;
61182	:douta	=	16'h	a389;
61183	:douta	=	16'h	a389;
61184	:douta	=	16'h	8c95;
61185	:douta	=	16'h	84b7;
61186	:douta	=	16'h	9d5a;
61187	:douta	=	16'h	1861;
61188	:douta	=	16'h	2904;
61189	:douta	=	16'h	2904;
61190	:douta	=	16'h	2904;
61191	:douta	=	16'h	20e3;
61192	:douta	=	16'h	2904;
61193	:douta	=	16'h	28e3;
61194	:douta	=	16'h	28e3;
61195	:douta	=	16'h	2904;
61196	:douta	=	16'h	2904;
61197	:douta	=	16'h	2904;
61198	:douta	=	16'h	20e3;
61199	:douta	=	16'h	20e3;
61200	:douta	=	16'h	20e3;
61201	:douta	=	16'h	20e3;
61202	:douta	=	16'h	28e3;
61203	:douta	=	16'h	20a3;
61204	:douta	=	16'h	20a3;
61205	:douta	=	16'h	20c2;
61206	:douta	=	16'h	20c2;
61207	:douta	=	16'h	20c2;
61208	:douta	=	16'h	28e3;
61209	:douta	=	16'h	28e3;
61210	:douta	=	16'h	28e3;
61211	:douta	=	16'h	28e3;
61212	:douta	=	16'h	28e3;
61213	:douta	=	16'h	30e3;
61214	:douta	=	16'h	3103;
61215	:douta	=	16'h	3103;
61216	:douta	=	16'h	3103;
61217	:douta	=	16'h	3923;
61218	:douta	=	16'h	3923;
61219	:douta	=	16'h	3944;
61220	:douta	=	16'h	4164;
61221	:douta	=	16'h	4164;
61222	:douta	=	16'h	4164;
61223	:douta	=	16'h	4964;
61224	:douta	=	16'h	4a28;
61225	:douta	=	16'h	2947;
61226	:douta	=	16'h	0885;
61227	:douta	=	16'h	6204;
61228	:douta	=	16'h	59c4;
61229	:douta	=	16'h	59c4;
61230	:douta	=	16'h	59e4;
61231	:douta	=	16'h	6204;
61232	:douta	=	16'h	6204;
61233	:douta	=	16'h	6a25;
61234	:douta	=	16'h	6a24;
61235	:douta	=	16'h	6a44;
61236	:douta	=	16'h	6a44;
61237	:douta	=	16'h	7288;
61238	:douta	=	16'h	ad10;
61239	:douta	=	16'h	7a85;
61240	:douta	=	16'h	7a85;
61241	:douta	=	16'h	7a85;
61242	:douta	=	16'h	8286;
61243	:douta	=	16'h	82a5;
61244	:douta	=	16'h	82a6;
61245	:douta	=	16'h	82c6;
61246	:douta	=	16'h	82c6;
61247	:douta	=	16'h	82c6;
61248	:douta	=	16'h	8ac6;
61249	:douta	=	16'h	8ae7;
61250	:douta	=	16'h	8ae7;
61251	:douta	=	16'h	8b07;
61252	:douta	=	16'h	9307;
61253	:douta	=	16'h	8b07;
61254	:douta	=	16'h	9327;
61255	:douta	=	16'h	9b47;
61256	:douta	=	16'h	9b47;
61257	:douta	=	16'h	9b27;
61258	:douta	=	16'h	b3eb;
61259	:douta	=	16'h	de77;
61260	:douta	=	16'h	d636;
61261	:douta	=	16'h	e6b7;
61262	:douta	=	16'h	e6b7;
61263	:douta	=	16'h	de76;
61264	:douta	=	16'h	de98;
61265	:douta	=	16'h	7a23;
61266	:douta	=	16'h	b3e8;
61267	:douta	=	16'h	abc8;
61268	:douta	=	16'h	b3c7;
61269	:douta	=	16'h	b3c7;
61270	:douta	=	16'h	b3e8;
61271	:douta	=	16'h	b3e8;
61272	:douta	=	16'h	bbe8;
61273	:douta	=	16'h	bc08;
61274	:douta	=	16'h	bc08;
61275	:douta	=	16'h	bc08;
61276	:douta	=	16'h	bc08;
61277	:douta	=	16'h	c408;
61278	:douta	=	16'h	bc08;
61279	:douta	=	16'h	c428;
61280	:douta	=	16'h	c428;
61281	:douta	=	16'h	c448;
61282	:douta	=	16'h	c448;
61283	:douta	=	16'h	c448;
61284	:douta	=	16'h	c449;
61285	:douta	=	16'h	c428;
61286	:douta	=	16'h	c448;
61287	:douta	=	16'h	c448;
61288	:douta	=	16'h	c448;
61289	:douta	=	16'h	c448;
61290	:douta	=	16'h	c448;
61291	:douta	=	16'h	c448;
61292	:douta	=	16'h	c449;
61293	:douta	=	16'h	c449;
61294	:douta	=	16'h	c468;
61295	:douta	=	16'h	c448;
61296	:douta	=	16'h	cc69;
61297	:douta	=	16'h	cc49;
61298	:douta	=	16'h	cc49;
61299	:douta	=	16'h	cc69;
61300	:douta	=	16'h	cc69;
61301	:douta	=	16'h	cc69;
61302	:douta	=	16'h	cc68;
61303	:douta	=	16'h	cc68;
61304	:douta	=	16'h	cc68;
61305	:douta	=	16'h	cc69;
61306	:douta	=	16'h	cc68;
61307	:douta	=	16'h	cc89;
61308	:douta	=	16'h	cc69;
61309	:douta	=	16'h	cc69;
61310	:douta	=	16'h	cc89;
61311	:douta	=	16'h	cc69;
61312	:douta	=	16'h	cc69;
61313	:douta	=	16'h	cc69;
61314	:douta	=	16'h	cc69;
61315	:douta	=	16'h	cc69;
61316	:douta	=	16'h	cc89;
61317	:douta	=	16'h	cc89;
61318	:douta	=	16'h	cc69;
61319	:douta	=	16'h	cc69;
61320	:douta	=	16'h	cc89;
61321	:douta	=	16'h	cc89;
61322	:douta	=	16'h	cc69;
61323	:douta	=	16'h	cc69;
61324	:douta	=	16'h	cc8a;
61325	:douta	=	16'h	cc89;
61326	:douta	=	16'h	cc89;
61327	:douta	=	16'h	cc89;
61328	:douta	=	16'h	cc89;
61329	:douta	=	16'h	cc89;
61330	:douta	=	16'h	cc89;
61331	:douta	=	16'h	cc89;
61332	:douta	=	16'h	cc89;
61333	:douta	=	16'h	cc69;
61334	:douta	=	16'h	cc89;
61335	:douta	=	16'h	cc89;
61336	:douta	=	16'h	cc69;
61337	:douta	=	16'h	cc89;
61338	:douta	=	16'h	cc89;
61339	:douta	=	16'h	cc69;
61340	:douta	=	16'h	cc69;
61341	:douta	=	16'h	cc69;
61342	:douta	=	16'h	cc69;
61343	:douta	=	16'h	cc89;
61344	:douta	=	16'h	cc89;
61345	:douta	=	16'h	cc89;
61346	:douta	=	16'h	cc89;
61347	:douta	=	16'h	b595;
61348	:douta	=	16'h	e675;
61349	:douta	=	16'h	cc49;
61350	:douta	=	16'h	cc69;
61351	:douta	=	16'h	cc6a;
61352	:douta	=	16'h	cc69;
61353	:douta	=	16'h	cc69;
61354	:douta	=	16'h	cc69;
61355	:douta	=	16'h	cc6a;
61356	:douta	=	16'h	cc6a;
61357	:douta	=	16'h	cc6a;
61358	:douta	=	16'h	cc6a;
61359	:douta	=	16'h	cc69;
61360	:douta	=	16'h	cc69;
61361	:douta	=	16'h	cc69;
61362	:douta	=	16'h	cc6a;
61363	:douta	=	16'h	cc49;
61364	:douta	=	16'h	cc69;
61365	:douta	=	16'h	cc69;
61366	:douta	=	16'h	cc49;
61367	:douta	=	16'h	c449;
61368	:douta	=	16'h	cc49;
61369	:douta	=	16'h	cc69;
61370	:douta	=	16'h	cc49;
61371	:douta	=	16'h	cc49;
61372	:douta	=	16'h	c449;
61373	:douta	=	16'h	c449;
61374	:douta	=	16'h	cc49;
61375	:douta	=	16'h	c449;
61376	:douta	=	16'h	c449;
61377	:douta	=	16'h	c469;
61378	:douta	=	16'h	c449;
61379	:douta	=	16'h	c449;
61380	:douta	=	16'h	c469;
61381	:douta	=	16'h	c449;
61382	:douta	=	16'h	c449;
61383	:douta	=	16'h	c449;
61384	:douta	=	16'h	c44a;
61385	:douta	=	16'h	c44a;
61386	:douta	=	16'h	c429;
61387	:douta	=	16'h	c429;
61388	:douta	=	16'h	c44a;
61389	:douta	=	16'h	bc29;
61390	:douta	=	16'h	bc29;
61391	:douta	=	16'h	c429;
61392	:douta	=	16'h	c429;
61393	:douta	=	16'h	c429;
61394	:douta	=	16'h	c42a;
61395	:douta	=	16'h	c40a;
61396	:douta	=	16'h	bc09;
61397	:douta	=	16'h	bc2a;
61398	:douta	=	16'h	bc2a;
61399	:douta	=	16'h	bc2a;
61400	:douta	=	16'h	bc09;
61401	:douta	=	16'h	bc09;
61402	:douta	=	16'h	bc09;
61403	:douta	=	16'h	bc09;
61404	:douta	=	16'h	bc09;
61405	:douta	=	16'h	bc09;
61406	:douta	=	16'h	bc09;
61407	:douta	=	16'h	bc09;
61408	:douta	=	16'h	bc09;
61409	:douta	=	16'h	bbe9;
61410	:douta	=	16'h	bc09;
61411	:douta	=	16'h	b3e9;
61412	:douta	=	16'h	b3e9;
61413	:douta	=	16'h	b3e9;
61414	:douta	=	16'h	b3e9;
61415	:douta	=	16'h	b3e9;
61416	:douta	=	16'h	b3e9;
61417	:douta	=	16'h	b3e9;
61418	:douta	=	16'h	b3e9;
61419	:douta	=	16'h	b3c9;
61420	:douta	=	16'h	b3e9;
61421	:douta	=	16'h	b3c9;
61422	:douta	=	16'h	b3ca;
61423	:douta	=	16'h	abc9;
61424	:douta	=	16'h	abc9;
61425	:douta	=	16'h	abc9;
61426	:douta	=	16'h	b3ca;
61427	:douta	=	16'h	abc9;
61428	:douta	=	16'h	abc9;
61429	:douta	=	16'h	aba9;
61430	:douta	=	16'h	aba9;
61431	:douta	=	16'h	abc9;
61432	:douta	=	16'h	aba9;
61433	:douta	=	16'h	aba9;
61434	:douta	=	16'h	aba9;
61435	:douta	=	16'h	aba9;
61436	:douta	=	16'h	aba9;
61437	:douta	=	16'h	a389;
61438	:douta	=	16'h	a389;
61439	:douta	=	16'h	a389;
61440	:douta	=	16'h	8c96;
61441	:douta	=	16'h	8cd8;
61442	:douta	=	16'h	84b7;
61443	:douta	=	16'h	20a2;
61444	:douta	=	16'h	2904;
61445	:douta	=	16'h	2904;
61446	:douta	=	16'h	2904;
61447	:douta	=	16'h	28e3;
61448	:douta	=	16'h	28e3;
61449	:douta	=	16'h	2904;
61450	:douta	=	16'h	2904;
61451	:douta	=	16'h	2904;
61452	:douta	=	16'h	2904;
61453	:douta	=	16'h	28e3;
61454	:douta	=	16'h	20e4;
61455	:douta	=	16'h	20e3;
61456	:douta	=	16'h	20e3;
61457	:douta	=	16'h	20e3;
61458	:douta	=	16'h	2904;
61459	:douta	=	16'h	20a2;
61460	:douta	=	16'h	20a3;
61461	:douta	=	16'h	20c2;
61462	:douta	=	16'h	20c2;
61463	:douta	=	16'h	20c2;
61464	:douta	=	16'h	28c3;
61465	:douta	=	16'h	28e3;
61466	:douta	=	16'h	28e3;
61467	:douta	=	16'h	28e3;
61468	:douta	=	16'h	28e3;
61469	:douta	=	16'h	30e3;
61470	:douta	=	16'h	3103;
61471	:douta	=	16'h	3103;
61472	:douta	=	16'h	3903;
61473	:douta	=	16'h	3123;
61474	:douta	=	16'h	3944;
61475	:douta	=	16'h	3944;
61476	:douta	=	16'h	4164;
61477	:douta	=	16'h	4164;
61478	:douta	=	16'h	4964;
61479	:douta	=	16'h	4985;
61480	:douta	=	16'h	4a29;
61481	:douta	=	16'h	2127;
61482	:douta	=	16'h	0885;
61483	:douta	=	16'h	61c4;
61484	:douta	=	16'h	59e4;
61485	:douta	=	16'h	59c4;
61486	:douta	=	16'h	61e4;
61487	:douta	=	16'h	6204;
61488	:douta	=	16'h	6205;
61489	:douta	=	16'h	6a25;
61490	:douta	=	16'h	6a44;
61491	:douta	=	16'h	6a44;
61492	:douta	=	16'h	7245;
61493	:douta	=	16'h	6aa8;
61494	:douta	=	16'h	accf;
61495	:douta	=	16'h	7244;
61496	:douta	=	16'h	7a85;
61497	:douta	=	16'h	8285;
61498	:douta	=	16'h	7a85;
61499	:douta	=	16'h	82a5;
61500	:douta	=	16'h	82c6;
61501	:douta	=	16'h	82c6;
61502	:douta	=	16'h	82c6;
61503	:douta	=	16'h	82c6;
61504	:douta	=	16'h	8ae7;
61505	:douta	=	16'h	8ac6;
61506	:douta	=	16'h	8ae7;
61507	:douta	=	16'h	8b07;
61508	:douta	=	16'h	8b07;
61509	:douta	=	16'h	9327;
61510	:douta	=	16'h	9327;
61511	:douta	=	16'h	9b47;
61512	:douta	=	16'h	9b47;
61513	:douta	=	16'h	9b27;
61514	:douta	=	16'h	c48f;
61515	:douta	=	16'h	eef9;
61516	:douta	=	16'h	deb8;
61517	:douta	=	16'h	deb8;
61518	:douta	=	16'h	e6d9;
61519	:douta	=	16'h	ef3b;
61520	:douta	=	16'h	ce78;
61521	:douta	=	16'h	92c3;
61522	:douta	=	16'h	b3e8;
61523	:douta	=	16'h	b3c8;
61524	:douta	=	16'h	b3c7;
61525	:douta	=	16'h	b3c8;
61526	:douta	=	16'h	b3e8;
61527	:douta	=	16'h	b3e8;
61528	:douta	=	16'h	bc08;
61529	:douta	=	16'h	bc08;
61530	:douta	=	16'h	bc08;
61531	:douta	=	16'h	bc08;
61532	:douta	=	16'h	bc08;
61533	:douta	=	16'h	c428;
61534	:douta	=	16'h	bc08;
61535	:douta	=	16'h	c428;
61536	:douta	=	16'h	c428;
61537	:douta	=	16'h	c448;
61538	:douta	=	16'h	c428;
61539	:douta	=	16'h	c428;
61540	:douta	=	16'h	c449;
61541	:douta	=	16'h	c449;
61542	:douta	=	16'h	c449;
61543	:douta	=	16'h	c448;
61544	:douta	=	16'h	c448;
61545	:douta	=	16'h	c448;
61546	:douta	=	16'h	c448;
61547	:douta	=	16'h	c448;
61548	:douta	=	16'h	c448;
61549	:douta	=	16'h	cc49;
61550	:douta	=	16'h	cc69;
61551	:douta	=	16'h	c468;
61552	:douta	=	16'h	cc69;
61553	:douta	=	16'h	cc69;
61554	:douta	=	16'h	cc49;
61555	:douta	=	16'h	cc69;
61556	:douta	=	16'h	cc69;
61557	:douta	=	16'h	cc69;
61558	:douta	=	16'h	cc69;
61559	:douta	=	16'h	cc69;
61560	:douta	=	16'h	cc69;
61561	:douta	=	16'h	cc69;
61562	:douta	=	16'h	cc69;
61563	:douta	=	16'h	cc89;
61564	:douta	=	16'h	cc69;
61565	:douta	=	16'h	cc89;
61566	:douta	=	16'h	cc89;
61567	:douta	=	16'h	cc89;
61568	:douta	=	16'h	cc69;
61569	:douta	=	16'h	cc89;
61570	:douta	=	16'h	cc89;
61571	:douta	=	16'h	cc69;
61572	:douta	=	16'h	cc69;
61573	:douta	=	16'h	cc89;
61574	:douta	=	16'h	cc69;
61575	:douta	=	16'h	cc89;
61576	:douta	=	16'h	cc69;
61577	:douta	=	16'h	cc69;
61578	:douta	=	16'h	cc89;
61579	:douta	=	16'h	cc69;
61580	:douta	=	16'h	cc89;
61581	:douta	=	16'h	cc89;
61582	:douta	=	16'h	cc89;
61583	:douta	=	16'h	cc89;
61584	:douta	=	16'h	cc69;
61585	:douta	=	16'h	cc89;
61586	:douta	=	16'h	cc89;
61587	:douta	=	16'h	cc89;
61588	:douta	=	16'h	cc89;
61589	:douta	=	16'h	cc69;
61590	:douta	=	16'h	cc89;
61591	:douta	=	16'h	cc69;
61592	:douta	=	16'h	cc69;
61593	:douta	=	16'h	cc89;
61594	:douta	=	16'h	cc89;
61595	:douta	=	16'h	cc69;
61596	:douta	=	16'h	cc89;
61597	:douta	=	16'h	cc89;
61598	:douta	=	16'h	cc89;
61599	:douta	=	16'h	cc89;
61600	:douta	=	16'h	cc89;
61601	:douta	=	16'h	cc69;
61602	:douta	=	16'h	cc69;
61603	:douta	=	16'h	b5b5;
61604	:douta	=	16'h	e675;
61605	:douta	=	16'h	cc49;
61606	:douta	=	16'h	cc6a;
61607	:douta	=	16'h	cc6a;
61608	:douta	=	16'h	cc69;
61609	:douta	=	16'h	cc69;
61610	:douta	=	16'h	cc69;
61611	:douta	=	16'h	cc6a;
61612	:douta	=	16'h	cc69;
61613	:douta	=	16'h	cc69;
61614	:douta	=	16'h	cc69;
61615	:douta	=	16'h	cc49;
61616	:douta	=	16'h	cc69;
61617	:douta	=	16'h	cc69;
61618	:douta	=	16'h	cc69;
61619	:douta	=	16'h	cc69;
61620	:douta	=	16'h	cc69;
61621	:douta	=	16'h	cc69;
61622	:douta	=	16'h	cc69;
61623	:douta	=	16'h	cc69;
61624	:douta	=	16'h	cc69;
61625	:douta	=	16'h	cc49;
61626	:douta	=	16'h	cc69;
61627	:douta	=	16'h	c449;
61628	:douta	=	16'h	cc69;
61629	:douta	=	16'h	c449;
61630	:douta	=	16'h	c449;
61631	:douta	=	16'h	c449;
61632	:douta	=	16'h	c449;
61633	:douta	=	16'h	c449;
61634	:douta	=	16'h	c449;
61635	:douta	=	16'h	c449;
61636	:douta	=	16'h	c449;
61637	:douta	=	16'h	c449;
61638	:douta	=	16'h	c469;
61639	:douta	=	16'h	c449;
61640	:douta	=	16'h	c44a;
61641	:douta	=	16'h	c429;
61642	:douta	=	16'h	c44a;
61643	:douta	=	16'h	c429;
61644	:douta	=	16'h	c429;
61645	:douta	=	16'h	c429;
61646	:douta	=	16'h	c429;
61647	:douta	=	16'h	c429;
61648	:douta	=	16'h	bc29;
61649	:douta	=	16'h	c40a;
61650	:douta	=	16'h	bc09;
61651	:douta	=	16'h	c40a;
61652	:douta	=	16'h	c40a;
61653	:douta	=	16'h	bc09;
61654	:douta	=	16'h	bc09;
61655	:douta	=	16'h	bc09;
61656	:douta	=	16'h	bc2a;
61657	:douta	=	16'h	bc09;
61658	:douta	=	16'h	bc09;
61659	:douta	=	16'h	bc09;
61660	:douta	=	16'h	bc09;
61661	:douta	=	16'h	bc09;
61662	:douta	=	16'h	bc09;
61663	:douta	=	16'h	bc09;
61664	:douta	=	16'h	bc09;
61665	:douta	=	16'h	bbe9;
61666	:douta	=	16'h	bc09;
61667	:douta	=	16'h	bbe9;
61668	:douta	=	16'h	bbe9;
61669	:douta	=	16'h	b3e9;
61670	:douta	=	16'h	bbe9;
61671	:douta	=	16'h	b3e9;
61672	:douta	=	16'h	bbe9;
61673	:douta	=	16'h	b3c9;
61674	:douta	=	16'h	b3e9;
61675	:douta	=	16'h	b3c9;
61676	:douta	=	16'h	b3e9;
61677	:douta	=	16'h	b3c9;
61678	:douta	=	16'h	b3ca;
61679	:douta	=	16'h	b3c9;
61680	:douta	=	16'h	abc9;
61681	:douta	=	16'h	b3c9;
61682	:douta	=	16'h	b3ca;
61683	:douta	=	16'h	abc9;
61684	:douta	=	16'h	abc9;
61685	:douta	=	16'h	aba9;
61686	:douta	=	16'h	aba9;
61687	:douta	=	16'h	aba9;
61688	:douta	=	16'h	aba9;
61689	:douta	=	16'h	aba9;
61690	:douta	=	16'h	ab89;
61691	:douta	=	16'h	aba9;
61692	:douta	=	16'h	a389;
61693	:douta	=	16'h	a389;
61694	:douta	=	16'h	a389;
61695	:douta	=	16'h	a369;
61696	:douta	=	16'h	8476;
61697	:douta	=	16'h	955a;
61698	:douta	=	16'h	52cc;
61699	:douta	=	16'h	2924;
61700	:douta	=	16'h	2904;
61701	:douta	=	16'h	2904;
61702	:douta	=	16'h	2904;
61703	:douta	=	16'h	2904;
61704	:douta	=	16'h	2904;
61705	:douta	=	16'h	2904;
61706	:douta	=	16'h	2904;
61707	:douta	=	16'h	2904;
61708	:douta	=	16'h	2904;
61709	:douta	=	16'h	28e3;
61710	:douta	=	16'h	20e3;
61711	:douta	=	16'h	20e3;
61712	:douta	=	16'h	20e3;
61713	:douta	=	16'h	20e3;
61714	:douta	=	16'h	2904;
61715	:douta	=	16'h	20a3;
61716	:douta	=	16'h	20c2;
61717	:douta	=	16'h	20c2;
61718	:douta	=	16'h	20c3;
61719	:douta	=	16'h	28c3;
61720	:douta	=	16'h	28e3;
61721	:douta	=	16'h	28e3;
61722	:douta	=	16'h	28e3;
61723	:douta	=	16'h	28e3;
61724	:douta	=	16'h	28e3;
61725	:douta	=	16'h	3103;
61726	:douta	=	16'h	3103;
61727	:douta	=	16'h	3103;
61728	:douta	=	16'h	3103;
61729	:douta	=	16'h	3923;
61730	:douta	=	16'h	3944;
61731	:douta	=	16'h	3944;
61732	:douta	=	16'h	4144;
61733	:douta	=	16'h	4164;
61734	:douta	=	16'h	4984;
61735	:douta	=	16'h	4985;
61736	:douta	=	16'h	528b;
61737	:douta	=	16'h	10e5;
61738	:douta	=	16'h	10a4;
61739	:douta	=	16'h	61e4;
61740	:douta	=	16'h	59c4;
61741	:douta	=	16'h	59c4;
61742	:douta	=	16'h	61e4;
61743	:douta	=	16'h	6204;
61744	:douta	=	16'h	6a25;
61745	:douta	=	16'h	6a44;
61746	:douta	=	16'h	6a45;
61747	:douta	=	16'h	7245;
61748	:douta	=	16'h	7245;
61749	:douta	=	16'h	736b;
61750	:douta	=	16'h	9c0b;
61751	:douta	=	16'h	7203;
61752	:douta	=	16'h	7a85;
61753	:douta	=	16'h	7a85;
61754	:douta	=	16'h	82a5;
61755	:douta	=	16'h	82c6;
61756	:douta	=	16'h	82c6;
61757	:douta	=	16'h	82c6;
61758	:douta	=	16'h	82c6;
61759	:douta	=	16'h	82c6;
61760	:douta	=	16'h	8ac6;
61761	:douta	=	16'h	8ae7;
61762	:douta	=	16'h	8b07;
61763	:douta	=	16'h	8ae7;
61764	:douta	=	16'h	9307;
61765	:douta	=	16'h	9307;
61766	:douta	=	16'h	9307;
61767	:douta	=	16'h	9b47;
61768	:douta	=	16'h	9b68;
61769	:douta	=	16'h	9b47;
61770	:douta	=	16'h	a388;
61771	:douta	=	16'h	a38b;
61772	:douta	=	16'h	9b48;
61773	:douta	=	16'h	9b48;
61774	:douta	=	16'h	9b07;
61775	:douta	=	16'h	9b05;
61776	:douta	=	16'h	a326;
61777	:douta	=	16'h	abc8;
61778	:douta	=	16'h	aba8;
61779	:douta	=	16'h	b3c7;
61780	:douta	=	16'h	b3c8;
61781	:douta	=	16'h	b3e8;
61782	:douta	=	16'h	b3e8;
61783	:douta	=	16'h	b3e8;
61784	:douta	=	16'h	b3e8;
61785	:douta	=	16'h	bc08;
61786	:douta	=	16'h	bc08;
61787	:douta	=	16'h	bc28;
61788	:douta	=	16'h	bc29;
61789	:douta	=	16'h	bc29;
61790	:douta	=	16'h	bc29;
61791	:douta	=	16'h	bc28;
61792	:douta	=	16'h	c448;
61793	:douta	=	16'h	c428;
61794	:douta	=	16'h	c449;
61795	:douta	=	16'h	c449;
61796	:douta	=	16'h	c449;
61797	:douta	=	16'h	c449;
61798	:douta	=	16'h	c449;
61799	:douta	=	16'h	c428;
61800	:douta	=	16'h	c448;
61801	:douta	=	16'h	c448;
61802	:douta	=	16'h	c448;
61803	:douta	=	16'h	c448;
61804	:douta	=	16'h	cc69;
61805	:douta	=	16'h	cc69;
61806	:douta	=	16'h	c448;
61807	:douta	=	16'h	cc69;
61808	:douta	=	16'h	cc69;
61809	:douta	=	16'h	cc69;
61810	:douta	=	16'h	cc69;
61811	:douta	=	16'h	cc69;
61812	:douta	=	16'h	cc69;
61813	:douta	=	16'h	cc69;
61814	:douta	=	16'h	cc69;
61815	:douta	=	16'h	cc69;
61816	:douta	=	16'h	cc69;
61817	:douta	=	16'h	cc69;
61818	:douta	=	16'h	cc69;
61819	:douta	=	16'h	cc69;
61820	:douta	=	16'h	cc89;
61821	:douta	=	16'h	cc69;
61822	:douta	=	16'h	cc69;
61823	:douta	=	16'h	cc89;
61824	:douta	=	16'h	cc89;
61825	:douta	=	16'h	cc89;
61826	:douta	=	16'h	cc69;
61827	:douta	=	16'h	cc69;
61828	:douta	=	16'h	cc89;
61829	:douta	=	16'h	cc69;
61830	:douta	=	16'h	cc89;
61831	:douta	=	16'h	cc89;
61832	:douta	=	16'h	cc69;
61833	:douta	=	16'h	cc89;
61834	:douta	=	16'h	cc89;
61835	:douta	=	16'h	cc89;
61836	:douta	=	16'h	cc89;
61837	:douta	=	16'h	cc89;
61838	:douta	=	16'h	cc89;
61839	:douta	=	16'h	cc89;
61840	:douta	=	16'h	cc89;
61841	:douta	=	16'h	cc69;
61842	:douta	=	16'h	cc69;
61843	:douta	=	16'h	cc69;
61844	:douta	=	16'h	cc69;
61845	:douta	=	16'h	cc69;
61846	:douta	=	16'h	cc69;
61847	:douta	=	16'h	cc69;
61848	:douta	=	16'h	cc89;
61849	:douta	=	16'h	cc69;
61850	:douta	=	16'h	cc69;
61851	:douta	=	16'h	cc89;
61852	:douta	=	16'h	cc89;
61853	:douta	=	16'h	cc89;
61854	:douta	=	16'h	cc89;
61855	:douta	=	16'h	c489;
61856	:douta	=	16'h	c489;
61857	:douta	=	16'h	cc89;
61858	:douta	=	16'h	cc68;
61859	:douta	=	16'h	b5b5;
61860	:douta	=	16'h	e655;
61861	:douta	=	16'h	cc69;
61862	:douta	=	16'h	cc6a;
61863	:douta	=	16'h	cc6a;
61864	:douta	=	16'h	cc89;
61865	:douta	=	16'h	cc89;
61866	:douta	=	16'h	cc69;
61867	:douta	=	16'h	cc69;
61868	:douta	=	16'h	cc6a;
61869	:douta	=	16'h	cc69;
61870	:douta	=	16'h	cc69;
61871	:douta	=	16'h	cc69;
61872	:douta	=	16'h	cc69;
61873	:douta	=	16'h	cc69;
61874	:douta	=	16'h	cc49;
61875	:douta	=	16'h	cc49;
61876	:douta	=	16'h	cc69;
61877	:douta	=	16'h	cc69;
61878	:douta	=	16'h	cc49;
61879	:douta	=	16'h	c449;
61880	:douta	=	16'h	cc6a;
61881	:douta	=	16'h	cc6a;
61882	:douta	=	16'h	cc6a;
61883	:douta	=	16'h	cc49;
61884	:douta	=	16'h	c449;
61885	:douta	=	16'h	c449;
61886	:douta	=	16'h	cc6a;
61887	:douta	=	16'h	c44a;
61888	:douta	=	16'h	c449;
61889	:douta	=	16'h	c449;
61890	:douta	=	16'h	c449;
61891	:douta	=	16'h	c449;
61892	:douta	=	16'h	c469;
61893	:douta	=	16'h	c449;
61894	:douta	=	16'h	c449;
61895	:douta	=	16'h	c449;
61896	:douta	=	16'h	c429;
61897	:douta	=	16'h	c429;
61898	:douta	=	16'h	c429;
61899	:douta	=	16'h	c44a;
61900	:douta	=	16'h	c429;
61901	:douta	=	16'h	c429;
61902	:douta	=	16'h	c429;
61903	:douta	=	16'h	c429;
61904	:douta	=	16'h	c429;
61905	:douta	=	16'h	c429;
61906	:douta	=	16'h	c42a;
61907	:douta	=	16'h	bc09;
61908	:douta	=	16'h	c40a;
61909	:douta	=	16'h	bc09;
61910	:douta	=	16'h	bc2a;
61911	:douta	=	16'h	bc29;
61912	:douta	=	16'h	bc09;
61913	:douta	=	16'h	bc09;
61914	:douta	=	16'h	bc09;
61915	:douta	=	16'h	bc09;
61916	:douta	=	16'h	bc09;
61917	:douta	=	16'h	bc09;
61918	:douta	=	16'h	bc09;
61919	:douta	=	16'h	bc09;
61920	:douta	=	16'h	bc09;
61921	:douta	=	16'h	bc09;
61922	:douta	=	16'h	bbe9;
61923	:douta	=	16'h	b3e9;
61924	:douta	=	16'h	b3e9;
61925	:douta	=	16'h	bc09;
61926	:douta	=	16'h	b3e9;
61927	:douta	=	16'h	b3e9;
61928	:douta	=	16'h	b3e9;
61929	:douta	=	16'h	b3e9;
61930	:douta	=	16'h	b3e9;
61931	:douta	=	16'h	b3e9;
61932	:douta	=	16'h	abc9;
61933	:douta	=	16'h	b3ca;
61934	:douta	=	16'h	b3c9;
61935	:douta	=	16'h	b3c9;
61936	:douta	=	16'h	abc9;
61937	:douta	=	16'h	abc9;
61938	:douta	=	16'h	aba9;
61939	:douta	=	16'h	abc9;
61940	:douta	=	16'h	abc9;
61941	:douta	=	16'h	abc9;
61942	:douta	=	16'h	aba9;
61943	:douta	=	16'h	abc9;
61944	:douta	=	16'h	aba9;
61945	:douta	=	16'h	aba9;
61946	:douta	=	16'h	aba9;
61947	:douta	=	16'h	a389;
61948	:douta	=	16'h	a389;
61949	:douta	=	16'h	abaa;
61950	:douta	=	16'h	a389;
61951	:douta	=	16'h	a389;
61952	:douta	=	16'h	8496;
61953	:douta	=	16'h	8cd8;
61954	:douta	=	16'h	3186;
61955	:douta	=	16'h	2924;
61956	:douta	=	16'h	3124;
61957	:douta	=	16'h	3124;
61958	:douta	=	16'h	2904;
61959	:douta	=	16'h	2904;
61960	:douta	=	16'h	2904;
61961	:douta	=	16'h	2924;
61962	:douta	=	16'h	2924;
61963	:douta	=	16'h	2904;
61964	:douta	=	16'h	2904;
61965	:douta	=	16'h	20e3;
61966	:douta	=	16'h	20e4;
61967	:douta	=	16'h	20e3;
61968	:douta	=	16'h	2103;
61969	:douta	=	16'h	2103;
61970	:douta	=	16'h	2904;
61971	:douta	=	16'h	20c2;
61972	:douta	=	16'h	20e3;
61973	:douta	=	16'h	20c3;
61974	:douta	=	16'h	28e3;
61975	:douta	=	16'h	28e3;
61976	:douta	=	16'h	28e3;
61977	:douta	=	16'h	28e3;
61978	:douta	=	16'h	28e3;
61979	:douta	=	16'h	28e3;
61980	:douta	=	16'h	2903;
61981	:douta	=	16'h	3103;
61982	:douta	=	16'h	3103;
61983	:douta	=	16'h	3103;
61984	:douta	=	16'h	3103;
61985	:douta	=	16'h	3923;
61986	:douta	=	16'h	4144;
61987	:douta	=	16'h	4144;
61988	:douta	=	16'h	4964;
61989	:douta	=	16'h	4984;
61990	:douta	=	16'h	4964;
61991	:douta	=	16'h	49e7;
61992	:douta	=	16'h	5acd;
61993	:douta	=	16'h	10e5;
61994	:douta	=	16'h	20e5;
61995	:douta	=	16'h	59e4;
61996	:douta	=	16'h	59c4;
61997	:douta	=	16'h	59e4;
61998	:douta	=	16'h	61e4;
61999	:douta	=	16'h	6204;
62000	:douta	=	16'h	6a25;
62001	:douta	=	16'h	6a44;
62002	:douta	=	16'h	7245;
62003	:douta	=	16'h	7245;
62004	:douta	=	16'h	7244;
62005	:douta	=	16'h	83cd;
62006	:douta	=	16'h	938a;
62007	:douta	=	16'h	7a24;
62008	:douta	=	16'h	7a85;
62009	:douta	=	16'h	82a5;
62010	:douta	=	16'h	8285;
62011	:douta	=	16'h	82a5;
62012	:douta	=	16'h	82c6;
62013	:douta	=	16'h	82c6;
62014	:douta	=	16'h	82c6;
62015	:douta	=	16'h	82c6;
62016	:douta	=	16'h	8ae7;
62017	:douta	=	16'h	8b07;
62018	:douta	=	16'h	8ae7;
62019	:douta	=	16'h	8b07;
62020	:douta	=	16'h	9307;
62021	:douta	=	16'h	9327;
62022	:douta	=	16'h	9327;
62023	:douta	=	16'h	9b47;
62024	:douta	=	16'h	9b47;
62025	:douta	=	16'h	9b47;
62026	:douta	=	16'h	9b46;
62027	:douta	=	16'h	9b05;
62028	:douta	=	16'h	9b46;
62029	:douta	=	16'h	9b46;
62030	:douta	=	16'h	a367;
62031	:douta	=	16'h	a388;
62032	:douta	=	16'h	a387;
62033	:douta	=	16'h	aba8;
62034	:douta	=	16'h	b3a8;
62035	:douta	=	16'h	b3c8;
62036	:douta	=	16'h	b3c8;
62037	:douta	=	16'h	b3e8;
62038	:douta	=	16'h	b3e8;
62039	:douta	=	16'h	b3e8;
62040	:douta	=	16'h	b3e8;
62041	:douta	=	16'h	b408;
62042	:douta	=	16'h	bc08;
62043	:douta	=	16'h	bc08;
62044	:douta	=	16'h	bc29;
62045	:douta	=	16'h	bc28;
62046	:douta	=	16'h	bc28;
62047	:douta	=	16'h	bc28;
62048	:douta	=	16'h	c428;
62049	:douta	=	16'h	c428;
62050	:douta	=	16'h	c449;
62051	:douta	=	16'h	c449;
62052	:douta	=	16'h	c449;
62053	:douta	=	16'h	c449;
62054	:douta	=	16'h	c449;
62055	:douta	=	16'h	c449;
62056	:douta	=	16'h	c448;
62057	:douta	=	16'h	c448;
62058	:douta	=	16'h	c448;
62059	:douta	=	16'h	c448;
62060	:douta	=	16'h	c468;
62061	:douta	=	16'h	c448;
62062	:douta	=	16'h	cc69;
62063	:douta	=	16'h	c468;
62064	:douta	=	16'h	cc69;
62065	:douta	=	16'h	c468;
62066	:douta	=	16'h	cc69;
62067	:douta	=	16'h	cc69;
62068	:douta	=	16'h	cc69;
62069	:douta	=	16'h	cc69;
62070	:douta	=	16'h	cc69;
62071	:douta	=	16'h	cc69;
62072	:douta	=	16'h	cc69;
62073	:douta	=	16'h	cc69;
62074	:douta	=	16'h	cc69;
62075	:douta	=	16'h	cc69;
62076	:douta	=	16'h	cc89;
62077	:douta	=	16'h	cc69;
62078	:douta	=	16'h	cc89;
62079	:douta	=	16'h	cc89;
62080	:douta	=	16'h	cc89;
62081	:douta	=	16'h	cc89;
62082	:douta	=	16'h	cc89;
62083	:douta	=	16'h	cc89;
62084	:douta	=	16'h	cc89;
62085	:douta	=	16'h	cc69;
62086	:douta	=	16'h	cc69;
62087	:douta	=	16'h	cc69;
62088	:douta	=	16'h	cc69;
62089	:douta	=	16'h	cc89;
62090	:douta	=	16'h	cc69;
62091	:douta	=	16'h	cc69;
62092	:douta	=	16'h	cc89;
62093	:douta	=	16'h	cc89;
62094	:douta	=	16'h	cc89;
62095	:douta	=	16'h	cc89;
62096	:douta	=	16'h	cc89;
62097	:douta	=	16'h	cc89;
62098	:douta	=	16'h	cc89;
62099	:douta	=	16'h	cc89;
62100	:douta	=	16'h	cc69;
62101	:douta	=	16'h	cc69;
62102	:douta	=	16'h	cc89;
62103	:douta	=	16'h	cc69;
62104	:douta	=	16'h	cc69;
62105	:douta	=	16'h	cc69;
62106	:douta	=	16'h	cc89;
62107	:douta	=	16'h	cc69;
62108	:douta	=	16'h	cc89;
62109	:douta	=	16'h	cc89;
62110	:douta	=	16'h	cc89;
62111	:douta	=	16'h	cc89;
62112	:douta	=	16'h	c489;
62113	:douta	=	16'h	cc69;
62114	:douta	=	16'h	cc68;
62115	:douta	=	16'h	b5d5;
62116	:douta	=	16'h	e655;
62117	:douta	=	16'h	cc69;
62118	:douta	=	16'h	cc6a;
62119	:douta	=	16'h	cc6a;
62120	:douta	=	16'h	cc89;
62121	:douta	=	16'h	cc89;
62122	:douta	=	16'h	cc89;
62123	:douta	=	16'h	cc69;
62124	:douta	=	16'h	cc6a;
62125	:douta	=	16'h	cc69;
62126	:douta	=	16'h	cc69;
62127	:douta	=	16'h	cc49;
62128	:douta	=	16'h	cc49;
62129	:douta	=	16'h	cc69;
62130	:douta	=	16'h	cc69;
62131	:douta	=	16'h	cc69;
62132	:douta	=	16'h	cc69;
62133	:douta	=	16'h	cc69;
62134	:douta	=	16'h	cc69;
62135	:douta	=	16'h	cc49;
62136	:douta	=	16'h	c44a;
62137	:douta	=	16'h	cc6a;
62138	:douta	=	16'h	cc6a;
62139	:douta	=	16'h	c44a;
62140	:douta	=	16'h	c449;
62141	:douta	=	16'h	c449;
62142	:douta	=	16'h	c449;
62143	:douta	=	16'h	c469;
62144	:douta	=	16'h	c449;
62145	:douta	=	16'h	c469;
62146	:douta	=	16'h	c449;
62147	:douta	=	16'h	c449;
62148	:douta	=	16'h	c449;
62149	:douta	=	16'h	c449;
62150	:douta	=	16'h	c449;
62151	:douta	=	16'h	c429;
62152	:douta	=	16'h	c44a;
62153	:douta	=	16'h	c429;
62154	:douta	=	16'h	c429;
62155	:douta	=	16'h	c44a;
62156	:douta	=	16'h	c429;
62157	:douta	=	16'h	c429;
62158	:douta	=	16'h	c429;
62159	:douta	=	16'h	c429;
62160	:douta	=	16'h	bc29;
62161	:douta	=	16'h	c429;
62162	:douta	=	16'h	c40a;
62163	:douta	=	16'h	bc2a;
62164	:douta	=	16'h	bc09;
62165	:douta	=	16'h	bc2a;
62166	:douta	=	16'h	bc2a;
62167	:douta	=	16'h	bc2a;
62168	:douta	=	16'h	bc2a;
62169	:douta	=	16'h	bc09;
62170	:douta	=	16'h	bc2a;
62171	:douta	=	16'h	bc09;
62172	:douta	=	16'h	bc09;
62173	:douta	=	16'h	bc09;
62174	:douta	=	16'h	bc09;
62175	:douta	=	16'h	bc09;
62176	:douta	=	16'h	bc09;
62177	:douta	=	16'h	bbe9;
62178	:douta	=	16'h	bc09;
62179	:douta	=	16'h	bbe9;
62180	:douta	=	16'h	b3e9;
62181	:douta	=	16'h	bbe9;
62182	:douta	=	16'h	bbe9;
62183	:douta	=	16'h	b3e9;
62184	:douta	=	16'h	b3e9;
62185	:douta	=	16'h	b3e9;
62186	:douta	=	16'h	b3e9;
62187	:douta	=	16'h	b3e9;
62188	:douta	=	16'h	b3c9;
62189	:douta	=	16'h	b3ca;
62190	:douta	=	16'h	b3c9;
62191	:douta	=	16'h	b3ca;
62192	:douta	=	16'h	abc9;
62193	:douta	=	16'h	abc9;
62194	:douta	=	16'h	b3c9;
62195	:douta	=	16'h	abc9;
62196	:douta	=	16'h	aba9;
62197	:douta	=	16'h	aba9;
62198	:douta	=	16'h	aba9;
62199	:douta	=	16'h	aba9;
62200	:douta	=	16'h	aba9;
62201	:douta	=	16'h	aba9;
62202	:douta	=	16'h	aba9;
62203	:douta	=	16'h	a389;
62204	:douta	=	16'h	abaa;
62205	:douta	=	16'h	abaa;
62206	:douta	=	16'h	a389;
62207	:douta	=	16'h	a389;
62208	:douta	=	16'h	8cb7;
62209	:douta	=	16'h	4a8b;
62210	:douta	=	16'h	1861;
62211	:douta	=	16'h	2904;
62212	:douta	=	16'h	2924;
62213	:douta	=	16'h	2904;
62214	:douta	=	16'h	3124;
62215	:douta	=	16'h	2904;
62216	:douta	=	16'h	2904;
62217	:douta	=	16'h	2904;
62218	:douta	=	16'h	2924;
62219	:douta	=	16'h	2904;
62220	:douta	=	16'h	2904;
62221	:douta	=	16'h	2904;
62222	:douta	=	16'h	20e3;
62223	:douta	=	16'h	20e3;
62224	:douta	=	16'h	2103;
62225	:douta	=	16'h	20e3;
62226	:douta	=	16'h	28e3;
62227	:douta	=	16'h	20c2;
62228	:douta	=	16'h	20e3;
62229	:douta	=	16'h	20c3;
62230	:douta	=	16'h	20e3;
62231	:douta	=	16'h	28e3;
62232	:douta	=	16'h	28e3;
62233	:douta	=	16'h	28e3;
62234	:douta	=	16'h	28e3;
62235	:douta	=	16'h	2903;
62236	:douta	=	16'h	2903;
62237	:douta	=	16'h	3103;
62238	:douta	=	16'h	3124;
62239	:douta	=	16'h	3903;
62240	:douta	=	16'h	3923;
62241	:douta	=	16'h	3923;
62242	:douta	=	16'h	3923;
62243	:douta	=	16'h	4144;
62244	:douta	=	16'h	4964;
62245	:douta	=	16'h	4964;
62246	:douta	=	16'h	4984;
62247	:douta	=	16'h	4a28;
62248	:douta	=	16'h	528b;
62249	:douta	=	16'h	1085;
62250	:douta	=	16'h	3124;
62251	:douta	=	16'h	59c4;
62252	:douta	=	16'h	61e4;
62253	:douta	=	16'h	59e4;
62254	:douta	=	16'h	6a05;
62255	:douta	=	16'h	6204;
62256	:douta	=	16'h	6a24;
62257	:douta	=	16'h	6a25;
62258	:douta	=	16'h	7244;
62259	:douta	=	16'h	7245;
62260	:douta	=	16'h	7224;
62261	:douta	=	16'h	9491;
62262	:douta	=	16'h	7aa5;
62263	:douta	=	16'h	7244;
62264	:douta	=	16'h	82a5;
62265	:douta	=	16'h	82a5;
62266	:douta	=	16'h	8285;
62267	:douta	=	16'h	82a6;
62268	:douta	=	16'h	8ac6;
62269	:douta	=	16'h	82c6;
62270	:douta	=	16'h	8ac6;
62271	:douta	=	16'h	8ae6;
62272	:douta	=	16'h	9307;
62273	:douta	=	16'h	8ac6;
62274	:douta	=	16'h	8ae7;
62275	:douta	=	16'h	9307;
62276	:douta	=	16'h	9307;
62277	:douta	=	16'h	9327;
62278	:douta	=	16'h	9327;
62279	:douta	=	16'h	9b47;
62280	:douta	=	16'h	9b47;
62281	:douta	=	16'h	9b47;
62282	:douta	=	16'h	a368;
62283	:douta	=	16'h	a368;
62284	:douta	=	16'h	9b67;
62285	:douta	=	16'h	a368;
62286	:douta	=	16'h	a368;
62287	:douta	=	16'h	a388;
62288	:douta	=	16'h	a388;
62289	:douta	=	16'h	aba8;
62290	:douta	=	16'h	aba8;
62291	:douta	=	16'h	b3c8;
62292	:douta	=	16'h	b3c8;
62293	:douta	=	16'h	b3e8;
62294	:douta	=	16'h	b3e8;
62295	:douta	=	16'h	b3e8;
62296	:douta	=	16'h	bbe8;
62297	:douta	=	16'h	bbe8;
62298	:douta	=	16'h	bc08;
62299	:douta	=	16'h	bc08;
62300	:douta	=	16'h	bc29;
62301	:douta	=	16'h	bc08;
62302	:douta	=	16'h	bc29;
62303	:douta	=	16'h	bc28;
62304	:douta	=	16'h	bc29;
62305	:douta	=	16'h	c429;
62306	:douta	=	16'h	c449;
62307	:douta	=	16'h	c449;
62308	:douta	=	16'h	c449;
62309	:douta	=	16'h	c449;
62310	:douta	=	16'h	c449;
62311	:douta	=	16'h	c449;
62312	:douta	=	16'h	c449;
62313	:douta	=	16'h	c449;
62314	:douta	=	16'h	c448;
62315	:douta	=	16'h	c468;
62316	:douta	=	16'h	cc49;
62317	:douta	=	16'h	cc49;
62318	:douta	=	16'h	cc69;
62319	:douta	=	16'h	cc69;
62320	:douta	=	16'h	cc69;
62321	:douta	=	16'h	cc69;
62322	:douta	=	16'h	cc69;
62323	:douta	=	16'h	cc69;
62324	:douta	=	16'h	cc69;
62325	:douta	=	16'h	cc69;
62326	:douta	=	16'h	cc69;
62327	:douta	=	16'h	cc69;
62328	:douta	=	16'h	cc69;
62329	:douta	=	16'h	cc69;
62330	:douta	=	16'h	cc69;
62331	:douta	=	16'h	cc89;
62332	:douta	=	16'h	cc69;
62333	:douta	=	16'h	cc69;
62334	:douta	=	16'h	cc89;
62335	:douta	=	16'h	cc69;
62336	:douta	=	16'h	cc89;
62337	:douta	=	16'h	cc89;
62338	:douta	=	16'h	cc69;
62339	:douta	=	16'h	cc89;
62340	:douta	=	16'h	cc69;
62341	:douta	=	16'h	cc89;
62342	:douta	=	16'h	cc89;
62343	:douta	=	16'h	cc69;
62344	:douta	=	16'h	cc69;
62345	:douta	=	16'h	cc69;
62346	:douta	=	16'h	cc89;
62347	:douta	=	16'h	cc89;
62348	:douta	=	16'h	cc89;
62349	:douta	=	16'h	cc89;
62350	:douta	=	16'h	cc89;
62351	:douta	=	16'h	cc69;
62352	:douta	=	16'h	cc89;
62353	:douta	=	16'h	cc69;
62354	:douta	=	16'h	cc89;
62355	:douta	=	16'h	cc89;
62356	:douta	=	16'h	cc89;
62357	:douta	=	16'h	cc69;
62358	:douta	=	16'h	cc69;
62359	:douta	=	16'h	cc69;
62360	:douta	=	16'h	cc89;
62361	:douta	=	16'h	cc69;
62362	:douta	=	16'h	cc69;
62363	:douta	=	16'h	cc69;
62364	:douta	=	16'h	cc69;
62365	:douta	=	16'h	cc89;
62366	:douta	=	16'h	cc89;
62367	:douta	=	16'h	c489;
62368	:douta	=	16'h	cc6a;
62369	:douta	=	16'h	cc69;
62370	:douta	=	16'h	cc69;
62371	:douta	=	16'h	b5d5;
62372	:douta	=	16'h	e675;
62373	:douta	=	16'h	c448;
62374	:douta	=	16'h	c469;
62375	:douta	=	16'h	cc69;
62376	:douta	=	16'h	cc69;
62377	:douta	=	16'h	cc6a;
62378	:douta	=	16'h	cc69;
62379	:douta	=	16'h	cc69;
62380	:douta	=	16'h	cc6a;
62381	:douta	=	16'h	cc8a;
62382	:douta	=	16'h	cc6a;
62383	:douta	=	16'h	cc69;
62384	:douta	=	16'h	cc49;
62385	:douta	=	16'h	cc6a;
62386	:douta	=	16'h	cc6a;
62387	:douta	=	16'h	cc6a;
62388	:douta	=	16'h	cc69;
62389	:douta	=	16'h	cc49;
62390	:douta	=	16'h	cc49;
62391	:douta	=	16'h	cc6a;
62392	:douta	=	16'h	cc6a;
62393	:douta	=	16'h	c449;
62394	:douta	=	16'h	c449;
62395	:douta	=	16'h	c449;
62396	:douta	=	16'h	c46a;
62397	:douta	=	16'h	c449;
62398	:douta	=	16'h	c469;
62399	:douta	=	16'h	c449;
62400	:douta	=	16'h	c469;
62401	:douta	=	16'h	c449;
62402	:douta	=	16'h	c449;
62403	:douta	=	16'h	c449;
62404	:douta	=	16'h	c44a;
62405	:douta	=	16'h	c44a;
62406	:douta	=	16'h	c44a;
62407	:douta	=	16'h	c44a;
62408	:douta	=	16'h	c44a;
62409	:douta	=	16'h	c429;
62410	:douta	=	16'h	c429;
62411	:douta	=	16'h	c42a;
62412	:douta	=	16'h	c42a;
62413	:douta	=	16'h	c40a;
62414	:douta	=	16'h	bc2a;
62415	:douta	=	16'h	bc29;
62416	:douta	=	16'h	bc09;
62417	:douta	=	16'h	bc09;
62418	:douta	=	16'h	bc0a;
62419	:douta	=	16'h	bc0a;
62420	:douta	=	16'h	bc2a;
62421	:douta	=	16'h	bc09;
62422	:douta	=	16'h	bc09;
62423	:douta	=	16'h	bc2a;
62424	:douta	=	16'h	bc09;
62425	:douta	=	16'h	bc09;
62426	:douta	=	16'h	bc09;
62427	:douta	=	16'h	bc09;
62428	:douta	=	16'h	bc09;
62429	:douta	=	16'h	bc09;
62430	:douta	=	16'h	bc09;
62431	:douta	=	16'h	bc09;
62432	:douta	=	16'h	bc09;
62433	:douta	=	16'h	bc09;
62434	:douta	=	16'h	bc09;
62435	:douta	=	16'h	bc09;
62436	:douta	=	16'h	bbe9;
62437	:douta	=	16'h	bbe9;
62438	:douta	=	16'h	b3e9;
62439	:douta	=	16'h	b3e9;
62440	:douta	=	16'h	b3e9;
62441	:douta	=	16'h	b3c9;
62442	:douta	=	16'h	b3e9;
62443	:douta	=	16'h	b3c9;
62444	:douta	=	16'h	b3c9;
62445	:douta	=	16'h	abc9;
62446	:douta	=	16'h	b3ca;
62447	:douta	=	16'h	aba9;
62448	:douta	=	16'h	b3ca;
62449	:douta	=	16'h	b3ca;
62450	:douta	=	16'h	abc9;
62451	:douta	=	16'h	abc9;
62452	:douta	=	16'h	abc9;
62453	:douta	=	16'h	abc9;
62454	:douta	=	16'h	aba9;
62455	:douta	=	16'h	aba9;
62456	:douta	=	16'h	aba9;
62457	:douta	=	16'h	aba9;
62458	:douta	=	16'h	aba9;
62459	:douta	=	16'h	a389;
62460	:douta	=	16'h	ab89;
62461	:douta	=	16'h	a389;
62462	:douta	=	16'h	ab8a;
62463	:douta	=	16'h	a389;
62464	:douta	=	16'h	9519;
62465	:douta	=	16'h	2925;
62466	:douta	=	16'h	28e3;
62467	:douta	=	16'h	2904;
62468	:douta	=	16'h	2924;
62469	:douta	=	16'h	3124;
62470	:douta	=	16'h	2904;
62471	:douta	=	16'h	3124;
62472	:douta	=	16'h	2904;
62473	:douta	=	16'h	2904;
62474	:douta	=	16'h	2904;
62475	:douta	=	16'h	2904;
62476	:douta	=	16'h	28e4;
62477	:douta	=	16'h	2904;
62478	:douta	=	16'h	20e3;
62479	:douta	=	16'h	2103;
62480	:douta	=	16'h	20e3;
62481	:douta	=	16'h	20e4;
62482	:douta	=	16'h	20e3;
62483	:douta	=	16'h	20c3;
62484	:douta	=	16'h	20c3;
62485	:douta	=	16'h	20c3;
62486	:douta	=	16'h	28e3;
62487	:douta	=	16'h	28e3;
62488	:douta	=	16'h	28e3;
62489	:douta	=	16'h	28e3;
62490	:douta	=	16'h	2903;
62491	:douta	=	16'h	3123;
62492	:douta	=	16'h	3103;
62493	:douta	=	16'h	3103;
62494	:douta	=	16'h	3103;
62495	:douta	=	16'h	3903;
62496	:douta	=	16'h	3923;
62497	:douta	=	16'h	3923;
62498	:douta	=	16'h	3944;
62499	:douta	=	16'h	4144;
62500	:douta	=	16'h	4964;
62501	:douta	=	16'h	4964;
62502	:douta	=	16'h	51a5;
62503	:douta	=	16'h	4a49;
62504	:douta	=	16'h	4a2a;
62505	:douta	=	16'h	1084;
62506	:douta	=	16'h	3945;
62507	:douta	=	16'h	59c4;
62508	:douta	=	16'h	59e4;
62509	:douta	=	16'h	61e5;
62510	:douta	=	16'h	6a05;
62511	:douta	=	16'h	6a05;
62512	:douta	=	16'h	6a24;
62513	:douta	=	16'h	6a24;
62514	:douta	=	16'h	6a24;
62515	:douta	=	16'h	7245;
62516	:douta	=	16'h	7224;
62517	:douta	=	16'h	a4f2;
62518	:douta	=	16'h	7244;
62519	:douta	=	16'h	7a64;
62520	:douta	=	16'h	7a85;
62521	:douta	=	16'h	82a6;
62522	:douta	=	16'h	82a6;
62523	:douta	=	16'h	82a6;
62524	:douta	=	16'h	82c6;
62525	:douta	=	16'h	82c6;
62526	:douta	=	16'h	82a6;
62527	:douta	=	16'h	82c6;
62528	:douta	=	16'h	8ae7;
62529	:douta	=	16'h	8ae7;
62530	:douta	=	16'h	8ae7;
62531	:douta	=	16'h	8b07;
62532	:douta	=	16'h	9307;
62533	:douta	=	16'h	9327;
62534	:douta	=	16'h	9327;
62535	:douta	=	16'h	9327;
62536	:douta	=	16'h	9b47;
62537	:douta	=	16'h	9b47;
62538	:douta	=	16'h	a368;
62539	:douta	=	16'h	9b67;
62540	:douta	=	16'h	a368;
62541	:douta	=	16'h	9b67;
62542	:douta	=	16'h	a388;
62543	:douta	=	16'h	ab88;
62544	:douta	=	16'h	a388;
62545	:douta	=	16'h	aba8;
62546	:douta	=	16'h	aba8;
62547	:douta	=	16'h	b3c8;
62548	:douta	=	16'h	b3e8;
62549	:douta	=	16'h	b3e8;
62550	:douta	=	16'h	b3e8;
62551	:douta	=	16'h	bbe8;
62552	:douta	=	16'h	b3e8;
62553	:douta	=	16'h	bbe8;
62554	:douta	=	16'h	bc08;
62555	:douta	=	16'h	bc08;
62556	:douta	=	16'h	bc08;
62557	:douta	=	16'h	bc28;
62558	:douta	=	16'h	bc29;
62559	:douta	=	16'h	c428;
62560	:douta	=	16'h	c429;
62561	:douta	=	16'h	c449;
62562	:douta	=	16'h	c449;
62563	:douta	=	16'h	c449;
62564	:douta	=	16'h	c449;
62565	:douta	=	16'h	c449;
62566	:douta	=	16'h	c449;
62567	:douta	=	16'h	c449;
62568	:douta	=	16'h	c449;
62569	:douta	=	16'h	c449;
62570	:douta	=	16'h	c468;
62571	:douta	=	16'h	c448;
62572	:douta	=	16'h	cc49;
62573	:douta	=	16'h	cc69;
62574	:douta	=	16'h	cc69;
62575	:douta	=	16'h	cc69;
62576	:douta	=	16'h	cc69;
62577	:douta	=	16'h	cc6a;
62578	:douta	=	16'h	cc6a;
62579	:douta	=	16'h	cc69;
62580	:douta	=	16'h	cc69;
62581	:douta	=	16'h	cc69;
62582	:douta	=	16'h	cc69;
62583	:douta	=	16'h	cc69;
62584	:douta	=	16'h	cc69;
62585	:douta	=	16'h	cc6a;
62586	:douta	=	16'h	cc69;
62587	:douta	=	16'h	cc89;
62588	:douta	=	16'h	cc89;
62589	:douta	=	16'h	cc69;
62590	:douta	=	16'h	cc8a;
62591	:douta	=	16'h	cc6a;
62592	:douta	=	16'h	cc89;
62593	:douta	=	16'h	cc89;
62594	:douta	=	16'h	cc89;
62595	:douta	=	16'h	cc89;
62596	:douta	=	16'h	cc89;
62597	:douta	=	16'h	cc89;
62598	:douta	=	16'h	cc69;
62599	:douta	=	16'h	cc69;
62600	:douta	=	16'h	cc89;
62601	:douta	=	16'h	cc89;
62602	:douta	=	16'h	cc89;
62603	:douta	=	16'h	cc89;
62604	:douta	=	16'h	cc89;
62605	:douta	=	16'h	cc89;
62606	:douta	=	16'h	cc89;
62607	:douta	=	16'h	cc69;
62608	:douta	=	16'h	cc6a;
62609	:douta	=	16'h	cc69;
62610	:douta	=	16'h	cc89;
62611	:douta	=	16'h	cc69;
62612	:douta	=	16'h	cc89;
62613	:douta	=	16'h	cc89;
62614	:douta	=	16'h	cc69;
62615	:douta	=	16'h	cc69;
62616	:douta	=	16'h	cc69;
62617	:douta	=	16'h	cc69;
62618	:douta	=	16'h	cc69;
62619	:douta	=	16'h	cc89;
62620	:douta	=	16'h	cc89;
62621	:douta	=	16'h	cc89;
62622	:douta	=	16'h	cc69;
62623	:douta	=	16'h	c489;
62624	:douta	=	16'h	cc6a;
62625	:douta	=	16'h	cc69;
62626	:douta	=	16'h	cc69;
62627	:douta	=	16'h	b5b5;
62628	:douta	=	16'h	e655;
62629	:douta	=	16'h	cc69;
62630	:douta	=	16'h	c469;
62631	:douta	=	16'h	c469;
62632	:douta	=	16'h	cc69;
62633	:douta	=	16'h	cc69;
62634	:douta	=	16'h	cc69;
62635	:douta	=	16'h	cc69;
62636	:douta	=	16'h	cc8a;
62637	:douta	=	16'h	cc6a;
62638	:douta	=	16'h	cc6a;
62639	:douta	=	16'h	cc49;
62640	:douta	=	16'h	cc69;
62641	:douta	=	16'h	cc6a;
62642	:douta	=	16'h	cc6a;
62643	:douta	=	16'h	cc6a;
62644	:douta	=	16'h	cc49;
62645	:douta	=	16'h	cc69;
62646	:douta	=	16'h	cc69;
62647	:douta	=	16'h	c44a;
62648	:douta	=	16'h	c44a;
62649	:douta	=	16'h	c46a;
62650	:douta	=	16'h	c44a;
62651	:douta	=	16'h	c46a;
62652	:douta	=	16'h	c469;
62653	:douta	=	16'h	c469;
62654	:douta	=	16'h	c449;
62655	:douta	=	16'h	c46a;
62656	:douta	=	16'h	c469;
62657	:douta	=	16'h	c449;
62658	:douta	=	16'h	c449;
62659	:douta	=	16'h	c449;
62660	:douta	=	16'h	c44a;
62661	:douta	=	16'h	c44a;
62662	:douta	=	16'h	c44a;
62663	:douta	=	16'h	c44a;
62664	:douta	=	16'h	c429;
62665	:douta	=	16'h	c429;
62666	:douta	=	16'h	c429;
62667	:douta	=	16'h	c42a;
62668	:douta	=	16'h	c42a;
62669	:douta	=	16'h	c42a;
62670	:douta	=	16'h	c42a;
62671	:douta	=	16'h	bc29;
62672	:douta	=	16'h	bc29;
62673	:douta	=	16'h	bc29;
62674	:douta	=	16'h	bc09;
62675	:douta	=	16'h	bc09;
62676	:douta	=	16'h	bc2a;
62677	:douta	=	16'h	bc09;
62678	:douta	=	16'h	bc2a;
62679	:douta	=	16'h	bc09;
62680	:douta	=	16'h	bc09;
62681	:douta	=	16'h	bc09;
62682	:douta	=	16'h	bc09;
62683	:douta	=	16'h	bc2a;
62684	:douta	=	16'h	bc0a;
62685	:douta	=	16'h	bc09;
62686	:douta	=	16'h	bc09;
62687	:douta	=	16'h	bc09;
62688	:douta	=	16'h	bc09;
62689	:douta	=	16'h	bc09;
62690	:douta	=	16'h	bbe9;
62691	:douta	=	16'h	bbe9;
62692	:douta	=	16'h	bbe9;
62693	:douta	=	16'h	b3e9;
62694	:douta	=	16'h	b3e9;
62695	:douta	=	16'h	b3e9;
62696	:douta	=	16'h	b3e9;
62697	:douta	=	16'h	b3e9;
62698	:douta	=	16'h	b3c9;
62699	:douta	=	16'h	b3e9;
62700	:douta	=	16'h	b3c9;
62701	:douta	=	16'h	abc9;
62702	:douta	=	16'h	b3ca;
62703	:douta	=	16'h	abc9;
62704	:douta	=	16'h	b3c9;
62705	:douta	=	16'h	aba9;
62706	:douta	=	16'h	abc9;
62707	:douta	=	16'h	abc9;
62708	:douta	=	16'h	aba9;
62709	:douta	=	16'h	aba9;
62710	:douta	=	16'h	aba9;
62711	:douta	=	16'h	aba9;
62712	:douta	=	16'h	ab89;
62713	:douta	=	16'h	aba9;
62714	:douta	=	16'h	ab89;
62715	:douta	=	16'h	a389;
62716	:douta	=	16'h	ab89;
62717	:douta	=	16'h	a389;
62718	:douta	=	16'h	a38a;
62719	:douta	=	16'h	a389;
62720	:douta	=	16'h	9539;
62721	:douta	=	16'h	1881;
62722	:douta	=	16'h	2924;
62723	:douta	=	16'h	2924;
62724	:douta	=	16'h	3124;
62725	:douta	=	16'h	3124;
62726	:douta	=	16'h	3124;
62727	:douta	=	16'h	3124;
62728	:douta	=	16'h	2904;
62729	:douta	=	16'h	2904;
62730	:douta	=	16'h	2904;
62731	:douta	=	16'h	2904;
62732	:douta	=	16'h	2904;
62733	:douta	=	16'h	2103;
62734	:douta	=	16'h	20e4;
62735	:douta	=	16'h	2103;
62736	:douta	=	16'h	2904;
62737	:douta	=	16'h	2904;
62738	:douta	=	16'h	20a3;
62739	:douta	=	16'h	20c3;
62740	:douta	=	16'h	20e3;
62741	:douta	=	16'h	28e3;
62742	:douta	=	16'h	28e3;
62743	:douta	=	16'h	28e3;
62744	:douta	=	16'h	2904;
62745	:douta	=	16'h	28e3;
62746	:douta	=	16'h	28e3;
62747	:douta	=	16'h	28e3;
62748	:douta	=	16'h	3103;
62749	:douta	=	16'h	3123;
62750	:douta	=	16'h	3123;
62751	:douta	=	16'h	3923;
62752	:douta	=	16'h	3923;
62753	:douta	=	16'h	3943;
62754	:douta	=	16'h	3944;
62755	:douta	=	16'h	4144;
62756	:douta	=	16'h	4164;
62757	:douta	=	16'h	4984;
62758	:douta	=	16'h	4964;
62759	:douta	=	16'h	528b;
62760	:douta	=	16'h	39c8;
62761	:douta	=	16'h	18a4;
62762	:douta	=	16'h	51a5;
62763	:douta	=	16'h	59e4;
62764	:douta	=	16'h	59c5;
62765	:douta	=	16'h	61e4;
62766	:douta	=	16'h	6204;
62767	:douta	=	16'h	6204;
62768	:douta	=	16'h	6a25;
62769	:douta	=	16'h	6a25;
62770	:douta	=	16'h	7245;
62771	:douta	=	16'h	7245;
62772	:douta	=	16'h	7224;
62773	:douta	=	16'h	b594;
62774	:douta	=	16'h	7203;
62775	:douta	=	16'h	7a85;
62776	:douta	=	16'h	82a5;
62777	:douta	=	16'h	82a5;
62778	:douta	=	16'h	82a6;
62779	:douta	=	16'h	82c6;
62780	:douta	=	16'h	82c6;
62781	:douta	=	16'h	82c6;
62782	:douta	=	16'h	8ac6;
62783	:douta	=	16'h	8b07;
62784	:douta	=	16'h	8ae7;
62785	:douta	=	16'h	8b07;
62786	:douta	=	16'h	8ae7;
62787	:douta	=	16'h	8b07;
62788	:douta	=	16'h	9307;
62789	:douta	=	16'h	9328;
62790	:douta	=	16'h	9b28;
62791	:douta	=	16'h	9b47;
62792	:douta	=	16'h	9b47;
62793	:douta	=	16'h	9b68;
62794	:douta	=	16'h	9b47;
62795	:douta	=	16'h	9b67;
62796	:douta	=	16'h	9b67;
62797	:douta	=	16'h	9b67;
62798	:douta	=	16'h	a368;
62799	:douta	=	16'h	a367;
62800	:douta	=	16'h	a388;
62801	:douta	=	16'h	ab87;
62802	:douta	=	16'h	abc8;
62803	:douta	=	16'h	b3c8;
62804	:douta	=	16'h	b3e8;
62805	:douta	=	16'h	b3e8;
62806	:douta	=	16'h	bc09;
62807	:douta	=	16'h	b3e8;
62808	:douta	=	16'h	bbe8;
62809	:douta	=	16'h	bbe8;
62810	:douta	=	16'h	bbe8;
62811	:douta	=	16'h	bc28;
62812	:douta	=	16'h	bc29;
62813	:douta	=	16'h	c429;
62814	:douta	=	16'h	c429;
62815	:douta	=	16'h	c449;
62816	:douta	=	16'h	c449;
62817	:douta	=	16'h	c429;
62818	:douta	=	16'h	c449;
62819	:douta	=	16'h	c429;
62820	:douta	=	16'h	c449;
62821	:douta	=	16'h	c429;
62822	:douta	=	16'h	c429;
62823	:douta	=	16'h	c449;
62824	:douta	=	16'h	c428;
62825	:douta	=	16'h	c449;
62826	:douta	=	16'h	cc49;
62827	:douta	=	16'h	cc49;
62828	:douta	=	16'h	cc69;
62829	:douta	=	16'h	cc69;
62830	:douta	=	16'h	c469;
62831	:douta	=	16'h	cc49;
62832	:douta	=	16'h	cc69;
62833	:douta	=	16'h	cc49;
62834	:douta	=	16'h	cc49;
62835	:douta	=	16'h	cc69;
62836	:douta	=	16'h	cc69;
62837	:douta	=	16'h	cc69;
62838	:douta	=	16'h	cc6a;
62839	:douta	=	16'h	cc69;
62840	:douta	=	16'h	cc6a;
62841	:douta	=	16'h	cc6a;
62842	:douta	=	16'h	cc6a;
62843	:douta	=	16'h	cc6a;
62844	:douta	=	16'h	cc6a;
62845	:douta	=	16'h	cc6a;
62846	:douta	=	16'h	cc6a;
62847	:douta	=	16'h	cc6a;
62848	:douta	=	16'h	cc8a;
62849	:douta	=	16'h	cc6a;
62850	:douta	=	16'h	cc89;
62851	:douta	=	16'h	cc69;
62852	:douta	=	16'h	cc69;
62853	:douta	=	16'h	cc69;
62854	:douta	=	16'h	cc89;
62855	:douta	=	16'h	cc89;
62856	:douta	=	16'h	cc69;
62857	:douta	=	16'h	cc89;
62858	:douta	=	16'h	cc89;
62859	:douta	=	16'h	cc69;
62860	:douta	=	16'h	cc69;
62861	:douta	=	16'h	cc69;
62862	:douta	=	16'h	cc6a;
62863	:douta	=	16'h	cc6a;
62864	:douta	=	16'h	cc6a;
62865	:douta	=	16'h	cc69;
62866	:douta	=	16'h	cc69;
62867	:douta	=	16'h	cc69;
62868	:douta	=	16'h	cc89;
62869	:douta	=	16'h	cc69;
62870	:douta	=	16'h	cc89;
62871	:douta	=	16'h	cc6a;
62872	:douta	=	16'h	cc6a;
62873	:douta	=	16'h	cc6a;
62874	:douta	=	16'h	cc6a;
62875	:douta	=	16'h	cc89;
62876	:douta	=	16'h	cc89;
62877	:douta	=	16'h	cc69;
62878	:douta	=	16'h	c489;
62879	:douta	=	16'h	cc6a;
62880	:douta	=	16'h	cc6a;
62881	:douta	=	16'h	cc69;
62882	:douta	=	16'h	cc69;
62883	:douta	=	16'h	b5b5;
62884	:douta	=	16'h	e655;
62885	:douta	=	16'h	c468;
62886	:douta	=	16'h	cc6a;
62887	:douta	=	16'h	cc6a;
62888	:douta	=	16'h	cc6a;
62889	:douta	=	16'h	cc6a;
62890	:douta	=	16'h	cc69;
62891	:douta	=	16'h	cc69;
62892	:douta	=	16'h	cc49;
62893	:douta	=	16'h	cc8a;
62894	:douta	=	16'h	cc69;
62895	:douta	=	16'h	cc49;
62896	:douta	=	16'h	cc49;
62897	:douta	=	16'h	cc6a;
62898	:douta	=	16'h	cc6a;
62899	:douta	=	16'h	cc6a;
62900	:douta	=	16'h	cc69;
62901	:douta	=	16'h	cc69;
62902	:douta	=	16'h	c469;
62903	:douta	=	16'h	c449;
62904	:douta	=	16'h	c449;
62905	:douta	=	16'h	c469;
62906	:douta	=	16'h	c449;
62907	:douta	=	16'h	c449;
62908	:douta	=	16'h	c449;
62909	:douta	=	16'h	c44a;
62910	:douta	=	16'h	c449;
62911	:douta	=	16'h	c449;
62912	:douta	=	16'h	c449;
62913	:douta	=	16'h	c469;
62914	:douta	=	16'h	c469;
62915	:douta	=	16'h	c44a;
62916	:douta	=	16'h	c44a;
62917	:douta	=	16'h	c44a;
62918	:douta	=	16'h	c44a;
62919	:douta	=	16'h	c429;
62920	:douta	=	16'h	c44a;
62921	:douta	=	16'h	c429;
62922	:douta	=	16'h	c42a;
62923	:douta	=	16'h	c42a;
62924	:douta	=	16'h	c42a;
62925	:douta	=	16'h	bc2a;
62926	:douta	=	16'h	bc2a;
62927	:douta	=	16'h	bc29;
62928	:douta	=	16'h	bc09;
62929	:douta	=	16'h	bc09;
62930	:douta	=	16'h	bc2a;
62931	:douta	=	16'h	bc29;
62932	:douta	=	16'h	bc09;
62933	:douta	=	16'h	bc2a;
62934	:douta	=	16'h	bc2a;
62935	:douta	=	16'h	bc09;
62936	:douta	=	16'h	bc09;
62937	:douta	=	16'h	bc09;
62938	:douta	=	16'h	bc09;
62939	:douta	=	16'h	bc09;
62940	:douta	=	16'h	bc09;
62941	:douta	=	16'h	bc09;
62942	:douta	=	16'h	bc09;
62943	:douta	=	16'h	bbe9;
62944	:douta	=	16'h	bc09;
62945	:douta	=	16'h	bbe9;
62946	:douta	=	16'h	bbe9;
62947	:douta	=	16'h	bbe9;
62948	:douta	=	16'h	bbe9;
62949	:douta	=	16'h	bbe9;
62950	:douta	=	16'h	b3e9;
62951	:douta	=	16'h	b3e9;
62952	:douta	=	16'h	b3e9;
62953	:douta	=	16'h	b3e9;
62954	:douta	=	16'h	b3c9;
62955	:douta	=	16'h	b3ca;
62956	:douta	=	16'h	b3c9;
62957	:douta	=	16'h	b3c9;
62958	:douta	=	16'h	abc9;
62959	:douta	=	16'h	b3c9;
62960	:douta	=	16'h	abc9;
62961	:douta	=	16'h	aba9;
62962	:douta	=	16'h	abc9;
62963	:douta	=	16'h	aba9;
62964	:douta	=	16'h	aba9;
62965	:douta	=	16'h	aba9;
62966	:douta	=	16'h	aba9;
62967	:douta	=	16'h	aba9;
62968	:douta	=	16'h	aba9;
62969	:douta	=	16'h	aba9;
62970	:douta	=	16'h	a389;
62971	:douta	=	16'h	a389;
62972	:douta	=	16'h	a389;
62973	:douta	=	16'h	a389;
62974	:douta	=	16'h	a38a;
62975	:douta	=	16'h	a369;
62976	:douta	=	16'h	7c55;
62977	:douta	=	16'h	28e3;
62978	:douta	=	16'h	3145;
62979	:douta	=	16'h	2925;
62980	:douta	=	16'h	3124;
62981	:douta	=	16'h	3124;
62982	:douta	=	16'h	3124;
62983	:douta	=	16'h	3124;
62984	:douta	=	16'h	2904;
62985	:douta	=	16'h	2904;
62986	:douta	=	16'h	2904;
62987	:douta	=	16'h	2904;
62988	:douta	=	16'h	28e4;
62989	:douta	=	16'h	28e3;
62990	:douta	=	16'h	20e3;
62991	:douta	=	16'h	28e3;
62992	:douta	=	16'h	2904;
62993	:douta	=	16'h	2904;
62994	:douta	=	16'h	20a2;
62995	:douta	=	16'h	20e3;
62996	:douta	=	16'h	20e3;
62997	:douta	=	16'h	28e3;
62998	:douta	=	16'h	28e3;
62999	:douta	=	16'h	2903;
63000	:douta	=	16'h	2903;
63001	:douta	=	16'h	2903;
63002	:douta	=	16'h	2903;
63003	:douta	=	16'h	28e3;
63004	:douta	=	16'h	3103;
63005	:douta	=	16'h	3123;
63006	:douta	=	16'h	3123;
63007	:douta	=	16'h	3923;
63008	:douta	=	16'h	3923;
63009	:douta	=	16'h	3943;
63010	:douta	=	16'h	3943;
63011	:douta	=	16'h	4144;
63012	:douta	=	16'h	4964;
63013	:douta	=	16'h	4964;
63014	:douta	=	16'h	4984;
63015	:douta	=	16'h	5a8b;
63016	:douta	=	16'h	3987;
63017	:douta	=	16'h	20e4;
63018	:douta	=	16'h	59c5;
63019	:douta	=	16'h	59e4;
63020	:douta	=	16'h	59c4;
63021	:douta	=	16'h	6205;
63022	:douta	=	16'h	6204;
63023	:douta	=	16'h	6204;
63024	:douta	=	16'h	6a25;
63025	:douta	=	16'h	7245;
63026	:douta	=	16'h	7245;
63027	:douta	=	16'h	7225;
63028	:douta	=	16'h	7224;
63029	:douta	=	16'h	b594;
63030	:douta	=	16'h	7224;
63031	:douta	=	16'h	7a84;
63032	:douta	=	16'h	7a85;
63033	:douta	=	16'h	7a85;
63034	:douta	=	16'h	82a6;
63035	:douta	=	16'h	82c6;
63036	:douta	=	16'h	82c6;
63037	:douta	=	16'h	82c6;
63038	:douta	=	16'h	82c6;
63039	:douta	=	16'h	8ae7;
63040	:douta	=	16'h	8b07;
63041	:douta	=	16'h	8b07;
63042	:douta	=	16'h	9307;
63043	:douta	=	16'h	9307;
63044	:douta	=	16'h	9327;
63045	:douta	=	16'h	9307;
63046	:douta	=	16'h	9328;
63047	:douta	=	16'h	9b47;
63048	:douta	=	16'h	9b68;
63049	:douta	=	16'h	9b68;
63050	:douta	=	16'h	9b67;
63051	:douta	=	16'h	9b67;
63052	:douta	=	16'h	a368;
63053	:douta	=	16'h	9b67;
63054	:douta	=	16'h	a388;
63055	:douta	=	16'h	a388;
63056	:douta	=	16'h	a388;
63057	:douta	=	16'h	aba8;
63058	:douta	=	16'h	aba8;
63059	:douta	=	16'h	b3c8;
63060	:douta	=	16'h	b3e7;
63061	:douta	=	16'h	b3e8;
63062	:douta	=	16'h	bc08;
63063	:douta	=	16'h	bbe8;
63064	:douta	=	16'h	bc09;
63065	:douta	=	16'h	bbe8;
63066	:douta	=	16'h	bc09;
63067	:douta	=	16'h	bc08;
63068	:douta	=	16'h	bc29;
63069	:douta	=	16'h	bc29;
63070	:douta	=	16'h	bc29;
63071	:douta	=	16'h	c429;
63072	:douta	=	16'h	c449;
63073	:douta	=	16'h	c449;
63074	:douta	=	16'h	c449;
63075	:douta	=	16'h	c449;
63076	:douta	=	16'h	c449;
63077	:douta	=	16'h	c429;
63078	:douta	=	16'h	c429;
63079	:douta	=	16'h	c449;
63080	:douta	=	16'h	c428;
63081	:douta	=	16'h	c449;
63082	:douta	=	16'h	cc49;
63083	:douta	=	16'h	c449;
63084	:douta	=	16'h	c469;
63085	:douta	=	16'h	c469;
63086	:douta	=	16'h	c449;
63087	:douta	=	16'h	c449;
63088	:douta	=	16'h	c469;
63089	:douta	=	16'h	cc69;
63090	:douta	=	16'h	cc69;
63091	:douta	=	16'h	cc69;
63092	:douta	=	16'h	cc69;
63093	:douta	=	16'h	cc6a;
63094	:douta	=	16'h	cc49;
63095	:douta	=	16'h	cc69;
63096	:douta	=	16'h	cc69;
63097	:douta	=	16'h	cc6a;
63098	:douta	=	16'h	cc6a;
63099	:douta	=	16'h	cc6a;
63100	:douta	=	16'h	cc6a;
63101	:douta	=	16'h	cc6a;
63102	:douta	=	16'h	cc6a;
63103	:douta	=	16'h	cc69;
63104	:douta	=	16'h	cc8a;
63105	:douta	=	16'h	cc8a;
63106	:douta	=	16'h	cc89;
63107	:douta	=	16'h	cc69;
63108	:douta	=	16'h	cc69;
63109	:douta	=	16'h	cc69;
63110	:douta	=	16'h	cc69;
63111	:douta	=	16'h	cc89;
63112	:douta	=	16'h	cc69;
63113	:douta	=	16'h	cc89;
63114	:douta	=	16'h	cc69;
63115	:douta	=	16'h	cc89;
63116	:douta	=	16'h	cc69;
63117	:douta	=	16'h	cc6a;
63118	:douta	=	16'h	cc6a;
63119	:douta	=	16'h	cc69;
63120	:douta	=	16'h	cc6a;
63121	:douta	=	16'h	cc69;
63122	:douta	=	16'h	cc69;
63123	:douta	=	16'h	cc89;
63124	:douta	=	16'h	cc89;
63125	:douta	=	16'h	cc69;
63126	:douta	=	16'h	cc89;
63127	:douta	=	16'h	cc6a;
63128	:douta	=	16'h	cc6a;
63129	:douta	=	16'h	cc6a;
63130	:douta	=	16'h	cc89;
63131	:douta	=	16'h	cc89;
63132	:douta	=	16'h	cc6a;
63133	:douta	=	16'h	cc8a;
63134	:douta	=	16'h	cc8a;
63135	:douta	=	16'h	c469;
63136	:douta	=	16'h	cc6a;
63137	:douta	=	16'h	cc69;
63138	:douta	=	16'h	cc69;
63139	:douta	=	16'h	b5b5;
63140	:douta	=	16'h	e655;
63141	:douta	=	16'h	cc49;
63142	:douta	=	16'h	c469;
63143	:douta	=	16'h	c469;
63144	:douta	=	16'h	cc6a;
63145	:douta	=	16'h	cc69;
63146	:douta	=	16'h	cc6a;
63147	:douta	=	16'h	cc69;
63148	:douta	=	16'h	cc69;
63149	:douta	=	16'h	cc8a;
63150	:douta	=	16'h	cc6a;
63151	:douta	=	16'h	cc49;
63152	:douta	=	16'h	c449;
63153	:douta	=	16'h	c449;
63154	:douta	=	16'h	cc6a;
63155	:douta	=	16'h	c44a;
63156	:douta	=	16'h	cc69;
63157	:douta	=	16'h	cc69;
63158	:douta	=	16'h	c449;
63159	:douta	=	16'h	cc6a;
63160	:douta	=	16'h	c44a;
63161	:douta	=	16'h	c46a;
63162	:douta	=	16'h	c469;
63163	:douta	=	16'h	c46a;
63164	:douta	=	16'h	c449;
63165	:douta	=	16'h	c44a;
63166	:douta	=	16'h	c449;
63167	:douta	=	16'h	c449;
63168	:douta	=	16'h	c449;
63169	:douta	=	16'h	c449;
63170	:douta	=	16'h	c449;
63171	:douta	=	16'h	c429;
63172	:douta	=	16'h	c429;
63173	:douta	=	16'h	c44a;
63174	:douta	=	16'h	c429;
63175	:douta	=	16'h	c44a;
63176	:douta	=	16'h	c44a;
63177	:douta	=	16'h	c44a;
63178	:douta	=	16'h	c44a;
63179	:douta	=	16'h	c42a;
63180	:douta	=	16'h	c42a;
63181	:douta	=	16'h	bc2a;
63182	:douta	=	16'h	bc2a;
63183	:douta	=	16'h	c42a;
63184	:douta	=	16'h	bc09;
63185	:douta	=	16'h	bc2a;
63186	:douta	=	16'h	bc09;
63187	:douta	=	16'h	bc09;
63188	:douta	=	16'h	bc2a;
63189	:douta	=	16'h	bc09;
63190	:douta	=	16'h	bc2a;
63191	:douta	=	16'h	bc09;
63192	:douta	=	16'h	bc09;
63193	:douta	=	16'h	bc29;
63194	:douta	=	16'h	bc09;
63195	:douta	=	16'h	bc0a;
63196	:douta	=	16'h	bc09;
63197	:douta	=	16'h	bc09;
63198	:douta	=	16'h	bc09;
63199	:douta	=	16'h	bbe9;
63200	:douta	=	16'h	bc09;
63201	:douta	=	16'h	bbe9;
63202	:douta	=	16'h	bc09;
63203	:douta	=	16'h	bbe9;
63204	:douta	=	16'h	b3c9;
63205	:douta	=	16'h	b3e9;
63206	:douta	=	16'h	b3e9;
63207	:douta	=	16'h	b3e9;
63208	:douta	=	16'h	b3e9;
63209	:douta	=	16'h	b3e9;
63210	:douta	=	16'h	b3c9;
63211	:douta	=	16'h	b3ea;
63212	:douta	=	16'h	b3ca;
63213	:douta	=	16'h	b3c9;
63214	:douta	=	16'h	abc9;
63215	:douta	=	16'h	abc9;
63216	:douta	=	16'h	abc9;
63217	:douta	=	16'h	aba9;
63218	:douta	=	16'h	abc9;
63219	:douta	=	16'h	abca;
63220	:douta	=	16'h	aba9;
63221	:douta	=	16'h	aba9;
63222	:douta	=	16'h	aba9;
63223	:douta	=	16'h	aba9;
63224	:douta	=	16'h	aba9;
63225	:douta	=	16'h	ab89;
63226	:douta	=	16'h	aba9;
63227	:douta	=	16'h	a389;
63228	:douta	=	16'h	a389;
63229	:douta	=	16'h	ab89;
63230	:douta	=	16'h	a369;
63231	:douta	=	16'h	a389;
63232	:douta	=	16'h	4229;
63233	:douta	=	16'h	2924;
63234	:douta	=	16'h	3145;
63235	:douta	=	16'h	3125;
63236	:douta	=	16'h	3124;
63237	:douta	=	16'h	3124;
63238	:douta	=	16'h	3124;
63239	:douta	=	16'h	2924;
63240	:douta	=	16'h	2904;
63241	:douta	=	16'h	2904;
63242	:douta	=	16'h	2904;
63243	:douta	=	16'h	2904;
63244	:douta	=	16'h	28e4;
63245	:douta	=	16'h	28e3;
63246	:douta	=	16'h	2104;
63247	:douta	=	16'h	2103;
63248	:douta	=	16'h	2904;
63249	:douta	=	16'h	2924;
63250	:douta	=	16'h	20a2;
63251	:douta	=	16'h	20e3;
63252	:douta	=	16'h	28e3;
63253	:douta	=	16'h	28e3;
63254	:douta	=	16'h	28e3;
63255	:douta	=	16'h	2903;
63256	:douta	=	16'h	28e3;
63257	:douta	=	16'h	2903;
63258	:douta	=	16'h	28e3;
63259	:douta	=	16'h	28e3;
63260	:douta	=	16'h	3103;
63261	:douta	=	16'h	3923;
63262	:douta	=	16'h	3123;
63263	:douta	=	16'h	3923;
63264	:douta	=	16'h	3923;
63265	:douta	=	16'h	3944;
63266	:douta	=	16'h	4144;
63267	:douta	=	16'h	4143;
63268	:douta	=	16'h	4984;
63269	:douta	=	16'h	4984;
63270	:douta	=	16'h	49a5;
63271	:douta	=	16'h	4a4a;
63272	:douta	=	16'h	2105;
63273	:douta	=	16'h	3924;
63274	:douta	=	16'h	61e4;
63275	:douta	=	16'h	59e4;
63276	:douta	=	16'h	59e4;
63277	:douta	=	16'h	6205;
63278	:douta	=	16'h	6225;
63279	:douta	=	16'h	6a25;
63280	:douta	=	16'h	6a45;
63281	:douta	=	16'h	6a45;
63282	:douta	=	16'h	6a25;
63283	:douta	=	16'h	7224;
63284	:douta	=	16'h	72a8;
63285	:douta	=	16'h	b572;
63286	:douta	=	16'h	7a44;
63287	:douta	=	16'h	7a85;
63288	:douta	=	16'h	82a5;
63289	:douta	=	16'h	82a5;
63290	:douta	=	16'h	82a6;
63291	:douta	=	16'h	82c6;
63292	:douta	=	16'h	82c6;
63293	:douta	=	16'h	8ac7;
63294	:douta	=	16'h	8ac7;
63295	:douta	=	16'h	8ae7;
63296	:douta	=	16'h	8b07;
63297	:douta	=	16'h	8ae7;
63298	:douta	=	16'h	9307;
63299	:douta	=	16'h	9327;
63300	:douta	=	16'h	9327;
63301	:douta	=	16'h	9328;
63302	:douta	=	16'h	9327;
63303	:douta	=	16'h	9b47;
63304	:douta	=	16'h	9b47;
63305	:douta	=	16'h	9b68;
63306	:douta	=	16'h	9b68;
63307	:douta	=	16'h	9b68;
63308	:douta	=	16'h	a368;
63309	:douta	=	16'h	9b67;
63310	:douta	=	16'h	a388;
63311	:douta	=	16'h	a387;
63312	:douta	=	16'h	a388;
63313	:douta	=	16'h	ab87;
63314	:douta	=	16'h	aba8;
63315	:douta	=	16'h	b3c8;
63316	:douta	=	16'h	b3e8;
63317	:douta	=	16'h	b408;
63318	:douta	=	16'h	b408;
63319	:douta	=	16'h	b408;
63320	:douta	=	16'h	b3e8;
63321	:douta	=	16'h	bc09;
63322	:douta	=	16'h	bc09;
63323	:douta	=	16'h	bc09;
63324	:douta	=	16'h	bc09;
63325	:douta	=	16'h	bc09;
63326	:douta	=	16'h	bc29;
63327	:douta	=	16'h	bc29;
63328	:douta	=	16'h	bc49;
63329	:douta	=	16'h	bc49;
63330	:douta	=	16'h	c449;
63331	:douta	=	16'h	c449;
63332	:douta	=	16'h	c449;
63333	:douta	=	16'h	c449;
63334	:douta	=	16'h	c449;
63335	:douta	=	16'h	c449;
63336	:douta	=	16'h	c469;
63337	:douta	=	16'h	c469;
63338	:douta	=	16'h	c449;
63339	:douta	=	16'h	c469;
63340	:douta	=	16'h	c46a;
63341	:douta	=	16'h	c46a;
63342	:douta	=	16'h	c469;
63343	:douta	=	16'h	cc8a;
63344	:douta	=	16'h	cc6a;
63345	:douta	=	16'h	cc6a;
63346	:douta	=	16'h	c469;
63347	:douta	=	16'h	cc6a;
63348	:douta	=	16'h	cc6a;
63349	:douta	=	16'h	c469;
63350	:douta	=	16'h	cc6a;
63351	:douta	=	16'h	cc69;
63352	:douta	=	16'h	cc6a;
63353	:douta	=	16'h	cc8a;
63354	:douta	=	16'h	cc8a;
63355	:douta	=	16'h	cc69;
63356	:douta	=	16'h	cc6a;
63357	:douta	=	16'h	cc6a;
63358	:douta	=	16'h	cc6a;
63359	:douta	=	16'h	cc6a;
63360	:douta	=	16'h	cc8a;
63361	:douta	=	16'h	cc8a;
63362	:douta	=	16'h	cc89;
63363	:douta	=	16'h	cc69;
63364	:douta	=	16'h	cc69;
63365	:douta	=	16'h	cc89;
63366	:douta	=	16'h	cc69;
63367	:douta	=	16'h	cc89;
63368	:douta	=	16'h	cc69;
63369	:douta	=	16'h	cc69;
63370	:douta	=	16'h	cc69;
63371	:douta	=	16'h	cc69;
63372	:douta	=	16'h	cc69;
63373	:douta	=	16'h	cc69;
63374	:douta	=	16'h	cc69;
63375	:douta	=	16'h	cc69;
63376	:douta	=	16'h	cc69;
63377	:douta	=	16'h	cc69;
63378	:douta	=	16'h	cc69;
63379	:douta	=	16'h	cc69;
63380	:douta	=	16'h	c489;
63381	:douta	=	16'h	cc69;
63382	:douta	=	16'h	cc6a;
63383	:douta	=	16'h	cc6a;
63384	:douta	=	16'h	cc69;
63385	:douta	=	16'h	cc69;
63386	:douta	=	16'h	cc6a;
63387	:douta	=	16'h	cc69;
63388	:douta	=	16'h	cc6a;
63389	:douta	=	16'h	cc6a;
63390	:douta	=	16'h	cc8a;
63391	:douta	=	16'h	cc6a;
63392	:douta	=	16'h	cc6a;
63393	:douta	=	16'h	cc6a;
63394	:douta	=	16'h	cc6a;
63395	:douta	=	16'h	b5d5;
63396	:douta	=	16'h	e654;
63397	:douta	=	16'h	cc49;
63398	:douta	=	16'h	cc6a;
63399	:douta	=	16'h	cc6a;
63400	:douta	=	16'h	c469;
63401	:douta	=	16'h	cc69;
63402	:douta	=	16'h	cc69;
63403	:douta	=	16'h	cc69;
63404	:douta	=	16'h	cc69;
63405	:douta	=	16'h	cc6a;
63406	:douta	=	16'h	cc69;
63407	:douta	=	16'h	cc69;
63408	:douta	=	16'h	cc49;
63409	:douta	=	16'h	cc6a;
63410	:douta	=	16'h	c44a;
63411	:douta	=	16'h	c46a;
63412	:douta	=	16'h	cc69;
63413	:douta	=	16'h	cc69;
63414	:douta	=	16'h	c46a;
63415	:douta	=	16'h	c469;
63416	:douta	=	16'h	c46a;
63417	:douta	=	16'h	c449;
63418	:douta	=	16'h	c449;
63419	:douta	=	16'h	c449;
63420	:douta	=	16'h	c46a;
63421	:douta	=	16'h	c469;
63422	:douta	=	16'h	c44a;
63423	:douta	=	16'h	c469;
63424	:douta	=	16'h	c469;
63425	:douta	=	16'h	c44a;
63426	:douta	=	16'h	c44a;
63427	:douta	=	16'h	c44a;
63428	:douta	=	16'h	c44a;
63429	:douta	=	16'h	c44a;
63430	:douta	=	16'h	c42a;
63431	:douta	=	16'h	c44a;
63432	:douta	=	16'h	c42a;
63433	:douta	=	16'h	c44a;
63434	:douta	=	16'h	bc2a;
63435	:douta	=	16'h	c44a;
63436	:douta	=	16'h	c42a;
63437	:douta	=	16'h	c42a;
63438	:douta	=	16'h	bc2a;
63439	:douta	=	16'h	bc2a;
63440	:douta	=	16'h	bc2a;
63441	:douta	=	16'h	bc2a;
63442	:douta	=	16'h	bc29;
63443	:douta	=	16'h	bc2a;
63444	:douta	=	16'h	bc2a;
63445	:douta	=	16'h	bc09;
63446	:douta	=	16'h	bc0a;
63447	:douta	=	16'h	bc0a;
63448	:douta	=	16'h	bc0a;
63449	:douta	=	16'h	bc09;
63450	:douta	=	16'h	bc0a;
63451	:douta	=	16'h	bc09;
63452	:douta	=	16'h	bc09;
63453	:douta	=	16'h	bc09;
63454	:douta	=	16'h	bc09;
63455	:douta	=	16'h	bbe9;
63456	:douta	=	16'h	bbe9;
63457	:douta	=	16'h	bc09;
63458	:douta	=	16'h	b3e9;
63459	:douta	=	16'h	bbe9;
63460	:douta	=	16'h	bbe9;
63461	:douta	=	16'h	b3e9;
63462	:douta	=	16'h	b3e9;
63463	:douta	=	16'h	b3e9;
63464	:douta	=	16'h	b3e9;
63465	:douta	=	16'h	b3ca;
63466	:douta	=	16'h	b3ca;
63467	:douta	=	16'h	b3c9;
63468	:douta	=	16'h	b3c9;
63469	:douta	=	16'h	b3c9;
63470	:douta	=	16'h	b3e9;
63471	:douta	=	16'h	abc9;
63472	:douta	=	16'h	abc9;
63473	:douta	=	16'h	aba9;
63474	:douta	=	16'h	aba9;
63475	:douta	=	16'h	aba9;
63476	:douta	=	16'h	aba9;
63477	:douta	=	16'h	aba9;
63478	:douta	=	16'h	aba9;
63479	:douta	=	16'h	aba9;
63480	:douta	=	16'h	aba9;
63481	:douta	=	16'h	aba9;
63482	:douta	=	16'h	a389;
63483	:douta	=	16'h	a389;
63484	:douta	=	16'h	a389;
63485	:douta	=	16'h	a389;
63486	:douta	=	16'h	a369;
63487	:douta	=	16'h	a389;
63488	:douta	=	16'h	2124;
63489	:douta	=	16'h	2924;
63490	:douta	=	16'h	3145;
63491	:douta	=	16'h	3125;
63492	:douta	=	16'h	2924;
63493	:douta	=	16'h	3145;
63494	:douta	=	16'h	3124;
63495	:douta	=	16'h	2904;
63496	:douta	=	16'h	2924;
63497	:douta	=	16'h	2904;
63498	:douta	=	16'h	2904;
63499	:douta	=	16'h	2904;
63500	:douta	=	16'h	2904;
63501	:douta	=	16'h	20e3;
63502	:douta	=	16'h	2104;
63503	:douta	=	16'h	2104;
63504	:douta	=	16'h	28e3;
63505	:douta	=	16'h	2904;
63506	:douta	=	16'h	20c3;
63507	:douta	=	16'h	20c3;
63508	:douta	=	16'h	20e3;
63509	:douta	=	16'h	28e3;
63510	:douta	=	16'h	28e3;
63511	:douta	=	16'h	2903;
63512	:douta	=	16'h	2903;
63513	:douta	=	16'h	3103;
63514	:douta	=	16'h	3103;
63515	:douta	=	16'h	3103;
63516	:douta	=	16'h	3103;
63517	:douta	=	16'h	3123;
63518	:douta	=	16'h	3123;
63519	:douta	=	16'h	3923;
63520	:douta	=	16'h	3923;
63521	:douta	=	16'h	3944;
63522	:douta	=	16'h	4144;
63523	:douta	=	16'h	4143;
63524	:douta	=	16'h	4984;
63525	:douta	=	16'h	4984;
63526	:douta	=	16'h	4185;
63527	:douta	=	16'h	4229;
63528	:douta	=	16'h	18e5;
63529	:douta	=	16'h	4145;
63530	:douta	=	16'h	6205;
63531	:douta	=	16'h	59e4;
63532	:douta	=	16'h	6205;
63533	:douta	=	16'h	6205;
63534	:douta	=	16'h	6205;
63535	:douta	=	16'h	6205;
63536	:douta	=	16'h	6a25;
63537	:douta	=	16'h	6a45;
63538	:douta	=	16'h	6a25;
63539	:douta	=	16'h	7224;
63540	:douta	=	16'h	72ea;
63541	:douta	=	16'h	ad10;
63542	:douta	=	16'h	8285;
63543	:douta	=	16'h	8285;
63544	:douta	=	16'h	7a85;
63545	:douta	=	16'h	82a6;
63546	:douta	=	16'h	82c6;
63547	:douta	=	16'h	82c6;
63548	:douta	=	16'h	82c6;
63549	:douta	=	16'h	8ae7;
63550	:douta	=	16'h	8ac7;
63551	:douta	=	16'h	8ac6;
63552	:douta	=	16'h	8b07;
63553	:douta	=	16'h	8b07;
63554	:douta	=	16'h	9307;
63555	:douta	=	16'h	9307;
63556	:douta	=	16'h	9307;
63557	:douta	=	16'h	9b28;
63558	:douta	=	16'h	9327;
63559	:douta	=	16'h	9b47;
63560	:douta	=	16'h	9b68;
63561	:douta	=	16'h	9b68;
63562	:douta	=	16'h	9b68;
63563	:douta	=	16'h	9b68;
63564	:douta	=	16'h	9b68;
63565	:douta	=	16'h	9b67;
63566	:douta	=	16'h	a368;
63567	:douta	=	16'h	a388;
63568	:douta	=	16'h	a388;
63569	:douta	=	16'h	aba8;
63570	:douta	=	16'h	abc8;
63571	:douta	=	16'h	b3e8;
63572	:douta	=	16'h	b3e8;
63573	:douta	=	16'h	b3e8;
63574	:douta	=	16'h	bc08;
63575	:douta	=	16'h	b3e8;
63576	:douta	=	16'h	bc29;
63577	:douta	=	16'h	bc08;
63578	:douta	=	16'h	bc09;
63579	:douta	=	16'h	bc09;
63580	:douta	=	16'h	bc09;
63581	:douta	=	16'h	bc09;
63582	:douta	=	16'h	bc09;
63583	:douta	=	16'h	bc29;
63584	:douta	=	16'h	bc49;
63585	:douta	=	16'h	bc49;
63586	:douta	=	16'h	c449;
63587	:douta	=	16'h	bc29;
63588	:douta	=	16'h	bc49;
63589	:douta	=	16'h	c449;
63590	:douta	=	16'h	c449;
63591	:douta	=	16'h	c449;
63592	:douta	=	16'h	c469;
63593	:douta	=	16'h	c469;
63594	:douta	=	16'h	c46a;
63595	:douta	=	16'h	c46a;
63596	:douta	=	16'h	cc6a;
63597	:douta	=	16'h	c46a;
63598	:douta	=	16'h	c469;
63599	:douta	=	16'h	c469;
63600	:douta	=	16'h	c469;
63601	:douta	=	16'h	cc6a;
63602	:douta	=	16'h	c469;
63603	:douta	=	16'h	cc6a;
63604	:douta	=	16'h	cc6a;
63605	:douta	=	16'h	cc6a;
63606	:douta	=	16'h	cc6a;
63607	:douta	=	16'h	cc69;
63608	:douta	=	16'h	cc8a;
63609	:douta	=	16'h	cc8a;
63610	:douta	=	16'h	cc8a;
63611	:douta	=	16'h	cc8a;
63612	:douta	=	16'h	cc69;
63613	:douta	=	16'h	cc6a;
63614	:douta	=	16'h	cc6a;
63615	:douta	=	16'h	cc6a;
63616	:douta	=	16'h	cc6a;
63617	:douta	=	16'h	cc6a;
63618	:douta	=	16'h	cc8a;
63619	:douta	=	16'h	cc6a;
63620	:douta	=	16'h	cc69;
63621	:douta	=	16'h	cc8a;
63622	:douta	=	16'h	cc6a;
63623	:douta	=	16'h	cc69;
63624	:douta	=	16'h	cc69;
63625	:douta	=	16'h	cc69;
63626	:douta	=	16'h	cc69;
63627	:douta	=	16'h	cc89;
63628	:douta	=	16'h	cc89;
63629	:douta	=	16'h	cc89;
63630	:douta	=	16'h	cc69;
63631	:douta	=	16'h	cc69;
63632	:douta	=	16'h	c468;
63633	:douta	=	16'h	cc69;
63634	:douta	=	16'h	cc89;
63635	:douta	=	16'h	cc89;
63636	:douta	=	16'h	cc69;
63637	:douta	=	16'h	c469;
63638	:douta	=	16'h	cc8a;
63639	:douta	=	16'h	cc6a;
63640	:douta	=	16'h	cc6a;
63641	:douta	=	16'h	cc6a;
63642	:douta	=	16'h	cc6a;
63643	:douta	=	16'h	cc6a;
63644	:douta	=	16'h	cc6a;
63645	:douta	=	16'h	cc6a;
63646	:douta	=	16'h	cc6a;
63647	:douta	=	16'h	cc6a;
63648	:douta	=	16'h	cc6a;
63649	:douta	=	16'h	cc6a;
63650	:douta	=	16'h	cc6a;
63651	:douta	=	16'h	b5d5;
63652	:douta	=	16'h	e634;
63653	:douta	=	16'h	cc69;
63654	:douta	=	16'h	c469;
63655	:douta	=	16'h	cc6a;
63656	:douta	=	16'h	cc6a;
63657	:douta	=	16'h	c469;
63658	:douta	=	16'h	cc6a;
63659	:douta	=	16'h	cc6a;
63660	:douta	=	16'h	cc69;
63661	:douta	=	16'h	cc69;
63662	:douta	=	16'h	cc69;
63663	:douta	=	16'h	cc69;
63664	:douta	=	16'h	cc69;
63665	:douta	=	16'h	cc49;
63666	:douta	=	16'h	cc6a;
63667	:douta	=	16'h	c449;
63668	:douta	=	16'h	c449;
63669	:douta	=	16'h	c449;
63670	:douta	=	16'h	c46a;
63671	:douta	=	16'h	c46a;
63672	:douta	=	16'h	c44a;
63673	:douta	=	16'h	c449;
63674	:douta	=	16'h	c46a;
63675	:douta	=	16'h	c469;
63676	:douta	=	16'h	c469;
63677	:douta	=	16'h	c469;
63678	:douta	=	16'h	c44a;
63679	:douta	=	16'h	c44a;
63680	:douta	=	16'h	c44a;
63681	:douta	=	16'h	c44a;
63682	:douta	=	16'h	c44a;
63683	:douta	=	16'h	c44a;
63684	:douta	=	16'h	c429;
63685	:douta	=	16'h	c429;
63686	:douta	=	16'h	c44a;
63687	:douta	=	16'h	c44a;
63688	:douta	=	16'h	c42a;
63689	:douta	=	16'h	c44a;
63690	:douta	=	16'h	c44a;
63691	:douta	=	16'h	c44a;
63692	:douta	=	16'h	c44a;
63693	:douta	=	16'h	bc2a;
63694	:douta	=	16'h	c42a;
63695	:douta	=	16'h	bc2a;
63696	:douta	=	16'h	c44a;
63697	:douta	=	16'h	bc2a;
63698	:douta	=	16'h	bc2a;
63699	:douta	=	16'h	bc2a;
63700	:douta	=	16'h	bc2a;
63701	:douta	=	16'h	bc0a;
63702	:douta	=	16'h	bc0a;
63703	:douta	=	16'h	bc0a;
63704	:douta	=	16'h	bc0a;
63705	:douta	=	16'h	bc09;
63706	:douta	=	16'h	bc09;
63707	:douta	=	16'h	bc09;
63708	:douta	=	16'h	bc09;
63709	:douta	=	16'h	bbe9;
63710	:douta	=	16'h	bc09;
63711	:douta	=	16'h	bc09;
63712	:douta	=	16'h	b3e9;
63713	:douta	=	16'h	bbe9;
63714	:douta	=	16'h	b3e9;
63715	:douta	=	16'h	bbe9;
63716	:douta	=	16'h	b3e9;
63717	:douta	=	16'h	b3e9;
63718	:douta	=	16'h	b3e9;
63719	:douta	=	16'h	b3e9;
63720	:douta	=	16'h	b3c9;
63721	:douta	=	16'h	b3e9;
63722	:douta	=	16'h	abc9;
63723	:douta	=	16'h	b3c9;
63724	:douta	=	16'h	b3ca;
63725	:douta	=	16'h	b3c9;
63726	:douta	=	16'h	abc9;
63727	:douta	=	16'h	b3e9;
63728	:douta	=	16'h	abc9;
63729	:douta	=	16'h	abca;
63730	:douta	=	16'h	abca;
63731	:douta	=	16'h	aba9;
63732	:douta	=	16'h	aba9;
63733	:douta	=	16'h	aba9;
63734	:douta	=	16'h	aba9;
63735	:douta	=	16'h	aba9;
63736	:douta	=	16'h	aba9;
63737	:douta	=	16'h	aba9;
63738	:douta	=	16'h	aba9;
63739	:douta	=	16'h	a389;
63740	:douta	=	16'h	aba9;
63741	:douta	=	16'h	a369;
63742	:douta	=	16'h	a389;
63743	:douta	=	16'h	a389;
63744	:douta	=	16'h	2082;
63745	:douta	=	16'h	2945;
63746	:douta	=	16'h	3145;
63747	:douta	=	16'h	2924;
63748	:douta	=	16'h	2924;
63749	:douta	=	16'h	2924;
63750	:douta	=	16'h	2904;
63751	:douta	=	16'h	2924;
63752	:douta	=	16'h	2904;
63753	:douta	=	16'h	2924;
63754	:douta	=	16'h	2904;
63755	:douta	=	16'h	2924;
63756	:douta	=	16'h	2904;
63757	:douta	=	16'h	2904;
63758	:douta	=	16'h	2104;
63759	:douta	=	16'h	2104;
63760	:douta	=	16'h	2104;
63761	:douta	=	16'h	28e3;
63762	:douta	=	16'h	20e3;
63763	:douta	=	16'h	20e3;
63764	:douta	=	16'h	20c3;
63765	:douta	=	16'h	28e3;
63766	:douta	=	16'h	2903;
63767	:douta	=	16'h	2903;
63768	:douta	=	16'h	2903;
63769	:douta	=	16'h	2904;
63770	:douta	=	16'h	3104;
63771	:douta	=	16'h	3104;
63772	:douta	=	16'h	3103;
63773	:douta	=	16'h	3123;
63774	:douta	=	16'h	3123;
63775	:douta	=	16'h	3923;
63776	:douta	=	16'h	3923;
63777	:douta	=	16'h	3923;
63778	:douta	=	16'h	4144;
63779	:douta	=	16'h	4123;
63780	:douta	=	16'h	4964;
63781	:douta	=	16'h	4984;
63782	:douta	=	16'h	49c6;
63783	:douta	=	16'h	39a8;
63784	:douta	=	16'h	10a4;
63785	:douta	=	16'h	51a5;
63786	:douta	=	16'h	59c5;
63787	:douta	=	16'h	59e5;
63788	:douta	=	16'h	59e5;
63789	:douta	=	16'h	6205;
63790	:douta	=	16'h	6205;
63791	:douta	=	16'h	6a25;
63792	:douta	=	16'h	7266;
63793	:douta	=	16'h	6a45;
63794	:douta	=	16'h	7266;
63795	:douta	=	16'h	7245;
63796	:douta	=	16'h	7bae;
63797	:douta	=	16'h	9c2d;
63798	:douta	=	16'h	7a85;
63799	:douta	=	16'h	7a85;
63800	:douta	=	16'h	7aa5;
63801	:douta	=	16'h	82a6;
63802	:douta	=	16'h	82c6;
63803	:douta	=	16'h	82c6;
63804	:douta	=	16'h	8ac6;
63805	:douta	=	16'h	82c6;
63806	:douta	=	16'h	8ac7;
63807	:douta	=	16'h	8ae7;
63808	:douta	=	16'h	8ae7;
63809	:douta	=	16'h	8ae6;
63810	:douta	=	16'h	9307;
63811	:douta	=	16'h	8b07;
63812	:douta	=	16'h	9327;
63813	:douta	=	16'h	9328;
63814	:douta	=	16'h	9b48;
63815	:douta	=	16'h	9b48;
63816	:douta	=	16'h	9b48;
63817	:douta	=	16'h	9b68;
63818	:douta	=	16'h	9b68;
63819	:douta	=	16'h	9b68;
63820	:douta	=	16'h	a368;
63821	:douta	=	16'h	a368;
63822	:douta	=	16'h	a388;
63823	:douta	=	16'h	a388;
63824	:douta	=	16'h	ab88;
63825	:douta	=	16'h	aba8;
63826	:douta	=	16'h	abc8;
63827	:douta	=	16'h	b3e8;
63828	:douta	=	16'h	b3e9;
63829	:douta	=	16'h	b3e9;
63830	:douta	=	16'h	bc08;
63831	:douta	=	16'h	bc08;
63832	:douta	=	16'h	bc29;
63833	:douta	=	16'h	bc29;
63834	:douta	=	16'h	bc29;
63835	:douta	=	16'h	bc29;
63836	:douta	=	16'h	bc29;
63837	:douta	=	16'h	bc29;
63838	:douta	=	16'h	bc29;
63839	:douta	=	16'h	bc29;
63840	:douta	=	16'h	bc29;
63841	:douta	=	16'h	bc29;
63842	:douta	=	16'h	bc29;
63843	:douta	=	16'h	c449;
63844	:douta	=	16'h	c449;
63845	:douta	=	16'h	c449;
63846	:douta	=	16'h	c449;
63847	:douta	=	16'h	c449;
63848	:douta	=	16'h	c469;
63849	:douta	=	16'h	c469;
63850	:douta	=	16'h	c469;
63851	:douta	=	16'h	c46a;
63852	:douta	=	16'h	c46a;
63853	:douta	=	16'h	c46a;
63854	:douta	=	16'h	c46a;
63855	:douta	=	16'h	c469;
63856	:douta	=	16'h	cc6a;
63857	:douta	=	16'h	cc6a;
63858	:douta	=	16'h	c469;
63859	:douta	=	16'h	c469;
63860	:douta	=	16'h	cc8a;
63861	:douta	=	16'h	cc6a;
63862	:douta	=	16'h	cc6a;
63863	:douta	=	16'h	cc6a;
63864	:douta	=	16'h	cc8a;
63865	:douta	=	16'h	cc6a;
63866	:douta	=	16'h	cc6a;
63867	:douta	=	16'h	cc8a;
63868	:douta	=	16'h	cc8a;
63869	:douta	=	16'h	c469;
63870	:douta	=	16'h	cc8a;
63871	:douta	=	16'h	cc6a;
63872	:douta	=	16'h	cc8a;
63873	:douta	=	16'h	cc8a;
63874	:douta	=	16'h	cc6a;
63875	:douta	=	16'h	cc6a;
63876	:douta	=	16'h	cc6a;
63877	:douta	=	16'h	cc6a;
63878	:douta	=	16'h	cc69;
63879	:douta	=	16'h	cc6a;
63880	:douta	=	16'h	cc6a;
63881	:douta	=	16'h	cc6a;
63882	:douta	=	16'h	cc89;
63883	:douta	=	16'h	cc69;
63884	:douta	=	16'h	cc69;
63885	:douta	=	16'h	cc69;
63886	:douta	=	16'h	cc69;
63887	:douta	=	16'h	cc6a;
63888	:douta	=	16'h	cc69;
63889	:douta	=	16'h	cc69;
63890	:douta	=	16'h	cc69;
63891	:douta	=	16'h	cc69;
63892	:douta	=	16'h	cc69;
63893	:douta	=	16'h	cc8a;
63894	:douta	=	16'h	cc6a;
63895	:douta	=	16'h	cc6a;
63896	:douta	=	16'h	cc6a;
63897	:douta	=	16'h	cc6a;
63898	:douta	=	16'h	cc6a;
63899	:douta	=	16'h	cc69;
63900	:douta	=	16'h	c469;
63901	:douta	=	16'h	c469;
63902	:douta	=	16'h	cc6a;
63903	:douta	=	16'h	cc8a;
63904	:douta	=	16'h	cc6a;
63905	:douta	=	16'h	cc69;
63906	:douta	=	16'h	cc69;
63907	:douta	=	16'h	bdd5;
63908	:douta	=	16'h	e634;
63909	:douta	=	16'h	c449;
63910	:douta	=	16'h	cc6a;
63911	:douta	=	16'h	cc6a;
63912	:douta	=	16'h	c46a;
63913	:douta	=	16'h	cc6a;
63914	:douta	=	16'h	c46a;
63915	:douta	=	16'h	c46a;
63916	:douta	=	16'h	cc6a;
63917	:douta	=	16'h	cc69;
63918	:douta	=	16'h	cc69;
63919	:douta	=	16'h	cc69;
63920	:douta	=	16'h	cc69;
63921	:douta	=	16'h	cc69;
63922	:douta	=	16'h	cc6a;
63923	:douta	=	16'h	cc6a;
63924	:douta	=	16'h	c46a;
63925	:douta	=	16'h	c46a;
63926	:douta	=	16'h	c46a;
63927	:douta	=	16'h	c469;
63928	:douta	=	16'h	c46a;
63929	:douta	=	16'h	c46a;
63930	:douta	=	16'h	c449;
63931	:douta	=	16'h	c44a;
63932	:douta	=	16'h	c44a;
63933	:douta	=	16'h	c44a;
63934	:douta	=	16'h	c44a;
63935	:douta	=	16'h	c44a;
63936	:douta	=	16'h	c429;
63937	:douta	=	16'h	c44a;
63938	:douta	=	16'h	c44a;
63939	:douta	=	16'h	c429;
63940	:douta	=	16'h	c44a;
63941	:douta	=	16'h	c429;
63942	:douta	=	16'h	c44a;
63943	:douta	=	16'h	c44a;
63944	:douta	=	16'h	c44a;
63945	:douta	=	16'h	c44a;
63946	:douta	=	16'h	c44a;
63947	:douta	=	16'h	c42a;
63948	:douta	=	16'h	bc2a;
63949	:douta	=	16'h	bc2a;
63950	:douta	=	16'h	bc2a;
63951	:douta	=	16'h	bc2a;
63952	:douta	=	16'h	bc2a;
63953	:douta	=	16'h	bc29;
63954	:douta	=	16'h	bc2a;
63955	:douta	=	16'h	bc2a;
63956	:douta	=	16'h	bc0a;
63957	:douta	=	16'h	bc0a;
63958	:douta	=	16'h	bc2a;
63959	:douta	=	16'h	bc0a;
63960	:douta	=	16'h	bc09;
63961	:douta	=	16'h	bc0a;
63962	:douta	=	16'h	bc09;
63963	:douta	=	16'h	bc09;
63964	:douta	=	16'h	bbe9;
63965	:douta	=	16'h	bc09;
63966	:douta	=	16'h	bc09;
63967	:douta	=	16'h	bc09;
63968	:douta	=	16'h	bc09;
63969	:douta	=	16'h	b3e9;
63970	:douta	=	16'h	bc09;
63971	:douta	=	16'h	b3e9;
63972	:douta	=	16'h	b3e9;
63973	:douta	=	16'h	b3e9;
63974	:douta	=	16'h	b3e9;
63975	:douta	=	16'h	b3e9;
63976	:douta	=	16'h	b3c9;
63977	:douta	=	16'h	b3ca;
63978	:douta	=	16'h	b3c9;
63979	:douta	=	16'h	b3ca;
63980	:douta	=	16'h	b3c9;
63981	:douta	=	16'h	aba9;
63982	:douta	=	16'h	abca;
63983	:douta	=	16'h	aba9;
63984	:douta	=	16'h	aba9;
63985	:douta	=	16'h	aba9;
63986	:douta	=	16'h	aba9;
63987	:douta	=	16'h	aba9;
63988	:douta	=	16'h	aba9;
63989	:douta	=	16'h	aba9;
63990	:douta	=	16'h	aba9;
63991	:douta	=	16'h	ab89;
63992	:douta	=	16'h	a389;
63993	:douta	=	16'h	ab89;
63994	:douta	=	16'h	a389;
63995	:douta	=	16'h	a389;
63996	:douta	=	16'h	a369;
63997	:douta	=	16'h	ab89;
63998	:douta	=	16'h	a369;
63999	:douta	=	16'h	a389;
64000	:douta	=	16'h	2904;
64001	:douta	=	16'h	3145;
64002	:douta	=	16'h	3125;
64003	:douta	=	16'h	2924;
64004	:douta	=	16'h	2904;
64005	:douta	=	16'h	2924;
64006	:douta	=	16'h	2924;
64007	:douta	=	16'h	2924;
64008	:douta	=	16'h	28e3;
64009	:douta	=	16'h	2924;
64010	:douta	=	16'h	2924;
64011	:douta	=	16'h	2904;
64012	:douta	=	16'h	2904;
64013	:douta	=	16'h	2104;
64014	:douta	=	16'h	2103;
64015	:douta	=	16'h	2104;
64016	:douta	=	16'h	2924;
64017	:douta	=	16'h	20e3;
64018	:douta	=	16'h	20e3;
64019	:douta	=	16'h	20e3;
64020	:douta	=	16'h	20c3;
64021	:douta	=	16'h	2903;
64022	:douta	=	16'h	2903;
64023	:douta	=	16'h	28e3;
64024	:douta	=	16'h	2903;
64025	:douta	=	16'h	2903;
64026	:douta	=	16'h	3124;
64027	:douta	=	16'h	3104;
64028	:douta	=	16'h	3103;
64029	:douta	=	16'h	3123;
64030	:douta	=	16'h	3923;
64031	:douta	=	16'h	3923;
64032	:douta	=	16'h	3923;
64033	:douta	=	16'h	3944;
64034	:douta	=	16'h	4124;
64035	:douta	=	16'h	4144;
64036	:douta	=	16'h	4964;
64037	:douta	=	16'h	4984;
64038	:douta	=	16'h	49c7;
64039	:douta	=	16'h	3187;
64040	:douta	=	16'h	0884;
64041	:douta	=	16'h	59c4;
64042	:douta	=	16'h	59c4;
64043	:douta	=	16'h	59e4;
64044	:douta	=	16'h	6205;
64045	:douta	=	16'h	6205;
64046	:douta	=	16'h	6a25;
64047	:douta	=	16'h	6a25;
64048	:douta	=	16'h	7266;
64049	:douta	=	16'h	7265;
64050	:douta	=	16'h	7265;
64051	:douta	=	16'h	7285;
64052	:douta	=	16'h	8430;
64053	:douta	=	16'h	93eb;
64054	:douta	=	16'h	7aa6;
64055	:douta	=	16'h	7aa5;
64056	:douta	=	16'h	82a6;
64057	:douta	=	16'h	82a6;
64058	:douta	=	16'h	82c6;
64059	:douta	=	16'h	82c6;
64060	:douta	=	16'h	82c6;
64061	:douta	=	16'h	8ac7;
64062	:douta	=	16'h	8ac7;
64063	:douta	=	16'h	8ae7;
64064	:douta	=	16'h	8b07;
64065	:douta	=	16'h	8b07;
64066	:douta	=	16'h	8b07;
64067	:douta	=	16'h	8b07;
64068	:douta	=	16'h	9327;
64069	:douta	=	16'h	9328;
64070	:douta	=	16'h	9b48;
64071	:douta	=	16'h	9b48;
64072	:douta	=	16'h	9b48;
64073	:douta	=	16'h	9b48;
64074	:douta	=	16'h	9b68;
64075	:douta	=	16'h	a388;
64076	:douta	=	16'h	a368;
64077	:douta	=	16'h	a368;
64078	:douta	=	16'h	a388;
64079	:douta	=	16'h	a388;
64080	:douta	=	16'h	a388;
64081	:douta	=	16'h	aba8;
64082	:douta	=	16'h	abc8;
64083	:douta	=	16'h	b3c8;
64084	:douta	=	16'h	b3e9;
64085	:douta	=	16'h	b3e9;
64086	:douta	=	16'h	bc09;
64087	:douta	=	16'h	b409;
64088	:douta	=	16'h	bc09;
64089	:douta	=	16'h	bc29;
64090	:douta	=	16'h	bc09;
64091	:douta	=	16'h	bc2a;
64092	:douta	=	16'h	bc2a;
64093	:douta	=	16'h	bc2a;
64094	:douta	=	16'h	bc29;
64095	:douta	=	16'h	bc29;
64096	:douta	=	16'h	c44a;
64097	:douta	=	16'h	bc29;
64098	:douta	=	16'h	bc49;
64099	:douta	=	16'h	bc49;
64100	:douta	=	16'h	bc49;
64101	:douta	=	16'h	c449;
64102	:douta	=	16'h	c449;
64103	:douta	=	16'h	c469;
64104	:douta	=	16'h	c469;
64105	:douta	=	16'h	c449;
64106	:douta	=	16'h	c469;
64107	:douta	=	16'h	c46a;
64108	:douta	=	16'h	c48a;
64109	:douta	=	16'h	c46a;
64110	:douta	=	16'h	cc8a;
64111	:douta	=	16'h	c469;
64112	:douta	=	16'h	c469;
64113	:douta	=	16'h	cc6a;
64114	:douta	=	16'h	c469;
64115	:douta	=	16'h	c48a;
64116	:douta	=	16'h	c48a;
64117	:douta	=	16'h	cc6a;
64118	:douta	=	16'h	cc6a;
64119	:douta	=	16'h	c469;
64120	:douta	=	16'h	cc6a;
64121	:douta	=	16'h	cc6a;
64122	:douta	=	16'h	cc6a;
64123	:douta	=	16'h	c469;
64124	:douta	=	16'h	cc6a;
64125	:douta	=	16'h	cc6a;
64126	:douta	=	16'h	cc8a;
64127	:douta	=	16'h	cc8a;
64128	:douta	=	16'h	cc6a;
64129	:douta	=	16'h	cc6a;
64130	:douta	=	16'h	cc6a;
64131	:douta	=	16'h	cc6a;
64132	:douta	=	16'h	cc6a;
64133	:douta	=	16'h	cc6a;
64134	:douta	=	16'h	cc6a;
64135	:douta	=	16'h	cc6a;
64136	:douta	=	16'h	c469;
64137	:douta	=	16'h	cc6a;
64138	:douta	=	16'h	cc6a;
64139	:douta	=	16'h	cc69;
64140	:douta	=	16'h	cc69;
64141	:douta	=	16'h	cc69;
64142	:douta	=	16'h	cc69;
64143	:douta	=	16'h	cc69;
64144	:douta	=	16'h	cc6a;
64145	:douta	=	16'h	cc6a;
64146	:douta	=	16'h	cc69;
64147	:douta	=	16'h	cc89;
64148	:douta	=	16'h	cc69;
64149	:douta	=	16'h	cc6a;
64150	:douta	=	16'h	cc6a;
64151	:douta	=	16'h	cc6a;
64152	:douta	=	16'h	cc6a;
64153	:douta	=	16'h	cc6a;
64154	:douta	=	16'h	cc6a;
64155	:douta	=	16'h	cc6a;
64156	:douta	=	16'h	c469;
64157	:douta	=	16'h	cc6a;
64158	:douta	=	16'h	cc6a;
64159	:douta	=	16'h	cc6a;
64160	:douta	=	16'h	cc6a;
64161	:douta	=	16'h	cc69;
64162	:douta	=	16'h	cc6a;
64163	:douta	=	16'h	bdd6;
64164	:douta	=	16'h	e634;
64165	:douta	=	16'h	c44a;
64166	:douta	=	16'h	cc6a;
64167	:douta	=	16'h	cc6a;
64168	:douta	=	16'h	cc6a;
64169	:douta	=	16'h	cc6a;
64170	:douta	=	16'h	c46a;
64171	:douta	=	16'h	c46a;
64172	:douta	=	16'h	cc6a;
64173	:douta	=	16'h	cc6a;
64174	:douta	=	16'h	cc69;
64175	:douta	=	16'h	cc69;
64176	:douta	=	16'h	cc69;
64177	:douta	=	16'h	c449;
64178	:douta	=	16'h	c44a;
64179	:douta	=	16'h	c44a;
64180	:douta	=	16'h	c469;
64181	:douta	=	16'h	c469;
64182	:douta	=	16'h	c46a;
64183	:douta	=	16'h	c449;
64184	:douta	=	16'h	c46a;
64185	:douta	=	16'h	c449;
64186	:douta	=	16'h	c449;
64187	:douta	=	16'h	c44a;
64188	:douta	=	16'h	c44a;
64189	:douta	=	16'h	c44a;
64190	:douta	=	16'h	c44a;
64191	:douta	=	16'h	c44a;
64192	:douta	=	16'h	c44a;
64193	:douta	=	16'h	c44a;
64194	:douta	=	16'h	c44a;
64195	:douta	=	16'h	c429;
64196	:douta	=	16'h	c44a;
64197	:douta	=	16'h	bc29;
64198	:douta	=	16'h	c44a;
64199	:douta	=	16'h	bc2a;
64200	:douta	=	16'h	c42a;
64201	:douta	=	16'h	c42a;
64202	:douta	=	16'h	c42a;
64203	:douta	=	16'h	bc2a;
64204	:douta	=	16'h	bc2a;
64205	:douta	=	16'h	bc0a;
64206	:douta	=	16'h	bc2a;
64207	:douta	=	16'h	bc2a;
64208	:douta	=	16'h	bc2a;
64209	:douta	=	16'h	c42a;
64210	:douta	=	16'h	bc2a;
64211	:douta	=	16'h	bc2a;
64212	:douta	=	16'h	bc0a;
64213	:douta	=	16'h	bc2a;
64214	:douta	=	16'h	bc2a;
64215	:douta	=	16'h	bc2a;
64216	:douta	=	16'h	bc0a;
64217	:douta	=	16'h	bc0a;
64218	:douta	=	16'h	bc09;
64219	:douta	=	16'h	bc0a;
64220	:douta	=	16'h	bc09;
64221	:douta	=	16'h	bbe9;
64222	:douta	=	16'h	bbe9;
64223	:douta	=	16'h	bbe9;
64224	:douta	=	16'h	bbe9;
64225	:douta	=	16'h	b3ea;
64226	:douta	=	16'h	b3e9;
64227	:douta	=	16'h	b3ea;
64228	:douta	=	16'h	b3e9;
64229	:douta	=	16'h	b3e9;
64230	:douta	=	16'h	b3e9;
64231	:douta	=	16'h	b3e9;
64232	:douta	=	16'h	b3e9;
64233	:douta	=	16'h	b3ca;
64234	:douta	=	16'h	b3ca;
64235	:douta	=	16'h	abc9;
64236	:douta	=	16'h	abc9;
64237	:douta	=	16'h	abca;
64238	:douta	=	16'h	abca;
64239	:douta	=	16'h	aba9;
64240	:douta	=	16'h	aba9;
64241	:douta	=	16'h	aba9;
64242	:douta	=	16'h	aba9;
64243	:douta	=	16'h	aba9;
64244	:douta	=	16'h	aba9;
64245	:douta	=	16'h	ab89;
64246	:douta	=	16'h	ab89;
64247	:douta	=	16'h	abaa;
64248	:douta	=	16'h	a389;
64249	:douta	=	16'h	abaa;
64250	:douta	=	16'h	a369;
64251	:douta	=	16'h	a369;
64252	:douta	=	16'h	a389;
64253	:douta	=	16'h	ab8a;
64254	:douta	=	16'h	a38a;
64255	:douta	=	16'h	a389;
64256	:douta	=	16'h	3146;
64257	:douta	=	16'h	3145;
64258	:douta	=	16'h	2945;
64259	:douta	=	16'h	2924;
64260	:douta	=	16'h	2904;
64261	:douta	=	16'h	2904;
64262	:douta	=	16'h	2924;
64263	:douta	=	16'h	2904;
64264	:douta	=	16'h	2904;
64265	:douta	=	16'h	2924;
64266	:douta	=	16'h	2924;
64267	:douta	=	16'h	2904;
64268	:douta	=	16'h	2904;
64269	:douta	=	16'h	2924;
64270	:douta	=	16'h	2104;
64271	:douta	=	16'h	2104;
64272	:douta	=	16'h	2924;
64273	:douta	=	16'h	20c3;
64274	:douta	=	16'h	20e3;
64275	:douta	=	16'h	20e3;
64276	:douta	=	16'h	20e3;
64277	:douta	=	16'h	28e3;
64278	:douta	=	16'h	2903;
64279	:douta	=	16'h	28e3;
64280	:douta	=	16'h	2904;
64281	:douta	=	16'h	2903;
64282	:douta	=	16'h	3123;
64283	:douta	=	16'h	3103;
64284	:douta	=	16'h	3124;
64285	:douta	=	16'h	3123;
64286	:douta	=	16'h	3923;
64287	:douta	=	16'h	3923;
64288	:douta	=	16'h	3944;
64289	:douta	=	16'h	3923;
64290	:douta	=	16'h	4164;
64291	:douta	=	16'h	4164;
64292	:douta	=	16'h	4964;
64293	:douta	=	16'h	4163;
64294	:douta	=	16'h	526a;
64295	:douta	=	16'h	1906;
64296	:douta	=	16'h	0884;
64297	:douta	=	16'h	59c4;
64298	:douta	=	16'h	59c4;
64299	:douta	=	16'h	59e5;
64300	:douta	=	16'h	59e4;
64301	:douta	=	16'h	6205;
64302	:douta	=	16'h	6a25;
64303	:douta	=	16'h	6a25;
64304	:douta	=	16'h	7246;
64305	:douta	=	16'h	7265;
64306	:douta	=	16'h	7286;
64307	:douta	=	16'h	7ae9;
64308	:douta	=	16'h	9d14;
64309	:douta	=	16'h	82e7;
64310	:douta	=	16'h	7a86;
64311	:douta	=	16'h	82a6;
64312	:douta	=	16'h	82a6;
64313	:douta	=	16'h	82c6;
64314	:douta	=	16'h	82c6;
64315	:douta	=	16'h	82c6;
64316	:douta	=	16'h	8ae6;
64317	:douta	=	16'h	8ac7;
64318	:douta	=	16'h	8ae7;
64319	:douta	=	16'h	8ae7;
64320	:douta	=	16'h	8b07;
64321	:douta	=	16'h	8b07;
64322	:douta	=	16'h	8ae7;
64323	:douta	=	16'h	8b07;
64324	:douta	=	16'h	9327;
64325	:douta	=	16'h	9328;
64326	:douta	=	16'h	9b48;
64327	:douta	=	16'h	9b28;
64328	:douta	=	16'h	9b48;
64329	:douta	=	16'h	9b48;
64330	:douta	=	16'h	a388;
64331	:douta	=	16'h	a388;
64332	:douta	=	16'h	9b67;
64333	:douta	=	16'h	a368;
64334	:douta	=	16'h	a388;
64335	:douta	=	16'h	a387;
64336	:douta	=	16'h	ab88;
64337	:douta	=	16'h	aba8;
64338	:douta	=	16'h	abc8;
64339	:douta	=	16'h	b3e8;
64340	:douta	=	16'h	b3e9;
64341	:douta	=	16'h	b409;
64342	:douta	=	16'h	b3e9;
64343	:douta	=	16'h	b409;
64344	:douta	=	16'h	bc09;
64345	:douta	=	16'h	bc2a;
64346	:douta	=	16'h	bc2a;
64347	:douta	=	16'h	bc2a;
64348	:douta	=	16'h	bc2a;
64349	:douta	=	16'h	c42a;
64350	:douta	=	16'h	c42a;
64351	:douta	=	16'h	bc29;
64352	:douta	=	16'h	bc29;
64353	:douta	=	16'h	bc29;
64354	:douta	=	16'h	bc29;
64355	:douta	=	16'h	c449;
64356	:douta	=	16'h	c449;
64357	:douta	=	16'h	c449;
64358	:douta	=	16'h	c449;
64359	:douta	=	16'h	c469;
64360	:douta	=	16'h	c449;
64361	:douta	=	16'h	c44a;
64362	:douta	=	16'h	c46a;
64363	:douta	=	16'h	c46a;
64364	:douta	=	16'h	cc6a;
64365	:douta	=	16'h	cc8b;
64366	:douta	=	16'h	c46a;
64367	:douta	=	16'h	c46a;
64368	:douta	=	16'h	c46a;
64369	:douta	=	16'h	c46a;
64370	:douta	=	16'h	c46a;
64371	:douta	=	16'h	c48a;
64372	:douta	=	16'h	c48a;
64373	:douta	=	16'h	cc8a;
64374	:douta	=	16'h	c469;
64375	:douta	=	16'h	cc89;
64376	:douta	=	16'h	cc8a;
64377	:douta	=	16'h	cc6a;
64378	:douta	=	16'h	cc6a;
64379	:douta	=	16'h	cc6a;
64380	:douta	=	16'h	cc6a;
64381	:douta	=	16'h	cc6a;
64382	:douta	=	16'h	cc6a;
64383	:douta	=	16'h	c469;
64384	:douta	=	16'h	cc8a;
64385	:douta	=	16'h	cc6a;
64386	:douta	=	16'h	cc69;
64387	:douta	=	16'h	cc89;
64388	:douta	=	16'h	cc69;
64389	:douta	=	16'h	cc8a;
64390	:douta	=	16'h	c469;
64391	:douta	=	16'h	cc6a;
64392	:douta	=	16'h	cc6a;
64393	:douta	=	16'h	cc6a;
64394	:douta	=	16'h	cc69;
64395	:douta	=	16'h	cc6a;
64396	:douta	=	16'h	cc69;
64397	:douta	=	16'h	cc69;
64398	:douta	=	16'h	cc69;
64399	:douta	=	16'h	cc6a;
64400	:douta	=	16'h	cc69;
64401	:douta	=	16'h	cc6a;
64402	:douta	=	16'h	cc6a;
64403	:douta	=	16'h	cc6a;
64404	:douta	=	16'h	cc69;
64405	:douta	=	16'h	cc6a;
64406	:douta	=	16'h	cc69;
64407	:douta	=	16'h	cc6a;
64408	:douta	=	16'h	c469;
64409	:douta	=	16'h	cc69;
64410	:douta	=	16'h	cc69;
64411	:douta	=	16'h	cc6a;
64412	:douta	=	16'h	cc6a;
64413	:douta	=	16'h	cc8a;
64414	:douta	=	16'h	cc6a;
64415	:douta	=	16'h	cc8a;
64416	:douta	=	16'h	cc6a;
64417	:douta	=	16'h	cc69;
64418	:douta	=	16'h	c46a;
64419	:douta	=	16'h	bdd6;
64420	:douta	=	16'h	e634;
64421	:douta	=	16'h	cc49;
64422	:douta	=	16'h	cc6a;
64423	:douta	=	16'h	cc6a;
64424	:douta	=	16'h	c46a;
64425	:douta	=	16'h	c46a;
64426	:douta	=	16'h	c46a;
64427	:douta	=	16'h	c46a;
64428	:douta	=	16'h	c46a;
64429	:douta	=	16'h	c469;
64430	:douta	=	16'h	c469;
64431	:douta	=	16'h	c449;
64432	:douta	=	16'h	c449;
64433	:douta	=	16'h	c46a;
64434	:douta	=	16'h	c469;
64435	:douta	=	16'h	c44a;
64436	:douta	=	16'h	c469;
64437	:douta	=	16'h	c449;
64438	:douta	=	16'h	c469;
64439	:douta	=	16'h	c469;
64440	:douta	=	16'h	c469;
64441	:douta	=	16'h	c44a;
64442	:douta	=	16'h	c429;
64443	:douta	=	16'h	c44a;
64444	:douta	=	16'h	c44a;
64445	:douta	=	16'h	c44a;
64446	:douta	=	16'h	c44a;
64447	:douta	=	16'h	c44a;
64448	:douta	=	16'h	c44a;
64449	:douta	=	16'h	c44a;
64450	:douta	=	16'h	c44a;
64451	:douta	=	16'h	c44a;
64452	:douta	=	16'h	c429;
64453	:douta	=	16'h	c44a;
64454	:douta	=	16'h	bc2a;
64455	:douta	=	16'h	c44a;
64456	:douta	=	16'h	c42a;
64457	:douta	=	16'h	bc2a;
64458	:douta	=	16'h	c44a;
64459	:douta	=	16'h	bc2a;
64460	:douta	=	16'h	c42a;
64461	:douta	=	16'h	bc2a;
64462	:douta	=	16'h	bc2a;
64463	:douta	=	16'h	bc2a;
64464	:douta	=	16'h	bc2a;
64465	:douta	=	16'h	bc29;
64466	:douta	=	16'h	bc2a;
64467	:douta	=	16'h	bc2a;
64468	:douta	=	16'h	bc2a;
64469	:douta	=	16'h	bc0a;
64470	:douta	=	16'h	bc2a;
64471	:douta	=	16'h	bc09;
64472	:douta	=	16'h	bc09;
64473	:douta	=	16'h	bc09;
64474	:douta	=	16'h	bc09;
64475	:douta	=	16'h	bc09;
64476	:douta	=	16'h	bc09;
64477	:douta	=	16'h	bc09;
64478	:douta	=	16'h	bbe9;
64479	:douta	=	16'h	b3ea;
64480	:douta	=	16'h	b40a;
64481	:douta	=	16'h	b3e9;
64482	:douta	=	16'h	b3ea;
64483	:douta	=	16'h	b3e9;
64484	:douta	=	16'h	b3e9;
64485	:douta	=	16'h	b3e9;
64486	:douta	=	16'h	b3ea;
64487	:douta	=	16'h	b3ca;
64488	:douta	=	16'h	b3ca;
64489	:douta	=	16'h	b3ca;
64490	:douta	=	16'h	b3ca;
64491	:douta	=	16'h	b3e9;
64492	:douta	=	16'h	b3e9;
64493	:douta	=	16'h	abca;
64494	:douta	=	16'h	abca;
64495	:douta	=	16'h	aba9;
64496	:douta	=	16'h	aba9;
64497	:douta	=	16'h	aba9;
64498	:douta	=	16'h	aba9;
64499	:douta	=	16'h	aba9;
64500	:douta	=	16'h	aba9;
64501	:douta	=	16'h	abaa;
64502	:douta	=	16'h	abaa;
64503	:douta	=	16'h	a389;
64504	:douta	=	16'h	abaa;
64505	:douta	=	16'h	ab89;
64506	:douta	=	16'h	ab89;
64507	:douta	=	16'h	a369;
64508	:douta	=	16'h	ab89;
64509	:douta	=	16'h	a389;
64510	:douta	=	16'h	a369;
64511	:douta	=	16'h	a389;
64512	:douta	=	16'h	3145;
64513	:douta	=	16'h	3145;
64514	:douta	=	16'h	2925;
64515	:douta	=	16'h	2924;
64516	:douta	=	16'h	2904;
64517	:douta	=	16'h	2904;
64518	:douta	=	16'h	2904;
64519	:douta	=	16'h	2904;
64520	:douta	=	16'h	2904;
64521	:douta	=	16'h	3124;
64522	:douta	=	16'h	2924;
64523	:douta	=	16'h	2904;
64524	:douta	=	16'h	2904;
64525	:douta	=	16'h	20e4;
64526	:douta	=	16'h	2104;
64527	:douta	=	16'h	2104;
64528	:douta	=	16'h	2104;
64529	:douta	=	16'h	20c3;
64530	:douta	=	16'h	20e3;
64531	:douta	=	16'h	20e3;
64532	:douta	=	16'h	20e3;
64533	:douta	=	16'h	2924;
64534	:douta	=	16'h	2903;
64535	:douta	=	16'h	2903;
64536	:douta	=	16'h	28e3;
64537	:douta	=	16'h	3124;
64538	:douta	=	16'h	3103;
64539	:douta	=	16'h	3103;
64540	:douta	=	16'h	3123;
64541	:douta	=	16'h	3123;
64542	:douta	=	16'h	3924;
64543	:douta	=	16'h	3923;
64544	:douta	=	16'h	3944;
64545	:douta	=	16'h	3944;
64546	:douta	=	16'h	4964;
64547	:douta	=	16'h	4164;
64548	:douta	=	16'h	4985;
64549	:douta	=	16'h	4964;
64550	:douta	=	16'h	5aab;
64551	:douta	=	16'h	18e5;
64552	:douta	=	16'h	1084;
64553	:douta	=	16'h	59c4;
64554	:douta	=	16'h	51c4;
64555	:douta	=	16'h	6205;
64556	:douta	=	16'h	59e5;
64557	:douta	=	16'h	6205;
64558	:douta	=	16'h	6a25;
64559	:douta	=	16'h	6a45;
64560	:douta	=	16'h	7246;
64561	:douta	=	16'h	7266;
64562	:douta	=	16'h	7265;
64563	:douta	=	16'h	732b;
64564	:douta	=	16'h	a576;
64565	:douta	=	16'h	7a86;
64566	:douta	=	16'h	82c7;
64567	:douta	=	16'h	82a6;
64568	:douta	=	16'h	82a6;
64569	:douta	=	16'h	82c6;
64570	:douta	=	16'h	82c6;
64571	:douta	=	16'h	8ae7;
64572	:douta	=	16'h	8ae7;
64573	:douta	=	16'h	8ae7;
64574	:douta	=	16'h	8ac7;
64575	:douta	=	16'h	8b07;
64576	:douta	=	16'h	8b07;
64577	:douta	=	16'h	8b07;
64578	:douta	=	16'h	8b07;
64579	:douta	=	16'h	9308;
64580	:douta	=	16'h	9327;
64581	:douta	=	16'h	9328;
64582	:douta	=	16'h	9b48;
64583	:douta	=	16'h	9b48;
64584	:douta	=	16'h	9b48;
64585	:douta	=	16'h	9b48;
64586	:douta	=	16'h	a368;
64587	:douta	=	16'h	a388;
64588	:douta	=	16'h	9b67;
64589	:douta	=	16'h	a368;
64590	:douta	=	16'h	a388;
64591	:douta	=	16'h	a387;
64592	:douta	=	16'h	a387;
64593	:douta	=	16'h	aba8;
64594	:douta	=	16'h	abc8;
64595	:douta	=	16'h	b3c9;
64596	:douta	=	16'h	b409;
64597	:douta	=	16'h	b409;
64598	:douta	=	16'h	b409;
64599	:douta	=	16'h	b409;
64600	:douta	=	16'h	b409;
64601	:douta	=	16'h	bc2a;
64602	:douta	=	16'h	bc2a;
64603	:douta	=	16'h	c42a;
64604	:douta	=	16'h	c42a;
64605	:douta	=	16'h	c44a;
64606	:douta	=	16'h	bc2a;
64607	:douta	=	16'h	c44a;
64608	:douta	=	16'h	bc29;
64609	:douta	=	16'h	bc29;
64610	:douta	=	16'h	bc29;
64611	:douta	=	16'h	c44a;
64612	:douta	=	16'h	bc49;
64613	:douta	=	16'h	c44a;
64614	:douta	=	16'h	c44a;
64615	:douta	=	16'h	c469;
64616	:douta	=	16'h	c449;
64617	:douta	=	16'h	c44a;
64618	:douta	=	16'h	cc6a;
64619	:douta	=	16'h	c46a;
64620	:douta	=	16'h	cc6a;
64621	:douta	=	16'h	c46a;
64622	:douta	=	16'h	c46a;
64623	:douta	=	16'h	c46a;
64624	:douta	=	16'h	c46a;
64625	:douta	=	16'h	c46a;
64626	:douta	=	16'h	c46a;
64627	:douta	=	16'h	c48a;
64628	:douta	=	16'h	c48a;
64629	:douta	=	16'h	cc8a;
64630	:douta	=	16'h	cc6a;
64631	:douta	=	16'h	cc6a;
64632	:douta	=	16'h	cc8a;
64633	:douta	=	16'h	cc6a;
64634	:douta	=	16'h	cc6a;
64635	:douta	=	16'h	cc8a;
64636	:douta	=	16'h	cc8a;
64637	:douta	=	16'h	cc6a;
64638	:douta	=	16'h	cc6a;
64639	:douta	=	16'h	cc6a;
64640	:douta	=	16'h	cc6a;
64641	:douta	=	16'h	cc6a;
64642	:douta	=	16'h	cc69;
64643	:douta	=	16'h	c489;
64644	:douta	=	16'h	c489;
64645	:douta	=	16'h	cc6a;
64646	:douta	=	16'h	cc6a;
64647	:douta	=	16'h	cc6a;
64648	:douta	=	16'h	cc69;
64649	:douta	=	16'h	cc6a;
64650	:douta	=	16'h	cc69;
64651	:douta	=	16'h	cc69;
64652	:douta	=	16'h	cc49;
64653	:douta	=	16'h	cc6a;
64654	:douta	=	16'h	cc69;
64655	:douta	=	16'h	cc69;
64656	:douta	=	16'h	cc6a;
64657	:douta	=	16'h	cc6a;
64658	:douta	=	16'h	cc69;
64659	:douta	=	16'h	cc69;
64660	:douta	=	16'h	cc69;
64661	:douta	=	16'h	cc6a;
64662	:douta	=	16'h	cc6a;
64663	:douta	=	16'h	cc6a;
64664	:douta	=	16'h	c469;
64665	:douta	=	16'h	c469;
64666	:douta	=	16'h	cc6a;
64667	:douta	=	16'h	cc6a;
64668	:douta	=	16'h	cc8a;
64669	:douta	=	16'h	cc8a;
64670	:douta	=	16'h	c469;
64671	:douta	=	16'h	cc8a;
64672	:douta	=	16'h	cc6a;
64673	:douta	=	16'h	cc69;
64674	:douta	=	16'h	c46a;
64675	:douta	=	16'h	bdd6;
64676	:douta	=	16'h	de33;
64677	:douta	=	16'h	c449;
64678	:douta	=	16'h	c46a;
64679	:douta	=	16'h	c46a;
64680	:douta	=	16'h	c46a;
64681	:douta	=	16'h	c46a;
64682	:douta	=	16'h	c46a;
64683	:douta	=	16'h	c46a;
64684	:douta	=	16'h	c46a;
64685	:douta	=	16'h	c469;
64686	:douta	=	16'h	c469;
64687	:douta	=	16'h	c469;
64688	:douta	=	16'h	c469;
64689	:douta	=	16'h	c46a;
64690	:douta	=	16'h	c449;
64691	:douta	=	16'h	c449;
64692	:douta	=	16'h	c469;
64693	:douta	=	16'h	c46a;
64694	:douta	=	16'h	c46a;
64695	:douta	=	16'h	c469;
64696	:douta	=	16'h	c449;
64697	:douta	=	16'h	c44a;
64698	:douta	=	16'h	c44a;
64699	:douta	=	16'h	c44a;
64700	:douta	=	16'h	c44a;
64701	:douta	=	16'h	c44a;
64702	:douta	=	16'h	c44a;
64703	:douta	=	16'h	c44a;
64704	:douta	=	16'h	c44a;
64705	:douta	=	16'h	c44a;
64706	:douta	=	16'h	c44a;
64707	:douta	=	16'h	c429;
64708	:douta	=	16'h	c44a;
64709	:douta	=	16'h	c42a;
64710	:douta	=	16'h	c42a;
64711	:douta	=	16'h	c42a;
64712	:douta	=	16'h	bc2a;
64713	:douta	=	16'h	c42a;
64714	:douta	=	16'h	c44a;
64715	:douta	=	16'h	bc2a;
64716	:douta	=	16'h	bc2a;
64717	:douta	=	16'h	bc2a;
64718	:douta	=	16'h	bc2a;
64719	:douta	=	16'h	bc2a;
64720	:douta	=	16'h	bc2a;
64721	:douta	=	16'h	bc2a;
64722	:douta	=	16'h	bc0a;
64723	:douta	=	16'h	bc2a;
64724	:douta	=	16'h	bc0a;
64725	:douta	=	16'h	bc0a;
64726	:douta	=	16'h	bc0a;
64727	:douta	=	16'h	bc0a;
64728	:douta	=	16'h	bc0a;
64729	:douta	=	16'h	bc0a;
64730	:douta	=	16'h	bc0a;
64731	:douta	=	16'h	bc09;
64732	:douta	=	16'h	bc09;
64733	:douta	=	16'h	b3ea;
64734	:douta	=	16'h	b40a;
64735	:douta	=	16'h	b3ea;
64736	:douta	=	16'h	b3e9;
64737	:douta	=	16'h	b40a;
64738	:douta	=	16'h	b3e9;
64739	:douta	=	16'h	b3e9;
64740	:douta	=	16'h	b3ea;
64741	:douta	=	16'h	b3ea;
64742	:douta	=	16'h	b3ca;
64743	:douta	=	16'h	b3ca;
64744	:douta	=	16'h	b3ca;
64745	:douta	=	16'h	b3ca;
64746	:douta	=	16'h	b3c9;
64747	:douta	=	16'h	abc9;
64748	:douta	=	16'h	abc9;
64749	:douta	=	16'h	abca;
64750	:douta	=	16'h	abca;
64751	:douta	=	16'h	abca;
64752	:douta	=	16'h	aba9;
64753	:douta	=	16'h	aba9;
64754	:douta	=	16'h	aba9;
64755	:douta	=	16'h	aba9;
64756	:douta	=	16'h	ab89;
64757	:douta	=	16'h	abaa;
64758	:douta	=	16'h	ab89;
64759	:douta	=	16'h	a389;
64760	:douta	=	16'h	a389;
64761	:douta	=	16'h	ab89;
64762	:douta	=	16'h	a389;
64763	:douta	=	16'h	a369;
64764	:douta	=	16'h	a389;
64765	:douta	=	16'h	a369;
64766	:douta	=	16'h	ab89;
64767	:douta	=	16'h	a369;
64768	:douta	=	16'h	2945;
64769	:douta	=	16'h	3145;
64770	:douta	=	16'h	3145;
64771	:douta	=	16'h	2944;
64772	:douta	=	16'h	2924;
64773	:douta	=	16'h	2924;
64774	:douta	=	16'h	2904;
64775	:douta	=	16'h	28e3;
64776	:douta	=	16'h	2924;
64777	:douta	=	16'h	2904;
64778	:douta	=	16'h	2904;
64779	:douta	=	16'h	2904;
64780	:douta	=	16'h	2104;
64781	:douta	=	16'h	2104;
64782	:douta	=	16'h	2104;
64783	:douta	=	16'h	20e4;
64784	:douta	=	16'h	2104;
64785	:douta	=	16'h	20c3;
64786	:douta	=	16'h	20e3;
64787	:douta	=	16'h	20e3;
64788	:douta	=	16'h	20e3;
64789	:douta	=	16'h	28e3;
64790	:douta	=	16'h	2903;
64791	:douta	=	16'h	2903;
64792	:douta	=	16'h	2904;
64793	:douta	=	16'h	3104;
64794	:douta	=	16'h	3103;
64795	:douta	=	16'h	3124;
64796	:douta	=	16'h	3123;
64797	:douta	=	16'h	3944;
64798	:douta	=	16'h	3944;
64799	:douta	=	16'h	3944;
64800	:douta	=	16'h	3944;
64801	:douta	=	16'h	4164;
64802	:douta	=	16'h	4965;
64803	:douta	=	16'h	4964;
64804	:douta	=	16'h	4984;
64805	:douta	=	16'h	4965;
64806	:douta	=	16'h	5aab;
64807	:douta	=	16'h	10a3;
64808	:douta	=	16'h	18c4;
64809	:douta	=	16'h	59c4;
64810	:douta	=	16'h	59c4;
64811	:douta	=	16'h	59e5;
64812	:douta	=	16'h	59e4;
64813	:douta	=	16'h	6205;
64814	:douta	=	16'h	6a25;
64815	:douta	=	16'h	6a45;
64816	:douta	=	16'h	6a45;
64817	:douta	=	16'h	7266;
64818	:douta	=	16'h	7265;
64819	:douta	=	16'h	7bcf;
64820	:douta	=	16'h	b617;
64821	:douta	=	16'h	7245;
64822	:douta	=	16'h	7a86;
64823	:douta	=	16'h	82a6;
64824	:douta	=	16'h	82c7;
64825	:douta	=	16'h	82c7;
64826	:douta	=	16'h	82c6;
64827	:douta	=	16'h	8ae7;
64828	:douta	=	16'h	8ac6;
64829	:douta	=	16'h	8ae6;
64830	:douta	=	16'h	8ae7;
64831	:douta	=	16'h	8b07;
64832	:douta	=	16'h	8b07;
64833	:douta	=	16'h	8b07;
64834	:douta	=	16'h	8b07;
64835	:douta	=	16'h	9308;
64836	:douta	=	16'h	9328;
64837	:douta	=	16'h	9348;
64838	:douta	=	16'h	9b48;
64839	:douta	=	16'h	9b48;
64840	:douta	=	16'h	9b48;
64841	:douta	=	16'h	9b69;
64842	:douta	=	16'h	9b68;
64843	:douta	=	16'h	9b48;
64844	:douta	=	16'h	a388;
64845	:douta	=	16'h	a388;
64846	:douta	=	16'h	a368;
64847	:douta	=	16'h	a3a8;
64848	:douta	=	16'h	a3a8;
64849	:douta	=	16'h	aba8;
64850	:douta	=	16'h	aba8;
64851	:douta	=	16'h	b3e9;
64852	:douta	=	16'h	b3e9;
64853	:douta	=	16'h	b3e9;
64854	:douta	=	16'h	b409;
64855	:douta	=	16'h	bc09;
64856	:douta	=	16'h	b409;
64857	:douta	=	16'h	bc2a;
64858	:douta	=	16'h	bc2a;
64859	:douta	=	16'h	bc2a;
64860	:douta	=	16'h	c42a;
64861	:douta	=	16'h	bc2a;
64862	:douta	=	16'h	bc2a;
64863	:douta	=	16'h	bc49;
64864	:douta	=	16'h	c44a;
64865	:douta	=	16'h	bc29;
64866	:douta	=	16'h	c44a;
64867	:douta	=	16'h	c44a;
64868	:douta	=	16'h	c44a;
64869	:douta	=	16'h	c44a;
64870	:douta	=	16'h	c44a;
64871	:douta	=	16'h	c44a;
64872	:douta	=	16'h	c44a;
64873	:douta	=	16'h	c44a;
64874	:douta	=	16'h	c46a;
64875	:douta	=	16'h	c48a;
64876	:douta	=	16'h	c46a;
64877	:douta	=	16'h	c46a;
64878	:douta	=	16'h	c46a;
64879	:douta	=	16'h	c48a;
64880	:douta	=	16'h	c46a;
64881	:douta	=	16'h	c46a;
64882	:douta	=	16'h	c46a;
64883	:douta	=	16'h	cc6a;
64884	:douta	=	16'h	c48a;
64885	:douta	=	16'h	c48a;
64886	:douta	=	16'h	cc6a;
64887	:douta	=	16'h	cc8a;
64888	:douta	=	16'h	cc6a;
64889	:douta	=	16'h	cc6a;
64890	:douta	=	16'h	cc8a;
64891	:douta	=	16'h	cc6a;
64892	:douta	=	16'h	cc6a;
64893	:douta	=	16'h	cc6a;
64894	:douta	=	16'h	cc8a;
64895	:douta	=	16'h	cc8a;
64896	:douta	=	16'h	cc6a;
64897	:douta	=	16'h	cc6a;
64898	:douta	=	16'h	c469;
64899	:douta	=	16'h	c489;
64900	:douta	=	16'h	cc89;
64901	:douta	=	16'h	c469;
64902	:douta	=	16'h	cc6a;
64903	:douta	=	16'h	cc6a;
64904	:douta	=	16'h	cc6a;
64905	:douta	=	16'h	cc6a;
64906	:douta	=	16'h	cc69;
64907	:douta	=	16'h	cc6a;
64908	:douta	=	16'h	cc6a;
64909	:douta	=	16'h	cc69;
64910	:douta	=	16'h	cc6a;
64911	:douta	=	16'h	cc6a;
64912	:douta	=	16'h	cc6a;
64913	:douta	=	16'h	cc6a;
64914	:douta	=	16'h	cc6a;
64915	:douta	=	16'h	cc6a;
64916	:douta	=	16'h	cc69;
64917	:douta	=	16'h	cc6a;
64918	:douta	=	16'h	cc6a;
64919	:douta	=	16'h	cc6a;
64920	:douta	=	16'h	cc6a;
64921	:douta	=	16'h	cc6a;
64922	:douta	=	16'h	cc6a;
64923	:douta	=	16'h	cc6a;
64924	:douta	=	16'h	cc6a;
64925	:douta	=	16'h	cc6a;
64926	:douta	=	16'h	cc6a;
64927	:douta	=	16'h	cc6a;
64928	:douta	=	16'h	cc6a;
64929	:douta	=	16'h	cc69;
64930	:douta	=	16'h	c46a;
64931	:douta	=	16'h	bdf6;
64932	:douta	=	16'h	de13;
64933	:douta	=	16'h	cc69;
64934	:douta	=	16'h	cc6a;
64935	:douta	=	16'h	cc6a;
64936	:douta	=	16'h	cc6a;
64937	:douta	=	16'h	cc8a;
64938	:douta	=	16'h	c46a;
64939	:douta	=	16'h	c469;
64940	:douta	=	16'h	c46a;
64941	:douta	=	16'h	c469;
64942	:douta	=	16'h	c46a;
64943	:douta	=	16'h	c469;
64944	:douta	=	16'h	c469;
64945	:douta	=	16'h	c469;
64946	:douta	=	16'h	c469;
64947	:douta	=	16'h	c469;
64948	:douta	=	16'h	c469;
64949	:douta	=	16'h	c469;
64950	:douta	=	16'h	c469;
64951	:douta	=	16'h	c44a;
64952	:douta	=	16'h	c44a;
64953	:douta	=	16'h	c44a;
64954	:douta	=	16'h	c44a;
64955	:douta	=	16'h	c44a;
64956	:douta	=	16'h	c429;
64957	:douta	=	16'h	c429;
64958	:douta	=	16'h	bc29;
64959	:douta	=	16'h	c44a;
64960	:douta	=	16'h	bc29;
64961	:douta	=	16'h	c44a;
64962	:douta	=	16'h	c44a;
64963	:douta	=	16'h	c44a;
64964	:douta	=	16'h	c42a;
64965	:douta	=	16'h	c42a;
64966	:douta	=	16'h	bc2a;
64967	:douta	=	16'h	c42a;
64968	:douta	=	16'h	bc2a;
64969	:douta	=	16'h	c42a;
64970	:douta	=	16'h	bc2a;
64971	:douta	=	16'h	bc2a;
64972	:douta	=	16'h	bc2a;
64973	:douta	=	16'h	bc2a;
64974	:douta	=	16'h	bc2a;
64975	:douta	=	16'h	bc2a;
64976	:douta	=	16'h	bc0a;
64977	:douta	=	16'h	bc0a;
64978	:douta	=	16'h	bc0a;
64979	:douta	=	16'h	bc09;
64980	:douta	=	16'h	bc2a;
64981	:douta	=	16'h	bc0a;
64982	:douta	=	16'h	bc0a;
64983	:douta	=	16'h	bc09;
64984	:douta	=	16'h	bc0a;
64985	:douta	=	16'h	b3e9;
64986	:douta	=	16'h	b40a;
64987	:douta	=	16'h	bc0a;
64988	:douta	=	16'h	b409;
64989	:douta	=	16'h	b40a;
64990	:douta	=	16'h	b3e9;
64991	:douta	=	16'h	b40a;
64992	:douta	=	16'h	b3e9;
64993	:douta	=	16'h	b3ea;
64994	:douta	=	16'h	b3ea;
64995	:douta	=	16'h	b3e9;
64996	:douta	=	16'h	b3e9;
64997	:douta	=	16'h	b3ca;
64998	:douta	=	16'h	b3e9;
64999	:douta	=	16'h	b3ca;
65000	:douta	=	16'h	abc9;
65001	:douta	=	16'h	b3e9;
65002	:douta	=	16'h	abc9;
65003	:douta	=	16'h	abc9;
65004	:douta	=	16'h	abc9;
65005	:douta	=	16'h	abc9;
65006	:douta	=	16'h	aba9;
65007	:douta	=	16'h	abc9;
65008	:douta	=	16'h	aba9;
65009	:douta	=	16'h	b3ca;
65010	:douta	=	16'h	ab8a;
65011	:douta	=	16'h	abaa;
65012	:douta	=	16'h	a389;
65013	:douta	=	16'h	abaa;
65014	:douta	=	16'h	abaa;
65015	:douta	=	16'h	a389;
65016	:douta	=	16'h	ab89;
65017	:douta	=	16'h	abaa;
65018	:douta	=	16'h	a389;
65019	:douta	=	16'h	a38a;
65020	:douta	=	16'h	a389;
65021	:douta	=	16'h	a369;
65022	:douta	=	16'h	a369;
65023	:douta	=	16'h	a38a;
65024	:douta	=	16'h	2945;
65025	:douta	=	16'h	3145;
65026	:douta	=	16'h	2924;
65027	:douta	=	16'h	2924;
65028	:douta	=	16'h	2104;
65029	:douta	=	16'h	2924;
65030	:douta	=	16'h	2924;
65031	:douta	=	16'h	2104;
65032	:douta	=	16'h	2104;
65033	:douta	=	16'h	3124;
65034	:douta	=	16'h	2904;
65035	:douta	=	16'h	2104;
65036	:douta	=	16'h	2104;
65037	:douta	=	16'h	20e4;
65038	:douta	=	16'h	2104;
65039	:douta	=	16'h	2104;
65040	:douta	=	16'h	20e3;
65041	:douta	=	16'h	20e3;
65042	:douta	=	16'h	20c3;
65043	:douta	=	16'h	28e3;
65044	:douta	=	16'h	28e3;
65045	:douta	=	16'h	2903;
65046	:douta	=	16'h	2903;
65047	:douta	=	16'h	2904;
65048	:douta	=	16'h	3104;
65049	:douta	=	16'h	3104;
65050	:douta	=	16'h	3124;
65051	:douta	=	16'h	3124;
65052	:douta	=	16'h	3124;
65053	:douta	=	16'h	3944;
65054	:douta	=	16'h	3944;
65055	:douta	=	16'h	3944;
65056	:douta	=	16'h	3944;
65057	:douta	=	16'h	4164;
65058	:douta	=	16'h	4164;
65059	:douta	=	16'h	4985;
65060	:douta	=	16'h	4985;
65061	:douta	=	16'h	4985;
65062	:douta	=	16'h	5aaa;
65063	:douta	=	16'h	0884;
65064	:douta	=	16'h	28e3;
65065	:douta	=	16'h	59c5;
65066	:douta	=	16'h	59c4;
65067	:douta	=	16'h	59e4;
65068	:douta	=	16'h	6205;
65069	:douta	=	16'h	6205;
65070	:douta	=	16'h	6a25;
65071	:douta	=	16'h	6a45;
65072	:douta	=	16'h	7266;
65073	:douta	=	16'h	7267;
65074	:douta	=	16'h	7266;
65075	:douta	=	16'h	8430;
65076	:douta	=	16'h	be17;
65077	:douta	=	16'h	7a44;
65078	:douta	=	16'h	82a6;
65079	:douta	=	16'h	82c7;
65080	:douta	=	16'h	82c7;
65081	:douta	=	16'h	82c7;
65082	:douta	=	16'h	82c6;
65083	:douta	=	16'h	8ae6;
65084	:douta	=	16'h	8ae7;
65085	:douta	=	16'h	8ae7;
65086	:douta	=	16'h	8ae7;
65087	:douta	=	16'h	8b07;
65088	:douta	=	16'h	8b07;
65089	:douta	=	16'h	8b07;
65090	:douta	=	16'h	8b07;
65091	:douta	=	16'h	8b07;
65092	:douta	=	16'h	9308;
65093	:douta	=	16'h	9348;
65094	:douta	=	16'h	9348;
65095	:douta	=	16'h	9b48;
65096	:douta	=	16'h	9b48;
65097	:douta	=	16'h	9b68;
65098	:douta	=	16'h	9b68;
65099	:douta	=	16'h	9b68;
65100	:douta	=	16'h	9b68;
65101	:douta	=	16'h	a368;
65102	:douta	=	16'h	a388;
65103	:douta	=	16'h	a388;
65104	:douta	=	16'h	a388;
65105	:douta	=	16'h	aba8;
65106	:douta	=	16'h	abc8;
65107	:douta	=	16'h	abe9;
65108	:douta	=	16'h	b3e9;
65109	:douta	=	16'h	b3e9;
65110	:douta	=	16'h	b409;
65111	:douta	=	16'h	b409;
65112	:douta	=	16'h	b409;
65113	:douta	=	16'h	bc0a;
65114	:douta	=	16'h	bc2a;
65115	:douta	=	16'h	bc2a;
65116	:douta	=	16'h	bc2a;
65117	:douta	=	16'h	bc2a;
65118	:douta	=	16'h	c42a;
65119	:douta	=	16'h	c44a;
65120	:douta	=	16'h	bc49;
65121	:douta	=	16'h	bc29;
65122	:douta	=	16'h	bc29;
65123	:douta	=	16'h	bc29;
65124	:douta	=	16'h	c44a;
65125	:douta	=	16'h	c44a;
65126	:douta	=	16'h	bc49;
65127	:douta	=	16'h	c44a;
65128	:douta	=	16'h	c44a;
65129	:douta	=	16'h	c46a;
65130	:douta	=	16'h	c46a;
65131	:douta	=	16'h	c46a;
65132	:douta	=	16'h	c46a;
65133	:douta	=	16'h	c46a;
65134	:douta	=	16'h	c44a;
65135	:douta	=	16'h	cc6a;
65136	:douta	=	16'h	c46a;
65137	:douta	=	16'h	c48a;
65138	:douta	=	16'h	c46a;
65139	:douta	=	16'h	cc6a;
65140	:douta	=	16'h	c48a;
65141	:douta	=	16'h	cc8a;
65142	:douta	=	16'h	cc6a;
65143	:douta	=	16'h	c46a;
65144	:douta	=	16'h	c469;
65145	:douta	=	16'h	c489;
65146	:douta	=	16'h	c48a;
65147	:douta	=	16'h	c48a;
65148	:douta	=	16'h	c48a;
65149	:douta	=	16'h	cc6a;
65150	:douta	=	16'h	cc8a;
65151	:douta	=	16'h	cc6a;
65152	:douta	=	16'h	cc6a;
65153	:douta	=	16'h	cc6a;
65154	:douta	=	16'h	c469;
65155	:douta	=	16'h	c489;
65156	:douta	=	16'h	cc69;
65157	:douta	=	16'h	c469;
65158	:douta	=	16'h	c469;
65159	:douta	=	16'h	cc6a;
65160	:douta	=	16'h	c469;
65161	:douta	=	16'h	cc6a;
65162	:douta	=	16'h	cc6a;
65163	:douta	=	16'h	c469;
65164	:douta	=	16'h	cc6a;
65165	:douta	=	16'h	cc6a;
65166	:douta	=	16'h	cc69;
65167	:douta	=	16'h	cc69;
65168	:douta	=	16'h	c469;
65169	:douta	=	16'h	cc6a;
65170	:douta	=	16'h	cc69;
65171	:douta	=	16'h	cc6a;
65172	:douta	=	16'h	cc6a;
65173	:douta	=	16'h	cc69;
65174	:douta	=	16'h	cc6a;
65175	:douta	=	16'h	cc6a;
65176	:douta	=	16'h	cc6a;
65177	:douta	=	16'h	cc6a;
65178	:douta	=	16'h	c46a;
65179	:douta	=	16'h	cc6a;
65180	:douta	=	16'h	cc6a;
65181	:douta	=	16'h	cc6a;
65182	:douta	=	16'h	cc6a;
65183	:douta	=	16'h	cc6a;
65184	:douta	=	16'h	cc6a;
65185	:douta	=	16'h	cc69;
65186	:douta	=	16'h	c46a;
65187	:douta	=	16'h	be16;
65188	:douta	=	16'h	de34;
65189	:douta	=	16'h	cc69;
65190	:douta	=	16'h	c46a;
65191	:douta	=	16'h	cc6a;
65192	:douta	=	16'h	c46a;
65193	:douta	=	16'h	c46a;
65194	:douta	=	16'h	c46a;
65195	:douta	=	16'h	c46a;
65196	:douta	=	16'h	c469;
65197	:douta	=	16'h	c46a;
65198	:douta	=	16'h	c46a;
65199	:douta	=	16'h	c46a;
65200	:douta	=	16'h	c469;
65201	:douta	=	16'h	c46a;
65202	:douta	=	16'h	c46a;
65203	:douta	=	16'h	c46a;
65204	:douta	=	16'h	c469;
65205	:douta	=	16'h	c469;
65206	:douta	=	16'h	c44a;
65207	:douta	=	16'h	c44a;
65208	:douta	=	16'h	c44a;
65209	:douta	=	16'h	c44a;
65210	:douta	=	16'h	c429;
65211	:douta	=	16'h	c44a;
65212	:douta	=	16'h	bc29;
65213	:douta	=	16'h	bc29;
65214	:douta	=	16'h	c44a;
65215	:douta	=	16'h	c44a;
65216	:douta	=	16'h	bc29;
65217	:douta	=	16'h	c42a;
65218	:douta	=	16'h	c42a;
65219	:douta	=	16'h	c42a;
65220	:douta	=	16'h	c42a;
65221	:douta	=	16'h	bc2a;
65222	:douta	=	16'h	c42a;
65223	:douta	=	16'h	c42a;
65224	:douta	=	16'h	bc2a;
65225	:douta	=	16'h	bc2a;
65226	:douta	=	16'h	bc2a;
65227	:douta	=	16'h	c42a;
65228	:douta	=	16'h	bc2a;
65229	:douta	=	16'h	bc2a;
65230	:douta	=	16'h	bc2a;
65231	:douta	=	16'h	bc2a;
65232	:douta	=	16'h	bc0a;
65233	:douta	=	16'h	bc2a;
65234	:douta	=	16'h	bc0a;
65235	:douta	=	16'h	bc0a;
65236	:douta	=	16'h	bc0a;
65237	:douta	=	16'h	bc0a;
65238	:douta	=	16'h	bc0a;
65239	:douta	=	16'h	bc0a;
65240	:douta	=	16'h	bc0a;
65241	:douta	=	16'h	bc0a;
65242	:douta	=	16'h	b40a;
65243	:douta	=	16'h	b40a;
65244	:douta	=	16'h	b3ea;
65245	:douta	=	16'h	b3ea;
65246	:douta	=	16'h	b40a;
65247	:douta	=	16'h	b40a;
65248	:douta	=	16'h	b40a;
65249	:douta	=	16'h	b3e9;
65250	:douta	=	16'h	b3ea;
65251	:douta	=	16'h	b40a;
65252	:douta	=	16'h	abc9;
65253	:douta	=	16'h	b3ea;
65254	:douta	=	16'h	b3ea;
65255	:douta	=	16'h	b3e9;
65256	:douta	=	16'h	b3e9;
65257	:douta	=	16'h	abc9;
65258	:douta	=	16'h	abc9;
65259	:douta	=	16'h	abc9;
65260	:douta	=	16'h	abc9;
65261	:douta	=	16'h	aba9;
65262	:douta	=	16'h	aba9;
65263	:douta	=	16'h	aba9;
65264	:douta	=	16'h	aba9;
65265	:douta	=	16'h	abaa;
65266	:douta	=	16'h	abaa;
65267	:douta	=	16'h	abaa;
65268	:douta	=	16'h	a389;
65269	:douta	=	16'h	a38a;
65270	:douta	=	16'h	a389;
65271	:douta	=	16'h	ab89;
65272	:douta	=	16'h	abaa;
65273	:douta	=	16'h	a389;
65274	:douta	=	16'h	a389;
65275	:douta	=	16'h	a389;
65276	:douta	=	16'h	a389;
65277	:douta	=	16'h	ab8a;
65278	:douta	=	16'h	a389;
65279	:douta	=	16'h	a38a;
65280	:douta	=	16'h	3145;
65281	:douta	=	16'h	2925;
65282	:douta	=	16'h	2924;
65283	:douta	=	16'h	2924;
65284	:douta	=	16'h	2924;
65285	:douta	=	16'h	2924;
65286	:douta	=	16'h	2104;
65287	:douta	=	16'h	2104;
65288	:douta	=	16'h	2104;
65289	:douta	=	16'h	2104;
65290	:douta	=	16'h	2924;
65291	:douta	=	16'h	2104;
65292	:douta	=	16'h	2104;
65293	:douta	=	16'h	2104;
65294	:douta	=	16'h	2924;
65295	:douta	=	16'h	2924;
65296	:douta	=	16'h	20e3;
65297	:douta	=	16'h	20e3;
65298	:douta	=	16'h	20e3;
65299	:douta	=	16'h	20e3;
65300	:douta	=	16'h	28e3;
65301	:douta	=	16'h	28e3;
65302	:douta	=	16'h	2903;
65303	:douta	=	16'h	28e3;
65304	:douta	=	16'h	3103;
65305	:douta	=	16'h	3124;
65306	:douta	=	16'h	3123;
65307	:douta	=	16'h	3124;
65308	:douta	=	16'h	3944;
65309	:douta	=	16'h	3924;
65310	:douta	=	16'h	3944;
65311	:douta	=	16'h	4144;
65312	:douta	=	16'h	4164;
65313	:douta	=	16'h	4164;
65314	:douta	=	16'h	4165;
65315	:douta	=	16'h	4185;
65316	:douta	=	16'h	4985;
65317	:douta	=	16'h	49c6;
65318	:douta	=	16'h	4228;
65319	:douta	=	16'h	1084;
65320	:douta	=	16'h	3944;
65321	:douta	=	16'h	59c5;
65322	:douta	=	16'h	59e4;
65323	:douta	=	16'h	59e4;
65324	:douta	=	16'h	59e4;
65325	:douta	=	16'h	6205;
65326	:douta	=	16'h	6a25;
65327	:douta	=	16'h	6a25;
65328	:douta	=	16'h	7266;
65329	:douta	=	16'h	7266;
65330	:douta	=	16'h	7244;
65331	:douta	=	16'h	94f4;
65332	:douta	=	16'h	b5b4;
65333	:douta	=	16'h	7a66;
65334	:douta	=	16'h	7aa6;
65335	:douta	=	16'h	82a7;
65336	:douta	=	16'h	82a7;
65337	:douta	=	16'h	82c7;
65338	:douta	=	16'h	8ac7;
65339	:douta	=	16'h	82c6;
65340	:douta	=	16'h	8ae6;
65341	:douta	=	16'h	8ae6;
65342	:douta	=	16'h	8ae7;
65343	:douta	=	16'h	8b07;
65344	:douta	=	16'h	9308;
65345	:douta	=	16'h	9308;
65346	:douta	=	16'h	9328;
65347	:douta	=	16'h	9328;
65348	:douta	=	16'h	9328;
65349	:douta	=	16'h	9348;
65350	:douta	=	16'h	9348;
65351	:douta	=	16'h	9b48;
65352	:douta	=	16'h	9b69;
65353	:douta	=	16'h	9b69;
65354	:douta	=	16'h	9b68;
65355	:douta	=	16'h	9b48;
65356	:douta	=	16'h	a369;
65357	:douta	=	16'h	a369;
65358	:douta	=	16'h	a388;
65359	:douta	=	16'h	a388;
65360	:douta	=	16'h	a3a8;
65361	:douta	=	16'h	abc8;
65362	:douta	=	16'h	aba8;
65363	:douta	=	16'h	b3e9;
65364	:douta	=	16'h	b3e9;
65365	:douta	=	16'h	b3e9;
65366	:douta	=	16'h	b409;
65367	:douta	=	16'h	b409;
65368	:douta	=	16'h	b409;
65369	:douta	=	16'h	b42a;
65370	:douta	=	16'h	bc2a;
65371	:douta	=	16'h	bc2a;
65372	:douta	=	16'h	bc2a;
65373	:douta	=	16'h	bc2a;
65374	:douta	=	16'h	bc2a;
65375	:douta	=	16'h	bc2a;
65376	:douta	=	16'h	c42a;
65377	:douta	=	16'h	bc2a;
65378	:douta	=	16'h	bc2a;
65379	:douta	=	16'h	c44a;
65380	:douta	=	16'h	c44a;
65381	:douta	=	16'h	c44a;
65382	:douta	=	16'h	c44a;
65383	:douta	=	16'h	c44a;
65384	:douta	=	16'h	c46b;
65385	:douta	=	16'h	c46b;
65386	:douta	=	16'h	c46a;
65387	:douta	=	16'h	c46a;
65388	:douta	=	16'h	c46a;
65389	:douta	=	16'h	c46a;
65390	:douta	=	16'h	c46a;
65391	:douta	=	16'h	c48a;
65392	:douta	=	16'h	cc6a;
65393	:douta	=	16'h	c46a;
65394	:douta	=	16'h	cc6a;
65395	:douta	=	16'h	c46a;
65396	:douta	=	16'h	c46a;
65397	:douta	=	16'h	c46a;
65398	:douta	=	16'h	cc8a;
65399	:douta	=	16'h	cc8a;
65400	:douta	=	16'h	cc8a;
65401	:douta	=	16'h	c48a;
65402	:douta	=	16'h	cc8a;
65403	:douta	=	16'h	c46a;
65404	:douta	=	16'h	c469;
65405	:douta	=	16'h	c489;
65406	:douta	=	16'h	c469;
65407	:douta	=	16'h	cc6a;
65408	:douta	=	16'h	c469;
65409	:douta	=	16'h	cc6a;
65410	:douta	=	16'h	cc8a;
65411	:douta	=	16'h	cc6a;
65412	:douta	=	16'h	c469;
65413	:douta	=	16'h	cc6a;
65414	:douta	=	16'h	cc6a;
65415	:douta	=	16'h	cc6a;
65416	:douta	=	16'h	cc6a;
65417	:douta	=	16'h	cc6a;
65418	:douta	=	16'h	c469;
65419	:douta	=	16'h	c469;
65420	:douta	=	16'h	cc6a;
65421	:douta	=	16'h	c469;
65422	:douta	=	16'h	c469;
65423	:douta	=	16'h	cc6a;
65424	:douta	=	16'h	cc6a;
65425	:douta	=	16'h	cc6a;
65426	:douta	=	16'h	cc6a;
65427	:douta	=	16'h	c46a;
65428	:douta	=	16'h	c46a;
65429	:douta	=	16'h	c46a;
65430	:douta	=	16'h	cc6a;
65431	:douta	=	16'h	cc6a;
65432	:douta	=	16'h	cc6a;
65433	:douta	=	16'h	cc6a;
65434	:douta	=	16'h	cc6a;
65435	:douta	=	16'h	cc6a;
65436	:douta	=	16'h	cc6a;
65437	:douta	=	16'h	cc6a;
65438	:douta	=	16'h	c469;
65439	:douta	=	16'h	c46a;
65440	:douta	=	16'h	cc6a;
65441	:douta	=	16'h	cc69;
65442	:douta	=	16'h	c46a;
65443	:douta	=	16'h	be16;
65444	:douta	=	16'h	de13;
65445	:douta	=	16'h	c44a;
65446	:douta	=	16'h	c46a;
65447	:douta	=	16'h	c469;
65448	:douta	=	16'h	c46a;
65449	:douta	=	16'h	c46a;
65450	:douta	=	16'h	c469;
65451	:douta	=	16'h	c469;
65452	:douta	=	16'h	c46a;
65453	:douta	=	16'h	c46a;
65454	:douta	=	16'h	c46a;
65455	:douta	=	16'h	c469;
65456	:douta	=	16'h	c469;
65457	:douta	=	16'h	c469;
65458	:douta	=	16'h	cc6a;
65459	:douta	=	16'h	c46a;
65460	:douta	=	16'h	c469;
65461	:douta	=	16'h	c44a;
65462	:douta	=	16'h	c44a;
65463	:douta	=	16'h	c44a;
65464	:douta	=	16'h	c44a;
65465	:douta	=	16'h	c44a;
65466	:douta	=	16'h	c44a;
65467	:douta	=	16'h	c44a;
65468	:douta	=	16'h	c44a;
65469	:douta	=	16'h	c44a;
65470	:douta	=	16'h	c44a;
65471	:douta	=	16'h	c44a;
65472	:douta	=	16'h	c44a;
65473	:douta	=	16'h	c42a;
65474	:douta	=	16'h	bc2a;
65475	:douta	=	16'h	c44a;
65476	:douta	=	16'h	c44a;
65477	:douta	=	16'h	c44a;
65478	:douta	=	16'h	bc2a;
65479	:douta	=	16'h	c42a;
65480	:douta	=	16'h	c42a;
65481	:douta	=	16'h	bc2a;
65482	:douta	=	16'h	bc2a;
65483	:douta	=	16'h	bc2a;
65484	:douta	=	16'h	bc0a;
65485	:douta	=	16'h	bc2a;
65486	:douta	=	16'h	bc2a;
65487	:douta	=	16'h	bc2a;
65488	:douta	=	16'h	bc0a;
65489	:douta	=	16'h	bc0a;
65490	:douta	=	16'h	bc0a;
65491	:douta	=	16'h	bc0a;
65492	:douta	=	16'h	bc0a;
65493	:douta	=	16'h	bc0a;
65494	:douta	=	16'h	bc09;
65495	:douta	=	16'h	bc09;
65496	:douta	=	16'h	bc0a;
65497	:douta	=	16'h	b40a;
65498	:douta	=	16'h	bc0a;
65499	:douta	=	16'h	b40a;
65500	:douta	=	16'h	b3ea;
65501	:douta	=	16'h	b3ea;
65502	:douta	=	16'h	b40a;
65503	:douta	=	16'h	b3ea;
65504	:douta	=	16'h	b40a;
65505	:douta	=	16'h	b3e9;
65506	:douta	=	16'h	b3ea;
65507	:douta	=	16'h	b3ea;
65508	:douta	=	16'h	b3e9;
65509	:douta	=	16'h	abc9;
65510	:douta	=	16'h	b3ca;
65511	:douta	=	16'h	abca;
65512	:douta	=	16'h	abca;
65513	:douta	=	16'h	b3ca;
65514	:douta	=	16'h	b3ca;
65515	:douta	=	16'h	abca;
65516	:douta	=	16'h	aba9;
65517	:douta	=	16'h	abca;
65518	:douta	=	16'h	aba9;
65519	:douta	=	16'h	aba9;
65520	:douta	=	16'h	abaa;
65521	:douta	=	16'h	abaa;
65522	:douta	=	16'h	abaa;
65523	:douta	=	16'h	abaa;
65524	:douta	=	16'h	abaa;
65525	:douta	=	16'h	abaa;
65526	:douta	=	16'h	abaa;
65527	:douta	=	16'h	ab89;
65528	:douta	=	16'h	a389;
65529	:douta	=	16'h	a389;
65530	:douta	=	16'h	a389;
65531	:douta	=	16'h	a389;
65532	:douta	=	16'h	a38a;
65533	:douta	=	16'h	a369;
65534	:douta	=	16'h	a38a;
65535	:douta	=	16'h	a369;
default :douta  =	16'h	0000;
endcase
end


endmodule 
